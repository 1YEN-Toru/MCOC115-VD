
module mcss_alu
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_206 ,
    DI,
    S,
    \rgf_c0bus_wb[4]_i_17 ,
    \rgf_c0bus_wb[4]_i_17_0 ,
    \rgf_c0bus_wb[8]_i_5 ,
    \rgf_c0bus_wb[8]_i_5_0 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \sr[6]_i_8 ,
    \sr[6]_i_8_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_206 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb[4]_i_17 ;
  input [3:0]\rgf_c0bus_wb[4]_i_17_0 ;
  input [3:0]\rgf_c0bus_wb[8]_i_5 ;
  input [3:0]\rgf_c0bus_wb[8]_i_5_0 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_8 ;
  input [1:0]\sr[6]_i_8_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb[4]_i_17 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_17_0 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_5 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_5_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire \sr[4]_i_206 ;
  wire [0:0]\sr[6]_i_8 ;
  wire [1:0]\sr[6]_i_8_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire [3:0]tout__1_carry__1_i_8;
  wire [3:0]tout__1_carry__2_i_8;
  wire [0:0]tout__1_carry__3_i_3__0;

  mcss_alu_art_52 art
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c0bus_wb[4]_i_17 (\rgf_c0bus_wb[4]_i_17 ),
        .\rgf_c0bus_wb[4]_i_17_0 (\rgf_c0bus_wb[4]_i_17_0 ),
        .\rgf_c0bus_wb[8]_i_5 (\rgf_c0bus_wb[8]_i_5 ),
        .\rgf_c0bus_wb[8]_i_5_0 (\rgf_c0bus_wb[8]_i_5_0 ),
        .\rgf_c0bus_wb_reg[15] (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15]_0 ),
        .\sr[4]_i_206 (\sr[4]_i_206 ),
        .\sr[6]_i_8 (\sr[6]_i_8 ),
        .\sr[6]_i_8_0 (\sr[6]_i_8_0 ),
        .tout__1_carry__0_i_8(tout__1_carry__0_i_8),
        .tout__1_carry__1_i_8(tout__1_carry__1_i_8),
        .tout__1_carry__2_i_8(tout__1_carry__2_i_8),
        .tout__1_carry__3_i_3__0(tout__1_carry__3_i_3__0));
endmodule

(* ORIG_REF_NAME = "mcss_alu" *) 
module mcss_alu_0
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3,
    \sr[4]_i_123 ,
    DI,
    S,
    \rgf_c1bus_wb[4]_i_5 ,
    \rgf_c1bus_wb[4]_i_5_0 ,
    \rgf_c1bus_wb[8]_i_4 ,
    \rgf_c1bus_wb[8]_i_4_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_2 ,
    \sr[6]_i_2_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_123 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb[4]_i_5 ;
  input [3:0]\rgf_c1bus_wb[4]_i_5_0 ;
  input [3:0]\rgf_c1bus_wb[8]_i_4 ;
  input [3:0]\rgf_c1bus_wb[8]_i_4_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_2 ;
  input [1:0]\sr[6]_i_2_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb[4]_i_5 ;
  wire [3:0]\rgf_c1bus_wb[4]_i_5_0 ;
  wire [3:0]\rgf_c1bus_wb[8]_i_4 ;
  wire [3:0]\rgf_c1bus_wb[8]_i_4_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire \sr[4]_i_123 ;
  wire [0:0]\sr[6]_i_2 ;
  wire [1:0]\sr[6]_i_2_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire [0:0]tout__1_carry__3_i_3;

  mcss_alu_art art
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c1bus_wb[4]_i_5 (\rgf_c1bus_wb[4]_i_5 ),
        .\rgf_c1bus_wb[4]_i_5_0 (\rgf_c1bus_wb[4]_i_5_0 ),
        .\rgf_c1bus_wb[8]_i_4 (\rgf_c1bus_wb[8]_i_4 ),
        .\rgf_c1bus_wb[8]_i_4_0 (\rgf_c1bus_wb[8]_i_4_0 ),
        .\rgf_c1bus_wb_reg[15] (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15]_0 ),
        .\sr[4]_i_123 (\sr[4]_i_123 ),
        .\sr[6]_i_2 (\sr[6]_i_2 ),
        .\sr[6]_i_2_0 (\sr[6]_i_2_0 ),
        .tout__1_carry__0_i_8__0(tout__1_carry__0_i_8__0),
        .tout__1_carry__1_i_8__0(tout__1_carry__1_i_8__0),
        .tout__1_carry__2_i_8__0(tout__1_carry__2_i_8__0),
        .tout__1_carry__3_i_3(tout__1_carry__3_i_3));
endmodule

module mcss_alu_add
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3,
    \sr[4]_i_123_0 ,
    DI,
    S,
    \rgf_c1bus_wb[4]_i_5 ,
    \rgf_c1bus_wb[4]_i_5_0 ,
    \rgf_c1bus_wb[8]_i_4 ,
    \rgf_c1bus_wb[8]_i_4_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_2 ,
    \sr[6]_i_2_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_123_0 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb[4]_i_5 ;
  input [3:0]\rgf_c1bus_wb[4]_i_5_0 ;
  input [3:0]\rgf_c1bus_wb[8]_i_4 ;
  input [3:0]\rgf_c1bus_wb[8]_i_4_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_2 ;
  input [1:0]\sr[6]_i_2_0 ;

  wire \<const0> ;
  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb[4]_i_5 ;
  wire [3:0]\rgf_c1bus_wb[4]_i_5_0 ;
  wire [3:0]\rgf_c1bus_wb[8]_i_4 ;
  wire [3:0]\rgf_c1bus_wb[8]_i_4_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire \sr[4]_i_122_n_0 ;
  wire \sr[4]_i_123_0 ;
  wire \sr[4]_i_123_n_0 ;
  wire \sr[4]_i_182_n_0 ;
  wire [0:0]\sr[6]_i_2 ;
  wire [1:0]\sr[6]_i_2_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire tout__1_carry__0_n_0;
  wire tout__1_carry__0_n_1;
  wire tout__1_carry__0_n_2;
  wire tout__1_carry__0_n_3;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire tout__1_carry__1_n_0;
  wire tout__1_carry__1_n_1;
  wire tout__1_carry__1_n_2;
  wire tout__1_carry__1_n_3;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire tout__1_carry__2_n_0;
  wire tout__1_carry__2_n_1;
  wire tout__1_carry__2_n_2;
  wire tout__1_carry__2_n_3;
  wire [0:0]tout__1_carry__3_i_3;
  wire tout__1_carry__3_n_3;
  wire tout__1_carry_n_0;
  wire tout__1_carry_n_1;
  wire tout__1_carry_n_2;
  wire tout__1_carry_n_3;
  wire [3:0]NLW_tout__1_carry__3_O_UNCONNECTED;

  GND GND
       (.G(\<const0> ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_122 
       (.I0(O[1]),
        .I1(O[2]),
        .I2(tout__1_carry__0_i_8__0[2]),
        .I3(tout__1_carry__2_i_8__0[1]),
        .O(\sr[4]_i_122_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_123 
       (.I0(tout__1_carry__2_i_8__0[0]),
        .I1(tout__1_carry__1_i_8__0[0]),
        .I2(tout__1_carry__2_i_8__0[3]),
        .I3(tout__1_carry__2_i_8__0[2]),
        .I4(\sr[4]_i_182_n_0 ),
        .O(\sr[4]_i_123_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_182 
       (.I0(O[0]),
        .I1(tout__1_carry__0_i_8__0[1]),
        .I2(tout__1_carry__0_i_8__0[3]),
        .I3(tout__1_carry__1_i_8__0[3]),
        .O(\sr[4]_i_182_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_47 
       (.I0(\sr[4]_i_122_n_0 ),
        .I1(O[3]),
        .I2(tout__1_carry__1_i_8__0[1]),
        .I3(tout__1_carry__0_i_8__0[0]),
        .I4(tout__1_carry__1_i_8__0[2]),
        .I5(\sr[4]_i_123_n_0 ),
        .O(\sr[4]_i_123_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry
       (.CI(\<const0> ),
        .CO({tout__1_carry_n_0,tout__1_carry_n_1,tout__1_carry_n_2,tout__1_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({DI,\<const0> }),
        .O(O),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__0
       (.CI(tout__1_carry_n_0),
        .CO({tout__1_carry__0_n_0,tout__1_carry__0_n_1,tout__1_carry__0_n_2,tout__1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb[4]_i_5 ),
        .O(tout__1_carry__0_i_8__0),
        .S(\rgf_c1bus_wb[4]_i_5_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__1
       (.CI(tout__1_carry__0_n_0),
        .CO({tout__1_carry__1_n_0,tout__1_carry__1_n_1,tout__1_carry__1_n_2,tout__1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb[8]_i_4 ),
        .O(tout__1_carry__1_i_8__0),
        .S(\rgf_c1bus_wb[8]_i_4_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__2
       (.CI(tout__1_carry__1_n_0),
        .CO({tout__1_carry__2_n_0,tout__1_carry__2_n_1,tout__1_carry__2_n_2,tout__1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c1bus_wb_reg[15] ),
        .O(tout__1_carry__2_i_8__0),
        .S(\rgf_c1bus_wb_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__3
       (.CI(tout__1_carry__2_n_0),
        .CO(tout__1_carry__3_n_3),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_2 }),
        .O({tout__1_carry__3_i_3,NLW_tout__1_carry__3_O_UNCONNECTED[0]}),
        .S({\<const0> ,\<const0> ,\sr[6]_i_2_0 }));
endmodule

(* ORIG_REF_NAME = "mcss_alu_add" *) 
module mcss_alu_add_53
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_206_0 ,
    DI,
    S,
    \rgf_c0bus_wb[4]_i_17 ,
    \rgf_c0bus_wb[4]_i_17_0 ,
    \rgf_c0bus_wb[8]_i_5 ,
    \rgf_c0bus_wb[8]_i_5_0 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \sr[6]_i_8 ,
    \sr[6]_i_8_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_206_0 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb[4]_i_17 ;
  input [3:0]\rgf_c0bus_wb[4]_i_17_0 ;
  input [3:0]\rgf_c0bus_wb[8]_i_5 ;
  input [3:0]\rgf_c0bus_wb[8]_i_5_0 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_8 ;
  input [1:0]\sr[6]_i_8_0 ;

  wire \<const0> ;
  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb[4]_i_17 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_17_0 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_5 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_5_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire \sr[4]_i_205_n_0 ;
  wire \sr[4]_i_206_0 ;
  wire \sr[4]_i_206_n_0 ;
  wire \sr[4]_i_233_n_0 ;
  wire [0:0]\sr[6]_i_8 ;
  wire [1:0]\sr[6]_i_8_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire tout__1_carry__0_n_0;
  wire tout__1_carry__0_n_1;
  wire tout__1_carry__0_n_2;
  wire tout__1_carry__0_n_3;
  wire [3:0]tout__1_carry__1_i_8;
  wire tout__1_carry__1_n_0;
  wire tout__1_carry__1_n_1;
  wire tout__1_carry__1_n_2;
  wire tout__1_carry__1_n_3;
  wire [3:0]tout__1_carry__2_i_8;
  wire tout__1_carry__2_n_0;
  wire tout__1_carry__2_n_1;
  wire tout__1_carry__2_n_2;
  wire tout__1_carry__2_n_3;
  wire [0:0]tout__1_carry__3_i_3__0;
  wire tout__1_carry__3_n_3;
  wire tout__1_carry_n_0;
  wire tout__1_carry_n_1;
  wire tout__1_carry_n_2;
  wire tout__1_carry_n_3;
  wire [3:0]NLW_tout__1_carry__3_O_UNCONNECTED;

  GND GND
       (.G(\<const0> ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_152 
       (.I0(\sr[4]_i_205_n_0 ),
        .I1(tout__1_carry__1_i_8[1]),
        .I2(tout__1_carry__2_i_8[3]),
        .I3(tout__1_carry__0_i_8[3]),
        .I4(tout__1_carry__1_i_8[3]),
        .I5(\sr[4]_i_206_n_0 ),
        .O(\sr[4]_i_206_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_205 
       (.I0(O[3]),
        .I1(tout__1_carry__2_i_8[1]),
        .I2(O[2]),
        .I3(tout__1_carry__0_i_8[1]),
        .O(\sr[4]_i_205_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_206 
       (.I0(tout__1_carry__2_i_8[2]),
        .I1(tout__1_carry__0_i_8[2]),
        .I2(tout__1_carry__1_i_8[0]),
        .I3(O[1]),
        .I4(\sr[4]_i_233_n_0 ),
        .O(\sr[4]_i_206_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_233 
       (.I0(tout__1_carry__1_i_8[2]),
        .I1(tout__1_carry__2_i_8[0]),
        .I2(O[0]),
        .I3(tout__1_carry__0_i_8[0]),
        .O(\sr[4]_i_233_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry
       (.CI(\<const0> ),
        .CO({tout__1_carry_n_0,tout__1_carry_n_1,tout__1_carry_n_2,tout__1_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({DI,\<const0> }),
        .O(O),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__0
       (.CI(tout__1_carry_n_0),
        .CO({tout__1_carry__0_n_0,tout__1_carry__0_n_1,tout__1_carry__0_n_2,tout__1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb[4]_i_17 ),
        .O(tout__1_carry__0_i_8),
        .S(\rgf_c0bus_wb[4]_i_17_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__1
       (.CI(tout__1_carry__0_n_0),
        .CO({tout__1_carry__1_n_0,tout__1_carry__1_n_1,tout__1_carry__1_n_2,tout__1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb[8]_i_5 ),
        .O(tout__1_carry__1_i_8),
        .S(\rgf_c0bus_wb[8]_i_5_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__2
       (.CI(tout__1_carry__1_n_0),
        .CO({tout__1_carry__2_n_0,tout__1_carry__2_n_1,tout__1_carry__2_n_2,tout__1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\rgf_c0bus_wb_reg[15] ),
        .O(tout__1_carry__2_i_8),
        .S(\rgf_c0bus_wb_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 tout__1_carry__3
       (.CI(tout__1_carry__2_n_0),
        .CO(tout__1_carry__3_n_3),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_8 }),
        .O({tout__1_carry__3_i_3__0,NLW_tout__1_carry__3_O_UNCONNECTED[0]}),
        .S({\<const0> ,\<const0> ,\sr[6]_i_8_0 }));
endmodule

module mcss_alu_art
   (O,
    tout__1_carry__0_i_8__0,
    tout__1_carry__1_i_8__0,
    tout__1_carry__2_i_8__0,
    tout__1_carry__3_i_3,
    \sr[4]_i_123 ,
    DI,
    S,
    \rgf_c1bus_wb[4]_i_5 ,
    \rgf_c1bus_wb[4]_i_5_0 ,
    \rgf_c1bus_wb[8]_i_4 ,
    \rgf_c1bus_wb[8]_i_4_0 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    \sr[6]_i_2 ,
    \sr[6]_i_2_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8__0;
  output [3:0]tout__1_carry__1_i_8__0;
  output [3:0]tout__1_carry__2_i_8__0;
  output [0:0]tout__1_carry__3_i_3;
  output \sr[4]_i_123 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c1bus_wb[4]_i_5 ;
  input [3:0]\rgf_c1bus_wb[4]_i_5_0 ;
  input [3:0]\rgf_c1bus_wb[8]_i_4 ;
  input [3:0]\rgf_c1bus_wb[8]_i_4_0 ;
  input [3:0]\rgf_c1bus_wb_reg[15] ;
  input [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_2 ;
  input [1:0]\sr[6]_i_2_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c1bus_wb[4]_i_5 ;
  wire [3:0]\rgf_c1bus_wb[4]_i_5_0 ;
  wire [3:0]\rgf_c1bus_wb[8]_i_4 ;
  wire [3:0]\rgf_c1bus_wb[8]_i_4_0 ;
  wire [3:0]\rgf_c1bus_wb_reg[15] ;
  wire [3:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire \sr[4]_i_123 ;
  wire [0:0]\sr[6]_i_2 ;
  wire [1:0]\sr[6]_i_2_0 ;
  wire [3:0]tout__1_carry__0_i_8__0;
  wire [3:0]tout__1_carry__1_i_8__0;
  wire [3:0]tout__1_carry__2_i_8__0;
  wire [0:0]tout__1_carry__3_i_3;

  mcss_alu_add add
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c1bus_wb[4]_i_5 (\rgf_c1bus_wb[4]_i_5 ),
        .\rgf_c1bus_wb[4]_i_5_0 (\rgf_c1bus_wb[4]_i_5_0 ),
        .\rgf_c1bus_wb[8]_i_4 (\rgf_c1bus_wb[8]_i_4 ),
        .\rgf_c1bus_wb[8]_i_4_0 (\rgf_c1bus_wb[8]_i_4_0 ),
        .\rgf_c1bus_wb_reg[15] (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15]_0 ),
        .\sr[4]_i_123_0 (\sr[4]_i_123 ),
        .\sr[6]_i_2 (\sr[6]_i_2 ),
        .\sr[6]_i_2_0 (\sr[6]_i_2_0 ),
        .tout__1_carry__0_i_8__0(tout__1_carry__0_i_8__0),
        .tout__1_carry__1_i_8__0(tout__1_carry__1_i_8__0),
        .tout__1_carry__2_i_8__0(tout__1_carry__2_i_8__0),
        .tout__1_carry__3_i_3(tout__1_carry__3_i_3));
endmodule

(* ORIG_REF_NAME = "mcss_alu_art" *) 
module mcss_alu_art_52
   (O,
    tout__1_carry__0_i_8,
    tout__1_carry__1_i_8,
    tout__1_carry__2_i_8,
    tout__1_carry__3_i_3__0,
    \sr[4]_i_206 ,
    DI,
    S,
    \rgf_c0bus_wb[4]_i_17 ,
    \rgf_c0bus_wb[4]_i_17_0 ,
    \rgf_c0bus_wb[8]_i_5 ,
    \rgf_c0bus_wb[8]_i_5_0 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \sr[6]_i_8 ,
    \sr[6]_i_8_0 );
  output [3:0]O;
  output [3:0]tout__1_carry__0_i_8;
  output [3:0]tout__1_carry__1_i_8;
  output [3:0]tout__1_carry__2_i_8;
  output [0:0]tout__1_carry__3_i_3__0;
  output \sr[4]_i_206 ;
  input [2:0]DI;
  input [3:0]S;
  input [3:0]\rgf_c0bus_wb[4]_i_17 ;
  input [3:0]\rgf_c0bus_wb[4]_i_17_0 ;
  input [3:0]\rgf_c0bus_wb[8]_i_5 ;
  input [3:0]\rgf_c0bus_wb[8]_i_5_0 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [0:0]\sr[6]_i_8 ;
  input [1:0]\sr[6]_i_8_0 ;

  wire [2:0]DI;
  wire [3:0]O;
  wire [3:0]S;
  wire [3:0]\rgf_c0bus_wb[4]_i_17 ;
  wire [3:0]\rgf_c0bus_wb[4]_i_17_0 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_5 ;
  wire [3:0]\rgf_c0bus_wb[8]_i_5_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire [3:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire \sr[4]_i_206 ;
  wire [0:0]\sr[6]_i_8 ;
  wire [1:0]\sr[6]_i_8_0 ;
  wire [3:0]tout__1_carry__0_i_8;
  wire [3:0]tout__1_carry__1_i_8;
  wire [3:0]tout__1_carry__2_i_8;
  wire [0:0]tout__1_carry__3_i_3__0;

  mcss_alu_add_53 add
       (.DI(DI),
        .O(O),
        .S(S),
        .\rgf_c0bus_wb[4]_i_17 (\rgf_c0bus_wb[4]_i_17 ),
        .\rgf_c0bus_wb[4]_i_17_0 (\rgf_c0bus_wb[4]_i_17_0 ),
        .\rgf_c0bus_wb[8]_i_5 (\rgf_c0bus_wb[8]_i_5 ),
        .\rgf_c0bus_wb[8]_i_5_0 (\rgf_c0bus_wb[8]_i_5_0 ),
        .\rgf_c0bus_wb_reg[15] (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15]_0 ),
        .\sr[4]_i_206_0 (\sr[4]_i_206 ),
        .\sr[6]_i_8 (\sr[6]_i_8 ),
        .\sr[6]_i_8_0 (\sr[6]_i_8_0 ),
        .tout__1_carry__0_i_8(tout__1_carry__0_i_8),
        .tout__1_carry__1_i_8(tout__1_carry__1_i_8),
        .tout__1_carry__2_i_8(tout__1_carry__2_i_8),
        .tout__1_carry__3_i_3__0(tout__1_carry__3_i_3__0));
endmodule

module mcss_fch
   (.out({ir0[15],ir0[14],ir0[13],ir0[12],ir0[11],ir0[10],ir0[9],ir0[7],ir0[2],ir0[1],ir0[0]}),
    .rst_n_fl_reg_0({ir1[15],ir1[14],ir1[13],ir1[12],ir1[11],ir1[10],ir1[9],ir1[5],ir1[2],ir1[1],ir1[0]}),
    fadr,
    fch_irq_req_fl,
    fch_term,
    O,
    \pc_reg[15] ,
    ctl_bcc_take0_fl,
    ctl_bcc_take1_fl,
    \bdatr[15] ,
    \cbus_i[15] ,
    p_2_in,
    rst_n_fl_reg_1,
    \stat_reg[2] ,
    \stat_reg[2]_0 ,
    \stat_reg[2]_1 ,
    \stat_reg[2]_2 ,
    \sr_reg[15] ,
    \stat_reg[2]_3 ,
    tout__1_carry_i_11_0,
    \tr_reg[4] ,
    rst_n_0,
    b1bus_sr,
    b1bus_sel_cr,
    rgf_selc1_stat_reg,
    \stat[2]_i_4 ,
    \stat_reg[0] ,
    \stat_reg[1] ,
    \sp_reg[15] ,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    fch_leir_nir_reg,
    \stat_reg[1]_0 ,
    \stat_reg[2]_4 ,
    bdatw,
    \bcmd[2]_INST_0_0 ,
    \bcmd[1]_INST_0_0 ,
    \tr_reg[4]_0 ,
    \rgf_c1bus_wb[15]_i_14_0 ,
    \stat_reg[2]_5 ,
    \stat_reg[2]_6 ,
    \stat_reg[2]_7 ,
    \bdatw[8]_INST_0_i_16_0 ,
    \bdatw[9]_INST_0_i_16_0 ,
    \stat_reg[2]_8 ,
    \bdatw[8]_INST_0_i_16_1 ,
    \sr_reg[6] ,
    \tr_reg[0] ,
    \bdatw[8]_INST_0_i_16_2 ,
    \rgf_c1bus_wb[15]_i_14_1 ,
    \badr[14]_INST_0_i_1 ,
    \bdatw[11]_INST_0_i_16_0 ,
    \stat_reg[2]_9 ,
    \tr_reg[0]_0 ,
    \stat_reg[0]_2 ,
    \stat_reg[2]_10 ,
    \stat_reg[1]_1 ,
    bbus_o,
    \stat_reg[0]_3 ,
    \rgf_c0bus_wb[15]_i_7_0 ,
    \stat_reg[1]_2 ,
    \bbus_o[2]_INST_0_i_1_0 ,
    \bbus_o[3]_INST_0_i_1_0 ,
    \bbus_o[1]_INST_0_i_1_0 ,
    \rgf_c0bus_wb[11]_i_11_0 ,
    \rgf_c0bus_wb[11]_i_3_0 ,
    \rgf_c0bus_wb[13]_i_10_0 ,
    \badr[15]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \bbus_o[0]_INST_0_i_1_0 ,
    \sr_reg[6]_0 ,
    \bbus_o[1]_INST_0_i_1_1 ,
    \bbus_o[1]_INST_0_i_1_2 ,
    \tr_reg[0]_1 ,
    ctl_sela0_rn,
    \stat_reg[0]_4 ,
    \stat_reg[2]_11 ,
    ccmd,
    \stat_reg[0]_5 ,
    \stat_reg[1]_3 ,
    \stat_reg[0]_6 ,
    \sr_reg[5] ,
    ctl_selb0_0,
    \stat_reg[0]_7 ,
    \stat_reg[0]_8 ,
    \stat_reg[0]_9 ,
    \stat_reg[0]_10 ,
    \stat_reg[1]_4 ,
    rst_n_fl_reg_2,
    ctl_selb0_rn,
    \stat_reg[1]_5 ,
    rst_n_fl_reg_3,
    \stat_reg[0]_11 ,
    ctl_selb1_0,
    \stat_reg[0]_12 ,
    rst_n_fl_reg_4,
    rst_n_fl_reg_5,
    rst_n_fl_reg_6,
    \stat_reg[0]_13 ,
    \stat_reg[0]_14 ,
    fch_leir_nir_reg_0,
    rst_n_fl_reg_7,
    rst_n_fl_reg_8,
    fch_leir_nir_reg_1,
    fch_leir_nir_reg_2,
    fch_leir_nir_reg_3,
    fch_leir_nir_reg_4,
    fch_leir_nir_reg_5,
    fch_leir_nir_reg_6,
    fch_leir_nir_reg_7,
    rst_n_fl_reg_9,
    \stat_reg[1]_6 ,
    \stat_reg[0]_15 ,
    ctl_sela0,
    \stat_reg[2]_12 ,
    \sr_reg[4] ,
    ctl_selb1_rn,
    \stat_reg[0]_16 ,
    \stat_reg[0]_17 ,
    \stat_reg[0]_18 ,
    ir0_id,
    fch_memacc1,
    .fdatx_5_sp_1(fdatx_5_sn_1),
    .fdatx_14_sp_1(fdatx_14_sn_1),
    .fdat_0_sp_1(fdat_0_sn_1),
    .fdat_12_sp_1(fdat_12_sn_1),
    .fdat_5_sp_1(fdat_5_sn_1),
    \stat_reg[1]_7 ,
    \sr_reg[4]_0 ,
    \stat_reg[2]_13 ,
    abus_o,
    \sr_reg[0] ,
    \stat_reg[0]_19 ,
    \sr_reg[0]_0 ,
    \sr_reg[0]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \grn_reg[4] ,
    \stat_reg[0]_20 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \sr_reg[0]_4 ,
    \stat_reg[2]_14 ,
    \stat_reg[2]_15 ,
    \stat_reg[2]_16 ,
    \sr_reg[0]_5 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[0]_11 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[0]_17 ,
    \sr_reg[0]_18 ,
    \sr_reg[0]_19 ,
    \grn_reg[4]_0 ,
    \stat_reg[0]_21 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \stat_reg[2]_17 ,
    \stat_reg[0]_22 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[4]_2 ,
    \stat_reg[0]_23 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_5 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_6 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_7 ,
    \sr_reg[0]_20 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[0]_23 ,
    \sr_reg[0]_24 ,
    \sr_reg[0]_25 ,
    \sr_reg[0]_26 ,
    \sr_reg[0]_27 ,
    \sr_reg[0]_28 ,
    \sr_reg[0]_29 ,
    \sr_reg[0]_30 ,
    \sr_reg[0]_31 ,
    \sr_reg[0]_32 ,
    \sr_reg[0]_33 ,
    \sr_reg[0]_34 ,
    \sr_reg[0]_35 ,
    \sr_reg[1] ,
    \sr_reg[1]_0 ,
    \sr_reg[1]_1 ,
    \sr_reg[1]_2 ,
    \sr_reg[1]_3 ,
    \sr_reg[1]_4 ,
    \sr_reg[1]_5 ,
    \sr_reg[1]_6 ,
    \sr_reg[1]_7 ,
    \sr_reg[1]_8 ,
    \sr_reg[1]_9 ,
    \sr_reg[1]_10 ,
    \sr_reg[1]_11 ,
    \sr_reg[1]_12 ,
    \sr_reg[1]_13 ,
    \stat_reg[2]_18 ,
    E,
    \stat_reg[0]_24 ,
    \stat_reg[0]_25 ,
    \stat_reg[0]_26 ,
    \stat_reg[0]_27 ,
    \stat_reg[0]_28 ,
    \stat_reg[0]_29 ,
    \stat_reg[0]_30 ,
    \stat_reg[0]_31 ,
    \stat_reg[0]_32 ,
    rst_n_fl_reg_10,
    rst_n_fl_reg_11,
    rst_n_fl_reg_12,
    \stat_reg[0]_33 ,
    \stat_reg[2]_19 ,
    \stat_reg[2]_20 ,
    fch_irq_req_fl_reg_0,
    a0bus_sel_cr,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4]_1 ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \tr_reg[15] ,
    b0bus_sr,
    \sr_reg[1]_14 ,
    \sr_reg[0]_36 ,
    \sr_reg[0]_37 ,
    \sr_reg[0]_38 ,
    \sr_reg[1]_15 ,
    \sr_reg[0]_39 ,
    \sr_reg[0]_40 ,
    \sr_reg[0]_41 ,
    \sr_reg[1]_16 ,
    \sr_reg[0]_42 ,
    \sr_reg[0]_43 ,
    \sr_reg[0]_44 ,
    \sr_reg[1]_17 ,
    \sr_reg[0]_45 ,
    \sr_reg[0]_46 ,
    \sr_reg[0]_47 ,
    \sr_reg[1]_18 ,
    \sr_reg[0]_48 ,
    \sr_reg[0]_49 ,
    \sr_reg[0]_50 ,
    \sr_reg[1]_19 ,
    \sr_reg[0]_51 ,
    \sr_reg[0]_52 ,
    \sr_reg[0]_53 ,
    \rgf_c0bus_wb[15]_i_8_0 ,
    \stat_reg[0]_34 ,
    \stat_reg[0]_35 ,
    \stat_reg[0]_36 ,
    \stat_reg[0]_37 ,
    \stat_reg[0]_38 ,
    \stat_reg[0]_39 ,
    \stat_reg[0]_40 ,
    \stat_reg[0]_41 ,
    \stat_reg[0]_42 ,
    \stat_reg[0]_43 ,
    \stat_reg[0]_44 ,
    badr,
    tout__1_carry_i_1__0_0,
    DI,
    \badr[15]_INST_0_i_1 ,
    \badr[15]_INST_0_i_1_0 ,
    \badr[15]_INST_0_i_1_1 ,
    \badr[14]_INST_0_i_2 ,
    \badr[15]_INST_0_i_2_0 ,
    \badr[15]_INST_0_i_2_1 ,
    \badr[15]_INST_0_i_2_2 ,
    a1bus_sr,
    a1bus_sel_cr,
    \sr_reg[0]_54 ,
    \sr_reg[1]_20 ,
    \sr_reg[0]_55 ,
    \sr_reg[0]_56 ,
    \badr[2]_INST_0_i_2 ,
    tout__1_carry_i_1_0,
    \badr[6]_INST_0_i_2 ,
    tout__1_carry__0_i_1_0,
    \badr[10]_INST_0_i_2 ,
    tout__1_carry__1_i_1_0,
    \badr[4]_INST_0_i_1 ,
    tout__1_carry__0_i_3__0_0,
    \pc0_reg[15]_0 ,
    \pc1_reg[15]_0 ,
    b0bus_sel_cr,
    \stat_reg[0]_45 ,
    b0bus_sel_0,
    \stat_reg[0]_46 ,
    a1bus_sel_0,
    \stat_reg[0]_47 ,
    \iv_reg[15] ,
    \tr_reg[15]_0 ,
    a0bus_sel_0,
    rgf_selc1_stat_reg_0,
    rgf_selc1_stat_reg_1,
    rgf_selc1_stat_reg_2,
    rgf_selc1_stat_reg_3,
    rgf_selc1_stat_reg_4,
    rgf_selc1_stat_reg_5,
    rgf_selc1_stat_reg_6,
    rgf_selc1_stat_reg_7,
    rgf_selc1_stat_reg_8,
    rgf_selc1_stat_reg_9,
    rgf_selc1_stat_reg_10,
    rgf_selc1_stat_reg_11,
    rgf_selc1_stat_reg_12,
    rgf_selc1_stat_reg_13,
    rgf_selc1_stat_reg_14,
    rgf_selc1_stat_reg_15,
    rgf_selc1_stat_reg_16,
    rgf_selc1_stat_reg_17,
    rgf_selc1_stat_reg_18,
    rgf_selc1_stat_reg_19,
    rgf_selc1_stat_reg_20,
    rgf_selc1_stat_reg_21,
    rgf_selc1_stat_reg_22,
    rgf_selc1_stat_reg_23,
    rgf_selc1_stat_reg_24,
    rgf_selc1_stat_reg_25,
    rgf_selc1_stat_reg_26,
    rgf_selc1_stat_reg_27,
    rgf_selc1_stat_reg_28,
    rgf_selc1_stat_reg_29,
    rgf_selc1_stat_reg_30,
    rgf_selc1_stat_reg_31,
    \sr_reg[0]_57 ,
    \sr_reg[0]_58 ,
    \sr_reg[0]_59 ,
    \sr_reg[1]_21 ,
    rst_n,
    clk,
    fch_irq_req,
    \pc0_reg[15]_1 ,
    S,
    \fadr[3] ,
    D,
    \pc1_reg[15]_1 ,
    ctl_bcc_take0_fl_reg_0,
    ctl_bcc_take1_fl_reg_0,
    \grn_reg[15] ,
    rgf_selc1_stat,
    Q,
    rgf_selc0_stat,
    \pc_reg[15]_0 ,
    \grn_reg[15]_0 ,
    \grn[15]_i_3__5 ,
    \sr[13]_i_5 ,
    \sr[13]_i_5_0 ,
    \sr_reg[4]_1 ,
    \sr_reg[5]_0 ,
    \sr_reg[15]_0 ,
    \sr_reg[6]_1 ,
    \pc_reg[15]_1 ,
    \pc_reg[14] ,
    \pc_reg[13] ,
    \sp_reg[15]_0 ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[1] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[2] ,
    \sp_reg[0] ,
    \sp_reg[0]_0 ,
    \sp[15]_i_2 ,
    \rgf_c1bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15]_0 ,
    a1bus_0,
    \bdatw[15] ,
    \stat_reg[0]_48 ,
    \bdatw[15]_0 ,
    \bdatw[15]_1 ,
    \bdatw[15]_2 ,
    \rgf_c1bus_wb_reg[14] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    \rgf_c1bus_wb[14]_i_3_0 ,
    \rgf_c1bus_wb_reg[13] ,
    \rgf_c1bus_wb[13]_i_5_0 ,
    bdatr,
    \rgf_c1bus_wb_reg[12] ,
    .bdatw_12_sp_1(bdatw_12_sn_1),
    \bdatw[12]_0 ,
    \rgf_c1bus_wb_reg[11] ,
    .bdatw_11_sp_1(bdatw_11_sn_1),
    \bdatw[11]_0 ,
    \rgf_c1bus_wb_reg[10] ,
    \sr[4]_i_52_0 ,
    .bdatw_10_sp_1(bdatw_10_sn_1),
    \bdatw[10]_0 ,
    \rgf_c1bus_wb_reg[9] ,
    .bdatw_9_sp_1(bdatw_9_sn_1),
    \bdatw[9]_0 ,
    \rgf_c1bus_wb_reg[8] ,
    .bdatw_8_sp_1(bdatw_8_sn_1),
    \bdatw[8]_0 ,
    \rgf_c1bus_wb[15]_i_10_0 ,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb_reg[7]_0 ,
    \rgf_c1bus_wb_reg[7]_1 ,
    \rgf_c1bus_wb_reg[6] ,
    \rgf_c1bus_wb_reg[6]_0 ,
    \rgf_c1bus_wb_reg[6]_1 ,
    \rgf_c1bus_wb[14]_i_3_1 ,
    .bdatw_6_sp_1(bdatw_6_sn_1),
    \rgf_c1bus_wb_reg[5] ,
    \rgf_c1bus_wb_reg[5]_0 ,
    \sr[4]_i_53_0 ,
    \sr[4]_i_53_1 ,
    tout__1_carry__0,
    .bdatw_5_sp_1(bdatw_5_sn_1),
    \sr[4]_i_10_0 ,
    \rgf_c1bus_wb_reg[13]_0 ,
    \rgf_c1bus_wb_reg[1] ,
    \rgf_c1bus_wb[9]_i_3_0 ,
    \rgf_c1bus_wb[9]_i_3_1 ,
    \sr[4]_i_9_0 ,
    \rgf_c1bus_wb_reg[15]_1 ,
    \sr[4]_i_41_0 ,
    \rgf_c1bus_wb_reg[3] ,
    \sr[4]_i_35_0 ,
    \rgf_c1bus_wb_reg[3]_0 ,
    \rgf_c1bus_wb_reg[3]_1 ,
    \sr[4]_i_91 ,
    \sr[4]_i_100_0 ,
    \sr[4]_i_10_1 ,
    \sr[4]_i_10_2 ,
    \rgf_c1bus_wb_reg[7]_2 ,
    \rgf_c1bus_wb_reg[11]_0 ,
    \sr[4]_i_35_1 ,
    \rgf_c1bus_wb[11]_i_6_0 ,
    \sr[4]_i_98_0 ,
    \sr[4]_i_98_1 ,
    \sr[4]_i_30_0 ,
    \sr[4]_i_30_1 ,
    \rgf_c1bus_wb_reg[8]_0 ,
    \rgf_c1bus_wb_reg[12]_0 ,
    \rgf_c1bus_wb_reg[4] ,
    \sr[4]_i_11_0 ,
    \rgf_c1bus_wb_reg[4]_0 ,
    \sr[6]_i_6_0 ,
    \rgf_c1bus_wb[4]_i_4_0 ,
    \rgf_c1bus_wb[4]_i_4_1 ,
    \rgf_c1bus_wb_reg[0] ,
    \sr[4]_i_36_0 ,
    \sr[4]_i_25_0 ,
    \rgf_c1bus_wb[4]_i_4_2 ,
    \rgf_c1bus_wb[4]_i_4_3 ,
    \rgf_c1bus_wb_reg[12]_1 ,
    \sr[4]_i_111_0 ,
    \sr[4]_i_36_1 ,
    \sr[4]_i_36_2 ,
    \rgf_c1bus_wb_reg[4]_1 ,
    \sr[6]_i_6_1 ,
    \rgf_c1bus_wb_reg[13]_1 ,
    \sr[4]_i_37_0 ,
    \sr[4]_i_39_0 ,
    \rgf_c1bus_wb[0]_i_4_0 ,
    \sr[4]_i_29_0 ,
    \rgf_c1bus_wb_reg[9]_0 ,
    \rgf_c1bus_wb[13]_i_2_0 ,
    \sr[4]_i_27_0 ,
    \rgf_c1bus_wb_reg[13]_2 ,
    \sr[4]_i_29_1 ,
    \sr[4]_i_29_2 ,
    \rgf_c1bus_wb[1]_i_2_0 ,
    \rgf_c1bus_wb_reg[2] ,
    \sr[4]_i_12_0 ,
    \rgf_c1bus_wb_reg[14]_1 ,
    \rgf_c1bus_wb_reg[14]_2 ,
    \sr[4]_i_29_3 ,
    \rgf_c1bus_wb_reg[10]_0 ,
    \sr[4]_i_44_0 ,
    \sr[4]_i_46_0 ,
    \sr[4]_i_43_0 ,
    \sr[4]_i_43_1 ,
    \rgf_c1bus_wb_reg[6]_2 ,
    \rgf_c1bus_wb_reg[6]_3 ,
    \sr[4]_i_43_2 ,
    \rgf_c1bus_wb_reg[14]_3 ,
    \sr[4]_i_46_1 ,
    \sr[4]_i_46_2 ,
    \rgf_c1bus_wb_reg[2]_0 ,
    \sr[4]_i_45_0 ,
    \sr[4]_i_34_0 ,
    \sr[4]_i_102_0 ,
    \rgf_c1bus_wb[9]_i_3_2 ,
    \rgf_c1bus_wb[15]_i_4_0 ,
    \sr[4]_i_33_0 ,
    \sr[4]_i_28_0 ,
    \sr[4]_i_28_1 ,
    \rgf_c1bus_wb_reg[7]_3 ,
    \rgf_c1bus_wb[11]_i_3_0 ,
    \sr[4]_i_100_1 ,
    \sr[4]_i_100_2 ,
    \rgf_c1bus_wb_reg[4]_2 ,
    \rgf_c1bus_wb_reg[13]_3 ,
    b1bus_b02,
    \rgf_c1bus_wb_reg[13]_4 ,
    \rgf_c1bus_wb_reg[13]_5 ,
    \sr[4]_i_102_1 ,
    \sr[4]_i_102_2 ,
    \sr[4]_i_102_3 ,
    \rgf_c1bus_wb[5]_i_9_0 ,
    \rgf_c1bus_wb[5]_i_9_1 ,
    \rgf_c1bus_wb[5]_i_9_2 ,
    \rgf_c1bus_wb_reg[1]_0 ,
    \rgf_c1bus_wb_reg[3]_2 ,
    \rgf_c1bus_wb[14]_i_28_0 ,
    \rgf_c1bus_wb[14]_i_28_1 ,
    \rgf_c1bus_wb[14]_i_28_2 ,
    \sr[6]_i_16 ,
    \sr[6]_i_16_0 ,
    \sr[6]_i_16_1 ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c0bus_wb_reg[15]_0 ,
    a0bus_0,
    \rgf_c0bus_wb_reg[14] ,
    .bbus_o_14_sp_1(bbus_o_14_sn_1),
    .bbus_o_13_sp_1(bbus_o_13_sn_1),
    \rgf_c0bus_wb_reg[12] ,
    \rgf_c0bus_wb_reg[11] ,
    \rgf_c0bus_wb_reg[11]_0 ,
    \sr[4]_i_72_0 ,
    \rgf_c0bus_wb_reg[10] ,
    \rgf_c0bus_wb_reg[10]_0 ,
    \rgf_c0bus_wb_reg[9] ,
    \rgf_c0bus_wb_reg[8] ,
    \sr[4]_i_71_0 ,
    \rgf_c0bus_wb_reg[10]_i_17_0 ,
    .bbus_o_7_sp_1(bbus_o_7_sn_1),
    cbus_i,
    \rgf_c0bus_wb_reg[7] ,
    \rgf_c0bus_wb_reg[7]_0 ,
    \sr[4]_i_69_0 ,
    \rgf_c0bus_wb_reg[10]_i_17_1 ,
    \rgf_c0bus_wb_reg[10]_i_17_2 ,
    .bbus_o_6_sp_1(bbus_o_6_sn_1),
    \rgf_c0bus_wb_reg[6] ,
    \sr[4]_i_70_0 ,
    \rgf_c0bus_wb_reg[5] ,
    \rgf_c0bus_wb_reg[10]_1 ,
    \sr[4]_i_6_0 ,
    \rgf_c0bus_wb_reg[7]_1 ,
    \sr[6]_i_5 ,
    \sr[4]_i_17_0 ,
    \rgf_c0bus_wb_reg[3] ,
    \rgf_c0bus_wb_reg[0] ,
    \rgf_c0bus_wb[0]_i_2_0 ,
    \sr[4]_i_66_0 ,
    \rgf_c0bus_wb[5]_i_2_0 ,
    \rgf_c0bus_wb_reg[2] ,
    \rgf_c0bus_wb_reg[2]_0 ,
    \rgf_c0bus_wb_reg[3]_0 ,
    \sr[4]_i_17_1 ,
    \sr[4]_i_18_0 ,
    \sr[4]_i_18_1 ,
    \sr[4]_i_18_2 ,
    \sr[4]_i_15_0 ,
    \rgf_c0bus_wb_reg[11]_1 ,
    \sr[4]_i_55_0 ,
    \rgf_c0bus_wb_reg[11]_2 ,
    \rgf_c0bus_wb_reg[11]_3 ,
    \rgf_c0bus_wb_reg[12]_0 ,
    \rgf_c0bus_wb_reg[13] ,
    \rgf_c0bus_wb_reg[14]_0 ,
    \sr[4]_i_16_0 ,
    \rgf_c0bus_wb[12]_i_3_0 ,
    \rgf_c0bus_wb[13]_i_2_0 ,
    \rgf_c0bus_wb_reg[4] ,
    \rgf_c0bus_wb_reg[4]_0 ,
    \rgf_c0bus_wb[12]_i_3_1 ,
    \rgf_c0bus_wb_reg[1] ,
    \rgf_c0bus_wb[5]_i_3_0 ,
    \sr[4]_i_67_0 ,
    \rgf_c0bus_wb_reg[8]_0 ,
    \rgf_c0bus_wb[1]_i_3_0 ,
    \rgf_c0bus_wb[9]_i_3_0 ,
    \rgf_c0bus_wb[10]_i_4_0 ,
    \rgf_c0bus_wb[10]_i_4_1 ,
    \rgf_c0bus_wb[11]_i_5_0 ,
    \rgf_c0bus_wb[13]_i_2_1 ,
    \rgf_c0bus_wb[13]_i_2_2 ,
    \sr[4]_i_58_0 ,
    \sr[4]_i_55_1 ,
    \sr[4]_i_55_2 ,
    \sr[4]_i_60_0 ,
    \sr[4]_i_65_0 ,
    \sr[4]_i_68_0 ,
    \rgf_c0bus_wb[9]_i_3_1 ,
    \rgf_c0bus_wb[5]_i_3_1 ,
    \rgf_c0bus_wb_reg[6]_0 ,
    \rgf_c0bus_wb_reg[6]_1 ,
    \rgf_c0bus_wb_reg[4]_1 ,
    \rgf_c0bus_wb_reg[4]_2 ,
    \rgf_c0bus_wb_reg[9]_0 ,
    \rgf_c0bus_wb_reg[9]_1 ,
    \rgf_c0bus_wb_reg[10]_2 ,
    \sr[4]_i_64_0 ,
    \sr[4]_i_60_1 ,
    \rgf_c0bus_wb_reg[10]_3 ,
    \rgf_c0bus_wb[4]_i_3_0 ,
    \rgf_c0bus_wb[4]_i_3_1 ,
    \rgf_c0bus_wb[5]_i_3_2 ,
    \sr[4]_i_68_1 ,
    \rgf_c0bus_wb[0]_i_2_1 ,
    \sr[4]_i_64_1 ,
    \sr[4]_i_60_2 ,
    \sr[4]_i_127_0 ,
    \sr[4]_i_127_1 ,
    \rgf_c0bus_wb_reg[7]_2 ,
    \rgf_c0bus_wb[14]_i_5_0 ,
    \rgf_c0bus_wb[5]_i_2_1 ,
    \rgf_c0bus_wb_reg[8]_1 ,
    \rgf_c0bus_wb_reg[8]_2 ,
    \rgf_c0bus_wb_reg[8]_3 ,
    \rgf_c0bus_wb_reg[8]_4 ,
    \rgf_c0bus_wb[4]_i_2_0 ,
    \rgf_c0bus_wb[4]_i_2_1 ,
    \sr[4]_i_128 ,
    \sr[4]_i_128_0 ,
    \rgf_c0bus_wb_reg[13]_0 ,
    p_1_in3_in,
    p_0_in2_in,
    \rgf_c0bus_wb_reg[13]_1 ,
    \sr[3]_i_3 ,
    .bbus_o_3_sp_1(bbus_o_3_sn_1),
    \bbus_o[3]_0 ,
    \rgf_c0bus_wb_reg[2]_1 ,
    .bbus_o_2_sp_1(bbus_o_2_sn_1),
    \bbus_o[2]_0 ,
    \rgf_c0bus_wb_reg[1]_0 ,
    .bbus_o_1_sp_1(bbus_o_1_sn_1),
    \bbus_o[1]_0 ,
    \rgf_c0bus_wb[4]_i_6_0 ,
    \rgf_c0bus_wb[4]_i_6_1 ,
    p_0_in,
    p_1_in,
    .bbus_o_0_sp_1(bbus_o_0_sn_1),
    \bbus_o[0]_0 ,
    \rgf_c0bus_wb[4]_i_5_0 ,
    \rgf_c0bus_wb_reg[5]_0 ,
    \rgf_c0bus_wb_reg[9]_2 ,
    \sr[4]_i_20_0 ,
    \rgf_selc0_rn_wb_reg[0] ,
    \rgf_selc0_rn_wb_reg[0]_0 ,
    ctl_fetch0_fl_reg_0,
    \stat_reg[0]_49 ,
    \stat_reg[0]_50 ,
    \stat[0]_i_8_0 ,
    \stat[0]_i_15_0 ,
    crdy,
    .ccmd_4_sp_1(ccmd_4_sn_1),
    \rgf_selc0_wb[1]_i_4_0 ,
    \ccmd[0]_INST_0_i_1_0 ,
    \ccmd[0]_INST_0_i_1_1 ,
    \stat_reg[0]_51 ,
    \fch_irq_lev[1]_i_2_0 ,
    irq_vec,
    brdy,
    ctl_fetch0_fl_reg_1,
    ctl_fetch0_fl_reg_2,
    \stat_reg[1]_8 ,
    \rgf_selc0_rn_wb_reg[0]_1 ,
    \rgf_selc0_wb[1]_i_4_1 ,
    \bdatw[15]_INST_0_i_67_0 ,
    \bcmd[1] ,
    \bcmd[1]_0 ,
    \sp[15]_i_8_0 ,
    \rgf_selc1_wb_reg[1] ,
    \stat[0]_i_2__1_0 ,
    \bbus_o[4]_INST_0_i_49_0 ,
    ctl_fetch1_fl_reg_i_6,
    \rgf_selc1_wb[1]_i_5_0 ,
    \read_cyc_reg[1] ,
    \rgf_selc1_wb_reg[1]_0 ,
    \sr[4]_i_3_0 ,
    \badr[15]_INST_0_i_25_0 ,
    \rgf_c1bus_wb[14]_i_53_0 ,
    \rgf_selc1_wb_reg[0] ,
    \ccmd[2]_INST_0_i_2_0 ,
    \badr[15]_INST_0_i_114_0 ,
    ctl_fetch1_fl_i_16,
    \rgf_selc0_rn_wb[0]_i_5_0 ,
    \stat_reg[0]_52 ,
    \read_cyc_reg[1]_0 ,
    \ccmd[2]_INST_0_i_3_0 ,
    ctl_fetch0_fl_i_8,
    \stat[0]_i_30_0 ,
    \ccmd[0]_INST_0_i_1_2 ,
    \stat_reg[2]_21 ,
    ctl_fetch0_fl_i_16,
    ctl_fetch0_fl_i_16_0,
    \stat_reg[0]_53 ,
    \ccmd[3]_INST_0_i_3_0 ,
    tout__1_carry_i_22_0,
    \rgf_selc1_rn_wb_reg[0] ,
    \rgf_selc1_rn_wb[1]_i_2_0 ,
    \rgf_selc1_rn_wb[1]_i_2_1 ,
    \stat_reg[0]_54 ,
    \rgf_selc1_rn_wb_reg[2] ,
    \stat_reg[0]_55 ,
    \badr[15]_INST_0_i_28_0 ,
    \iv_reg[15]_0 ,
    \stat[2]_i_2__1 ,
    \rgf_c1bus_wb[0]_i_16_0 ,
    \sr[15]_i_2 ,
    tout__1_carry_i_25_0,
    \rgf_selc1_wb[1]_i_5_1 ,
    \rgf_selc1_wb[1]_i_5_2 ,
    \stat_reg[0]_56 ,
    \ir1_id_fl_reg[20]_0 ,
    \nir_id_reg[21]_0 ,
    \ir1_id_fl_reg[21]_0 ,
    fdat,
    fdatx,
    fch_issu1_inferred_i_49_0,
    \nir_id_reg[24]_0 ,
    \rgf_c1bus_wb[4]_i_11_0 ,
    a1bus_b02,
    \rgf_c1bus_wb[4]_i_11_1 ,
    \rgf_c1bus_wb[4]_i_11_2 ,
    \sr[4]_i_18_3 ,
    \sr[4]_i_63_0 ,
    \sr[4]_i_63_1 ,
    \sr[4]_i_54_0 ,
    \sr[4]_i_54_1 ,
    \rgf_c0bus_wb[15]_i_4_0 ,
    \rgf_c0bus_wb_reg[5]_1 ,
    \rgf_c0bus_wb[11]_i_4_0 ,
    \rgf_c0bus_wb[2]_i_2_0 ,
    \rgf_c0bus_wb_reg[7]_3 ,
    \i_/rgf_c1bus_wb[4]_i_87 ,
    bank_sel,
    \i_/bdatw[12]_INST_0_i_64 ,
    \i_/bbus_o[4]_INST_0_i_22 ,
    \i_/bbus_o[4]_INST_0_i_22_0 ,
    \i_/bbus_o[4]_INST_0_i_23 ,
    \i_/bbus_o[4]_INST_0_i_23_0 ,
    \i_/bbus_o[0]_INST_0_i_18 ,
    \i_/bbus_o[4]_INST_0_i_20 ,
    \i_/bbus_o[4]_INST_0_i_21 ,
    \i_/bbus_o[4]_INST_0_i_21_0 ,
    \i_/bbus_o[4]_INST_0_i_20_0 ,
    \i_/rgf_c1bus_wb[4]_i_86 ,
    \i_/rgf_c1bus_wb[4]_i_96 ,
    \tr_reg[15]_1 ,
    cpuid,
    \rgf_c1bus_wb_reg[3]_3 ,
    \rgf_c1bus_wb_reg[0]_0 ,
    \rgf_c1bus_wb[0]_i_4_1 ,
    \rgf_c1bus_wb[1]_i_2_1 ,
    \rgf_c1bus_wb_reg[8]_1 ,
    \sr[6]_i_9_0 ,
    \sr[6]_i_6_2 ,
    \rgf_c1bus_wb_reg[8]_2 ,
    \sr[6]_i_9_1 ,
    \sr[6]_i_6_3 ,
    \rgf_c1bus_wb_reg[1]_1 ,
    \rgf_c1bus_wb_reg[13]_6 ,
    \rgf_c0bus_wb[12]_i_2_0 ,
    \rgf_c0bus_wb[13]_i_4_0 ,
    \rgf_c0bus_wb[15]_i_4_1 ,
    \rgf_c0bus_wb[15]_i_4_2 ,
    \sr[6]_i_5_0 ,
    SR,
    irq_lev);
  output [12:0]fadr;
  output fch_irq_req_fl;
  output fch_term;
  output [2:0]O;
  output [2:0]\pc_reg[15] ;
  output ctl_bcc_take0_fl;
  output ctl_bcc_take1_fl;
  output [15:0]\bdatr[15] ;
  output [15:0]\cbus_i[15] ;
  output p_2_in;
  output rst_n_fl_reg_1;
  output [2:0]\stat_reg[2] ;
  output [1:0]\stat_reg[2]_0 ;
  output [2:0]\stat_reg[2]_1 ;
  output [1:0]\stat_reg[2]_2 ;
  output [15:0]\sr_reg[15] ;
  output \stat_reg[2]_3 ;
  output tout__1_carry_i_11_0;
  output \tr_reg[4] ;
  output rst_n_0;
  output [14:0]b1bus_sr;
  output [5:0]b1bus_sel_cr;
  output [15:0]rgf_selc1_stat_reg;
  output \stat[2]_i_4 ;
  output \stat_reg[0] ;
  output \stat_reg[1] ;
  output [15:0]\sp_reg[15] ;
  output \stat_reg[0]_0 ;
  output \stat_reg[0]_1 ;
  output fch_leir_nir_reg;
  output \stat_reg[1]_0 ;
  output \stat_reg[2]_4 ;
  output [13:0]bdatw;
  output \bcmd[2]_INST_0_0 ;
  output \bcmd[1]_INST_0_0 ;
  output \tr_reg[4]_0 ;
  output \rgf_c1bus_wb[15]_i_14_0 ;
  output \stat_reg[2]_5 ;
  output \stat_reg[2]_6 ;
  output \stat_reg[2]_7 ;
  output \bdatw[8]_INST_0_i_16_0 ;
  output \bdatw[9]_INST_0_i_16_0 ;
  output \stat_reg[2]_8 ;
  output \bdatw[8]_INST_0_i_16_1 ;
  output \sr_reg[6] ;
  output \tr_reg[0] ;
  output \bdatw[8]_INST_0_i_16_2 ;
  output \rgf_c1bus_wb[15]_i_14_1 ;
  output \badr[14]_INST_0_i_1 ;
  output \bdatw[11]_INST_0_i_16_0 ;
  output \stat_reg[2]_9 ;
  output \tr_reg[0]_0 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[2]_10 ;
  output \stat_reg[1]_1 ;
  output [14:0]bbus_o;
  output \stat_reg[0]_3 ;
  output \rgf_c0bus_wb[15]_i_7_0 ;
  output \stat_reg[1]_2 ;
  output \bbus_o[2]_INST_0_i_1_0 ;
  output \bbus_o[3]_INST_0_i_1_0 ;
  output \bbus_o[1]_INST_0_i_1_0 ;
  output \rgf_c0bus_wb[11]_i_11_0 ;
  output \rgf_c0bus_wb[11]_i_3_0 ;
  output \rgf_c0bus_wb[13]_i_10_0 ;
  output \badr[15]_INST_0_i_2 ;
  output \badr[1]_INST_0_i_2 ;
  output \bbus_o[0]_INST_0_i_1_0 ;
  output \sr_reg[6]_0 ;
  output \bbus_o[1]_INST_0_i_1_1 ;
  output \bbus_o[1]_INST_0_i_1_2 ;
  output \tr_reg[0]_1 ;
  output [1:0]ctl_sela0_rn;
  output [2:0]\stat_reg[0]_4 ;
  output \stat_reg[2]_11 ;
  output [4:0]ccmd;
  output \stat_reg[0]_5 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[0]_6 ;
  output \sr_reg[5] ;
  output [0:0]ctl_selb0_0;
  output \stat_reg[0]_7 ;
  output \stat_reg[0]_8 ;
  output \stat_reg[0]_9 ;
  output \stat_reg[0]_10 ;
  output \stat_reg[1]_4 ;
  output rst_n_fl_reg_2;
  output [1:0]ctl_selb0_rn;
  output [2:0]\stat_reg[1]_5 ;
  output rst_n_fl_reg_3;
  output \stat_reg[0]_11 ;
  output [0:0]ctl_selb1_0;
  output \stat_reg[0]_12 ;
  output rst_n_fl_reg_4;
  output rst_n_fl_reg_5;
  output rst_n_fl_reg_6;
  output \stat_reg[0]_13 ;
  output \stat_reg[0]_14 ;
  output fch_leir_nir_reg_0;
  output rst_n_fl_reg_7;
  output rst_n_fl_reg_8;
  output fch_leir_nir_reg_1;
  output fch_leir_nir_reg_2;
  output fch_leir_nir_reg_3;
  output fch_leir_nir_reg_4;
  output fch_leir_nir_reg_5;
  output fch_leir_nir_reg_6;
  output fch_leir_nir_reg_7;
  output rst_n_fl_reg_9;
  output \stat_reg[1]_6 ;
  output [0:0]\stat_reg[0]_15 ;
  output [0:0]ctl_sela0;
  output [1:0]\stat_reg[2]_12 ;
  output \sr_reg[4] ;
  output [2:0]ctl_selb1_rn;
  output \stat_reg[0]_16 ;
  output \stat_reg[0]_17 ;
  output \stat_reg[0]_18 ;
  output [0:0]ir0_id;
  output fch_memacc1;
  output \stat_reg[1]_7 ;
  output \sr_reg[4]_0 ;
  output \stat_reg[2]_13 ;
  output [15:0]abus_o;
  output \sr_reg[0] ;
  output \stat_reg[0]_19 ;
  output \sr_reg[0]_0 ;
  output \sr_reg[0]_1 ;
  output \sr_reg[0]_2 ;
  output \sr_reg[0]_3 ;
  output \grn_reg[4] ;
  output \stat_reg[0]_20 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \sr_reg[0]_4 ;
  output \stat_reg[2]_14 ;
  output \stat_reg[2]_15 ;
  output \stat_reg[2]_16 ;
  output \sr_reg[0]_5 ;
  output \sr_reg[0]_6 ;
  output \sr_reg[0]_7 ;
  output \sr_reg[0]_8 ;
  output \sr_reg[0]_9 ;
  output \sr_reg[0]_10 ;
  output \sr_reg[0]_11 ;
  output \sr_reg[0]_12 ;
  output \sr_reg[0]_13 ;
  output \sr_reg[0]_14 ;
  output \sr_reg[0]_15 ;
  output \sr_reg[0]_16 ;
  output \sr_reg[0]_17 ;
  output \sr_reg[0]_18 ;
  output \sr_reg[0]_19 ;
  output \grn_reg[4]_0 ;
  output \stat_reg[0]_21 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \stat_reg[2]_17 ;
  output \stat_reg[0]_22 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[4]_2 ;
  output \stat_reg[0]_23 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_6 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_7 ;
  output \sr_reg[0]_20 ;
  output \sr_reg[0]_21 ;
  output \sr_reg[0]_22 ;
  output \sr_reg[0]_23 ;
  output \sr_reg[0]_24 ;
  output \sr_reg[0]_25 ;
  output \sr_reg[0]_26 ;
  output \sr_reg[0]_27 ;
  output \sr_reg[0]_28 ;
  output \sr_reg[0]_29 ;
  output \sr_reg[0]_30 ;
  output \sr_reg[0]_31 ;
  output \sr_reg[0]_32 ;
  output \sr_reg[0]_33 ;
  output \sr_reg[0]_34 ;
  output \sr_reg[0]_35 ;
  output \sr_reg[1] ;
  output \sr_reg[1]_0 ;
  output \sr_reg[1]_1 ;
  output \sr_reg[1]_2 ;
  output \sr_reg[1]_3 ;
  output \sr_reg[1]_4 ;
  output \sr_reg[1]_5 ;
  output \sr_reg[1]_6 ;
  output \sr_reg[1]_7 ;
  output \sr_reg[1]_8 ;
  output \sr_reg[1]_9 ;
  output \sr_reg[1]_10 ;
  output \sr_reg[1]_11 ;
  output \sr_reg[1]_12 ;
  output \sr_reg[1]_13 ;
  output \stat_reg[2]_18 ;
  output [0:0]E;
  output \stat_reg[0]_24 ;
  output \stat_reg[0]_25 ;
  output \stat_reg[0]_26 ;
  output \stat_reg[0]_27 ;
  output \stat_reg[0]_28 ;
  output \stat_reg[0]_29 ;
  output \stat_reg[0]_30 ;
  output \stat_reg[0]_31 ;
  output \stat_reg[0]_32 ;
  output rst_n_fl_reg_10;
  output rst_n_fl_reg_11;
  output rst_n_fl_reg_12;
  output \stat_reg[0]_33 ;
  output [0:0]\stat_reg[2]_19 ;
  output \stat_reg[2]_20 ;
  output fch_irq_req_fl_reg_0;
  output [3:0]a0bus_sel_cr;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4]_1 ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \tr_reg[15] ;
  output [15:0]b0bus_sr;
  output [0:0]\sr_reg[1]_14 ;
  output [0:0]\sr_reg[0]_36 ;
  output [0:0]\sr_reg[0]_37 ;
  output [0:0]\sr_reg[0]_38 ;
  output [0:0]\sr_reg[1]_15 ;
  output [0:0]\sr_reg[0]_39 ;
  output [0:0]\sr_reg[0]_40 ;
  output [0:0]\sr_reg[0]_41 ;
  output [0:0]\sr_reg[1]_16 ;
  output [0:0]\sr_reg[0]_42 ;
  output [0:0]\sr_reg[0]_43 ;
  output [0:0]\sr_reg[0]_44 ;
  output [0:0]\sr_reg[1]_17 ;
  output [0:0]\sr_reg[0]_45 ;
  output [0:0]\sr_reg[0]_46 ;
  output [0:0]\sr_reg[0]_47 ;
  output [0:0]\sr_reg[1]_18 ;
  output [0:0]\sr_reg[0]_48 ;
  output [0:0]\sr_reg[0]_49 ;
  output [0:0]\sr_reg[0]_50 ;
  output [0:0]\sr_reg[1]_19 ;
  output [0:0]\sr_reg[0]_51 ;
  output [0:0]\sr_reg[0]_52 ;
  output [0:0]\sr_reg[0]_53 ;
  output \rgf_c0bus_wb[15]_i_8_0 ;
  output \stat_reg[0]_34 ;
  output \stat_reg[0]_35 ;
  output \stat_reg[0]_36 ;
  output \stat_reg[0]_37 ;
  output \stat_reg[0]_38 ;
  output \stat_reg[0]_39 ;
  output \stat_reg[0]_40 ;
  output \stat_reg[0]_41 ;
  output \stat_reg[0]_42 ;
  output \stat_reg[0]_43 ;
  output \stat_reg[0]_44 ;
  output [14:0]badr;
  output [3:0]tout__1_carry_i_1__0_0;
  output [2:0]DI;
  output [1:0]\badr[15]_INST_0_i_1 ;
  output [0:0]\badr[15]_INST_0_i_1_0 ;
  output [0:0]\badr[15]_INST_0_i_1_1 ;
  output [2:0]\badr[14]_INST_0_i_2 ;
  output [3:0]\badr[15]_INST_0_i_2_0 ;
  output [0:0]\badr[15]_INST_0_i_2_1 ;
  output [1:0]\badr[15]_INST_0_i_2_2 ;
  output [15:0]a1bus_sr;
  output [4:0]a1bus_sel_cr;
  output [0:0]\sr_reg[0]_54 ;
  output [0:0]\sr_reg[1]_20 ;
  output [0:0]\sr_reg[0]_55 ;
  output [0:0]\sr_reg[0]_56 ;
  output [2:0]\badr[2]_INST_0_i_2 ;
  output [3:0]tout__1_carry_i_1_0;
  output [3:0]\badr[6]_INST_0_i_2 ;
  output [3:0]tout__1_carry__0_i_1_0;
  output [3:0]\badr[10]_INST_0_i_2 ;
  output [3:0]tout__1_carry__1_i_1_0;
  output [1:0]\badr[4]_INST_0_i_1 ;
  output [1:0]tout__1_carry__0_i_3__0_0;
  output [15:0]\pc0_reg[15]_0 ;
  output [15:0]\pc1_reg[15]_0 ;
  output [4:0]b0bus_sel_cr;
  output \stat_reg[0]_45 ;
  output [1:0]b0bus_sel_0;
  output \stat_reg[0]_46 ;
  output [3:0]a1bus_sel_0;
  output \stat_reg[0]_47 ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15]_0 ;
  output [3:0]a0bus_sel_0;
  output [15:0]rgf_selc1_stat_reg_0;
  output [15:0]rgf_selc1_stat_reg_1;
  output [15:0]rgf_selc1_stat_reg_2;
  output [15:0]rgf_selc1_stat_reg_3;
  output [15:0]rgf_selc1_stat_reg_4;
  output [15:0]rgf_selc1_stat_reg_5;
  output [15:0]rgf_selc1_stat_reg_6;
  output [15:0]rgf_selc1_stat_reg_7;
  output [15:0]rgf_selc1_stat_reg_8;
  output [15:0]rgf_selc1_stat_reg_9;
  output [15:0]rgf_selc1_stat_reg_10;
  output [15:0]rgf_selc1_stat_reg_11;
  output [15:0]rgf_selc1_stat_reg_12;
  output [15:0]rgf_selc1_stat_reg_13;
  output [15:0]rgf_selc1_stat_reg_14;
  output [15:0]rgf_selc1_stat_reg_15;
  output [15:0]rgf_selc1_stat_reg_16;
  output [15:0]rgf_selc1_stat_reg_17;
  output [15:0]rgf_selc1_stat_reg_18;
  output [15:0]rgf_selc1_stat_reg_19;
  output [15:0]rgf_selc1_stat_reg_20;
  output [15:0]rgf_selc1_stat_reg_21;
  output [15:0]rgf_selc1_stat_reg_22;
  output [15:0]rgf_selc1_stat_reg_23;
  output [15:0]rgf_selc1_stat_reg_24;
  output [15:0]rgf_selc1_stat_reg_25;
  output [15:0]rgf_selc1_stat_reg_26;
  output [15:0]rgf_selc1_stat_reg_27;
  output [15:0]rgf_selc1_stat_reg_28;
  output [15:0]rgf_selc1_stat_reg_29;
  output [15:0]rgf_selc1_stat_reg_30;
  output [15:0]rgf_selc1_stat_reg_31;
  output [0:0]\sr_reg[0]_57 ;
  output [0:0]\sr_reg[0]_58 ;
  output [0:0]\sr_reg[0]_59 ;
  output [0:0]\sr_reg[1]_21 ;
  input rst_n;
  input clk;
  input fch_irq_req;
  input [15:0]\pc0_reg[15]_1 ;
  input [0:0]S;
  input [0:0]\fadr[3] ;
  input [2:0]D;
  input [2:0]\pc1_reg[15]_1 ;
  input ctl_bcc_take0_fl_reg_0;
  input ctl_bcc_take1_fl_reg_0;
  input \grn_reg[15] ;
  input rgf_selc1_stat;
  input [15:0]Q;
  input rgf_selc0_stat;
  input [15:0]\pc_reg[15]_0 ;
  input [2:0]\grn_reg[15]_0 ;
  input [1:0]\grn[15]_i_3__5 ;
  input [2:0]\sr[13]_i_5 ;
  input [1:0]\sr[13]_i_5_0 ;
  input \sr_reg[4]_1 ;
  input \sr_reg[5]_0 ;
  input [15:0]\sr_reg[15]_0 ;
  input [0:0]\sr_reg[6]_1 ;
  input \pc_reg[15]_1 ;
  input \pc_reg[14] ;
  input \pc_reg[13] ;
  input \sp_reg[15]_0 ;
  input \sp_reg[14] ;
  input \sp_reg[13] ;
  input \sp_reg[12] ;
  input \sp_reg[11] ;
  input \sp_reg[10] ;
  input \sp_reg[9] ;
  input \sp_reg[8] ;
  input \sp_reg[7] ;
  input \sp_reg[6] ;
  input \sp_reg[5] ;
  input \sp_reg[1] ;
  input \sp_reg[3] ;
  input \sp_reg[4] ;
  input \sp_reg[2] ;
  input [0:0]\sp_reg[0] ;
  input [0:0]\sp_reg[0]_0 ;
  input \sp[15]_i_2 ;
  input [1:0]\rgf_c1bus_wb_reg[15] ;
  input \rgf_c1bus_wb_reg[15]_0 ;
  input [15:0]a1bus_0;
  input \bdatw[15] ;
  input \stat_reg[0]_48 ;
  input \bdatw[15]_0 ;
  input \bdatw[15]_1 ;
  input \bdatw[15]_2 ;
  input \rgf_c1bus_wb_reg[14] ;
  input \rgf_c1bus_wb_reg[14]_0 ;
  input \rgf_c1bus_wb[14]_i_3_0 ;
  input \rgf_c1bus_wb_reg[13] ;
  input \rgf_c1bus_wb[13]_i_5_0 ;
  input [4:0]bdatr;
  input \rgf_c1bus_wb_reg[12] ;
  input \bdatw[12]_0 ;
  input [1:0]\rgf_c1bus_wb_reg[11] ;
  input \bdatw[11]_0 ;
  input \rgf_c1bus_wb_reg[10] ;
  input \sr[4]_i_52_0 ;
  input \bdatw[10]_0 ;
  input \rgf_c1bus_wb_reg[9] ;
  input \bdatw[9]_0 ;
  input \rgf_c1bus_wb_reg[8] ;
  input \bdatw[8]_0 ;
  input \rgf_c1bus_wb[15]_i_10_0 ;
  input \rgf_c1bus_wb_reg[7] ;
  input \rgf_c1bus_wb_reg[7]_0 ;
  input [2:0]\rgf_c1bus_wb_reg[7]_1 ;
  input \rgf_c1bus_wb_reg[6] ;
  input \rgf_c1bus_wb_reg[6]_0 ;
  input \rgf_c1bus_wb_reg[6]_1 ;
  input \rgf_c1bus_wb[14]_i_3_1 ;
  input \rgf_c1bus_wb_reg[5] ;
  input \rgf_c1bus_wb_reg[5]_0 ;
  input \sr[4]_i_53_0 ;
  input \sr[4]_i_53_1 ;
  input tout__1_carry__0;
  input \sr[4]_i_10_0 ;
  input \rgf_c1bus_wb_reg[13]_0 ;
  input \rgf_c1bus_wb_reg[1] ;
  input \rgf_c1bus_wb[9]_i_3_0 ;
  input \rgf_c1bus_wb[9]_i_3_1 ;
  input \sr[4]_i_9_0 ;
  input \rgf_c1bus_wb_reg[15]_1 ;
  input \sr[4]_i_41_0 ;
  input \rgf_c1bus_wb_reg[3] ;
  input \sr[4]_i_35_0 ;
  input \rgf_c1bus_wb_reg[3]_0 ;
  input \rgf_c1bus_wb_reg[3]_1 ;
  input \sr[4]_i_91 ;
  input \sr[4]_i_100_0 ;
  input \sr[4]_i_10_1 ;
  input \sr[4]_i_10_2 ;
  input \rgf_c1bus_wb_reg[7]_2 ;
  input \rgf_c1bus_wb_reg[11]_0 ;
  input \sr[4]_i_35_1 ;
  input \rgf_c1bus_wb[11]_i_6_0 ;
  input \sr[4]_i_98_0 ;
  input \sr[4]_i_98_1 ;
  input \sr[4]_i_30_0 ;
  input \sr[4]_i_30_1 ;
  input \rgf_c1bus_wb_reg[8]_0 ;
  input \rgf_c1bus_wb_reg[12]_0 ;
  input \rgf_c1bus_wb_reg[4] ;
  input \sr[4]_i_11_0 ;
  input \rgf_c1bus_wb_reg[4]_0 ;
  input \sr[6]_i_6_0 ;
  input \rgf_c1bus_wb[4]_i_4_0 ;
  input \rgf_c1bus_wb[4]_i_4_1 ;
  input \rgf_c1bus_wb_reg[0] ;
  input \sr[4]_i_36_0 ;
  input \sr[4]_i_25_0 ;
  input \rgf_c1bus_wb[4]_i_4_2 ;
  input \rgf_c1bus_wb[4]_i_4_3 ;
  input \rgf_c1bus_wb_reg[12]_1 ;
  input \sr[4]_i_111_0 ;
  input \sr[4]_i_36_1 ;
  input \sr[4]_i_36_2 ;
  input \rgf_c1bus_wb_reg[4]_1 ;
  input \sr[6]_i_6_1 ;
  input \rgf_c1bus_wb_reg[13]_1 ;
  input \sr[4]_i_37_0 ;
  input \sr[4]_i_39_0 ;
  input \rgf_c1bus_wb[0]_i_4_0 ;
  input \sr[4]_i_29_0 ;
  input \rgf_c1bus_wb_reg[9]_0 ;
  input \rgf_c1bus_wb[13]_i_2_0 ;
  input \sr[4]_i_27_0 ;
  input \rgf_c1bus_wb_reg[13]_2 ;
  input \sr[4]_i_29_1 ;
  input \sr[4]_i_29_2 ;
  input \rgf_c1bus_wb[1]_i_2_0 ;
  input \rgf_c1bus_wb_reg[2] ;
  input \sr[4]_i_12_0 ;
  input \rgf_c1bus_wb_reg[14]_1 ;
  input \rgf_c1bus_wb_reg[14]_2 ;
  input \sr[4]_i_29_3 ;
  input \rgf_c1bus_wb_reg[10]_0 ;
  input \sr[4]_i_44_0 ;
  input \sr[4]_i_46_0 ;
  input \sr[4]_i_43_0 ;
  input \sr[4]_i_43_1 ;
  input \rgf_c1bus_wb_reg[6]_2 ;
  input \rgf_c1bus_wb_reg[6]_3 ;
  input \sr[4]_i_43_2 ;
  input \rgf_c1bus_wb_reg[14]_3 ;
  input \sr[4]_i_46_1 ;
  input \sr[4]_i_46_2 ;
  input \rgf_c1bus_wb_reg[2]_0 ;
  input \sr[4]_i_45_0 ;
  input \sr[4]_i_34_0 ;
  input \sr[4]_i_102_0 ;
  input \rgf_c1bus_wb[9]_i_3_2 ;
  input \rgf_c1bus_wb[15]_i_4_0 ;
  input \sr[4]_i_33_0 ;
  input \sr[4]_i_28_0 ;
  input \sr[4]_i_28_1 ;
  input \rgf_c1bus_wb_reg[7]_3 ;
  input \rgf_c1bus_wb[11]_i_3_0 ;
  input \sr[4]_i_100_1 ;
  input \sr[4]_i_100_2 ;
  input \rgf_c1bus_wb_reg[4]_2 ;
  input \rgf_c1bus_wb_reg[13]_3 ;
  input [4:0]b1bus_b02;
  input \rgf_c1bus_wb_reg[13]_4 ;
  input \rgf_c1bus_wb_reg[13]_5 ;
  input \sr[4]_i_102_1 ;
  input \sr[4]_i_102_2 ;
  input \sr[4]_i_102_3 ;
  input \rgf_c1bus_wb[5]_i_9_0 ;
  input \rgf_c1bus_wb[5]_i_9_1 ;
  input \rgf_c1bus_wb[5]_i_9_2 ;
  input \rgf_c1bus_wb_reg[1]_0 ;
  input [2:0]\rgf_c1bus_wb_reg[3]_2 ;
  input \rgf_c1bus_wb[14]_i_28_0 ;
  input \rgf_c1bus_wb[14]_i_28_1 ;
  input \rgf_c1bus_wb[14]_i_28_2 ;
  input \sr[6]_i_16 ;
  input \sr[6]_i_16_0 ;
  input \sr[6]_i_16_1 ;
  input [3:0]\rgf_c0bus_wb_reg[15] ;
  input \rgf_c0bus_wb_reg[15]_0 ;
  input [15:0]a0bus_0;
  input \rgf_c0bus_wb_reg[14] ;
  input \rgf_c0bus_wb_reg[12] ;
  input \rgf_c0bus_wb_reg[11] ;
  input [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  input \sr[4]_i_72_0 ;
  input \rgf_c0bus_wb_reg[10] ;
  input \rgf_c0bus_wb_reg[10]_0 ;
  input \rgf_c0bus_wb_reg[9] ;
  input \rgf_c0bus_wb_reg[8] ;
  input \sr[4]_i_71_0 ;
  input \rgf_c0bus_wb_reg[10]_i_17_0 ;
  input [9:0]cbus_i;
  input \rgf_c0bus_wb_reg[7] ;
  input [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  input \sr[4]_i_69_0 ;
  input \rgf_c0bus_wb_reg[10]_i_17_1 ;
  input \rgf_c0bus_wb_reg[10]_i_17_2 ;
  input \rgf_c0bus_wb_reg[6] ;
  input \sr[4]_i_70_0 ;
  input \rgf_c0bus_wb_reg[5] ;
  input \rgf_c0bus_wb_reg[10]_1 ;
  input \sr[4]_i_6_0 ;
  input \rgf_c0bus_wb_reg[7]_1 ;
  input \sr[6]_i_5 ;
  input \sr[4]_i_17_0 ;
  input [3:0]\rgf_c0bus_wb_reg[3] ;
  input \rgf_c0bus_wb_reg[0] ;
  input \rgf_c0bus_wb[0]_i_2_0 ;
  input \sr[4]_i_66_0 ;
  input \rgf_c0bus_wb[5]_i_2_0 ;
  input \rgf_c0bus_wb_reg[2] ;
  input \rgf_c0bus_wb_reg[2]_0 ;
  input \rgf_c0bus_wb_reg[3]_0 ;
  input \sr[4]_i_17_1 ;
  input \sr[4]_i_18_0 ;
  input \sr[4]_i_18_1 ;
  input \sr[4]_i_18_2 ;
  input \sr[4]_i_15_0 ;
  input \rgf_c0bus_wb_reg[11]_1 ;
  input \sr[4]_i_55_0 ;
  input \rgf_c0bus_wb_reg[11]_2 ;
  input \rgf_c0bus_wb_reg[11]_3 ;
  input \rgf_c0bus_wb_reg[12]_0 ;
  input \rgf_c0bus_wb_reg[13] ;
  input \rgf_c0bus_wb_reg[14]_0 ;
  input \sr[4]_i_16_0 ;
  input \rgf_c0bus_wb[12]_i_3_0 ;
  input \rgf_c0bus_wb[13]_i_2_0 ;
  input \rgf_c0bus_wb_reg[4] ;
  input \rgf_c0bus_wb_reg[4]_0 ;
  input \rgf_c0bus_wb[12]_i_3_1 ;
  input \rgf_c0bus_wb_reg[1] ;
  input \rgf_c0bus_wb[5]_i_3_0 ;
  input \sr[4]_i_67_0 ;
  input \rgf_c0bus_wb_reg[8]_0 ;
  input \rgf_c0bus_wb[1]_i_3_0 ;
  input \rgf_c0bus_wb[9]_i_3_0 ;
  input \rgf_c0bus_wb[10]_i_4_0 ;
  input \rgf_c0bus_wb[10]_i_4_1 ;
  input \rgf_c0bus_wb[11]_i_5_0 ;
  input \rgf_c0bus_wb[13]_i_2_1 ;
  input \rgf_c0bus_wb[13]_i_2_2 ;
  input \sr[4]_i_58_0 ;
  input \sr[4]_i_55_1 ;
  input \sr[4]_i_55_2 ;
  input \sr[4]_i_60_0 ;
  input \sr[4]_i_65_0 ;
  input \sr[4]_i_68_0 ;
  input \rgf_c0bus_wb[9]_i_3_1 ;
  input \rgf_c0bus_wb[5]_i_3_1 ;
  input \rgf_c0bus_wb_reg[6]_0 ;
  input \rgf_c0bus_wb_reg[6]_1 ;
  input \rgf_c0bus_wb_reg[4]_1 ;
  input \rgf_c0bus_wb_reg[4]_2 ;
  input \rgf_c0bus_wb_reg[9]_0 ;
  input \rgf_c0bus_wb_reg[9]_1 ;
  input \rgf_c0bus_wb_reg[10]_2 ;
  input \sr[4]_i_64_0 ;
  input \sr[4]_i_60_1 ;
  input \rgf_c0bus_wb_reg[10]_3 ;
  input \rgf_c0bus_wb[4]_i_3_0 ;
  input \rgf_c0bus_wb[4]_i_3_1 ;
  input \rgf_c0bus_wb[5]_i_3_2 ;
  input \sr[4]_i_68_1 ;
  input \rgf_c0bus_wb[0]_i_2_1 ;
  input \sr[4]_i_64_1 ;
  input \sr[4]_i_60_2 ;
  input \sr[4]_i_127_0 ;
  input \sr[4]_i_127_1 ;
  input \rgf_c0bus_wb_reg[7]_2 ;
  input \rgf_c0bus_wb[14]_i_5_0 ;
  input \rgf_c0bus_wb[5]_i_2_1 ;
  input \rgf_c0bus_wb_reg[8]_1 ;
  input \rgf_c0bus_wb_reg[8]_2 ;
  input \rgf_c0bus_wb_reg[8]_3 ;
  input \rgf_c0bus_wb_reg[8]_4 ;
  input \rgf_c0bus_wb[4]_i_2_0 ;
  input \rgf_c0bus_wb[4]_i_2_1 ;
  input \sr[4]_i_128 ;
  input \sr[4]_i_128_0 ;
  input \rgf_c0bus_wb_reg[13]_0 ;
  input [4:0]p_1_in3_in;
  input [4:0]p_0_in2_in;
  input \rgf_c0bus_wb_reg[13]_1 ;
  input \sr[3]_i_3 ;
  input \bbus_o[3]_0 ;
  input \rgf_c0bus_wb_reg[2]_1 ;
  input \bbus_o[2]_0 ;
  input \rgf_c0bus_wb_reg[1]_0 ;
  input \bbus_o[1]_0 ;
  input \rgf_c0bus_wb[4]_i_6_0 ;
  input \rgf_c0bus_wb[4]_i_6_1 ;
  input [0:0]p_0_in;
  input [0:0]p_1_in;
  input \bbus_o[0]_0 ;
  input \rgf_c0bus_wb[4]_i_5_0 ;
  input \rgf_c0bus_wb_reg[5]_0 ;
  input \rgf_c0bus_wb_reg[9]_2 ;
  input \sr[4]_i_20_0 ;
  input [2:0]\rgf_selc0_rn_wb_reg[0] ;
  input \rgf_selc0_rn_wb_reg[0]_0 ;
  input ctl_fetch0_fl_reg_0;
  input \stat_reg[0]_49 ;
  input \stat_reg[0]_50 ;
  input \stat[0]_i_8_0 ;
  input \stat[0]_i_15_0 ;
  input crdy;
  input \rgf_selc0_wb[1]_i_4_0 ;
  input \ccmd[0]_INST_0_i_1_0 ;
  input \ccmd[0]_INST_0_i_1_1 ;
  input \stat_reg[0]_51 ;
  input \fch_irq_lev[1]_i_2_0 ;
  input [5:0]irq_vec;
  input brdy;
  input ctl_fetch0_fl_reg_1;
  input ctl_fetch0_fl_reg_2;
  input \stat_reg[1]_8 ;
  input \rgf_selc0_rn_wb_reg[0]_1 ;
  input \rgf_selc0_wb[1]_i_4_1 ;
  input \bdatw[15]_INST_0_i_67_0 ;
  input \bcmd[1] ;
  input \bcmd[1]_0 ;
  input \sp[15]_i_8_0 ;
  input [2:0]\rgf_selc1_wb_reg[1] ;
  input \stat[0]_i_2__1_0 ;
  input \bbus_o[4]_INST_0_i_49_0 ;
  input ctl_fetch1_fl_reg_i_6;
  input \rgf_selc1_wb[1]_i_5_0 ;
  input \read_cyc_reg[1] ;
  input \rgf_selc1_wb_reg[1]_0 ;
  input \sr[4]_i_3_0 ;
  input \badr[15]_INST_0_i_25_0 ;
  input \rgf_c1bus_wb[14]_i_53_0 ;
  input \rgf_selc1_wb_reg[0] ;
  input \ccmd[2]_INST_0_i_2_0 ;
  input \badr[15]_INST_0_i_114_0 ;
  input ctl_fetch1_fl_i_16;
  input \rgf_selc0_rn_wb[0]_i_5_0 ;
  input \stat_reg[0]_52 ;
  input \read_cyc_reg[1]_0 ;
  input \ccmd[2]_INST_0_i_3_0 ;
  input ctl_fetch0_fl_i_8;
  input \stat[0]_i_30_0 ;
  input \ccmd[0]_INST_0_i_1_2 ;
  input \stat_reg[2]_21 ;
  input ctl_fetch0_fl_i_16;
  input ctl_fetch0_fl_i_16_0;
  input \stat_reg[0]_53 ;
  input \ccmd[3]_INST_0_i_3_0 ;
  input tout__1_carry_i_22_0;
  input \rgf_selc1_rn_wb_reg[0] ;
  input \rgf_selc1_rn_wb[1]_i_2_0 ;
  input \rgf_selc1_rn_wb[1]_i_2_1 ;
  input \stat_reg[0]_54 ;
  input \rgf_selc1_rn_wb_reg[2] ;
  input \stat_reg[0]_55 ;
  input \badr[15]_INST_0_i_28_0 ;
  input [15:0]\iv_reg[15]_0 ;
  input \stat[2]_i_2__1 ;
  input \rgf_c1bus_wb[0]_i_16_0 ;
  input \sr[15]_i_2 ;
  input tout__1_carry_i_25_0;
  input \rgf_selc1_wb[1]_i_5_1 ;
  input \rgf_selc1_wb[1]_i_5_2 ;
  input [1:0]\stat_reg[0]_56 ;
  input \ir1_id_fl_reg[20]_0 ;
  input [1:0]\nir_id_reg[21]_0 ;
  input \ir1_id_fl_reg[21]_0 ;
  input [15:0]fdat;
  input [15:0]fdatx;
  input fch_issu1_inferred_i_49_0;
  input \nir_id_reg[24]_0 ;
  input \rgf_c1bus_wb[4]_i_11_0 ;
  input [0:0]a1bus_b02;
  input \rgf_c1bus_wb[4]_i_11_1 ;
  input \rgf_c1bus_wb[4]_i_11_2 ;
  input \sr[4]_i_18_3 ;
  input \sr[4]_i_63_0 ;
  input \sr[4]_i_63_1 ;
  input \sr[4]_i_54_0 ;
  input \sr[4]_i_54_1 ;
  input \rgf_c0bus_wb[15]_i_4_0 ;
  input \rgf_c0bus_wb_reg[5]_1 ;
  input \rgf_c0bus_wb[11]_i_4_0 ;
  input \rgf_c0bus_wb[2]_i_2_0 ;
  input \rgf_c0bus_wb_reg[7]_3 ;
  input [15:0]\i_/rgf_c1bus_wb[4]_i_87 ;
  input [0:0]bank_sel;
  input [4:0]\i_/bdatw[12]_INST_0_i_64 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_22 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_22_0 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_23 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_23_0 ;
  input \i_/bbus_o[0]_INST_0_i_18 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_20 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_21 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_21_0 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_20_0 ;
  input [15:0]\i_/rgf_c1bus_wb[4]_i_86 ;
  input [14:0]\i_/rgf_c1bus_wb[4]_i_96 ;
  input [15:0]\tr_reg[15]_1 ;
  input [1:0]cpuid;
  input \rgf_c1bus_wb_reg[3]_3 ;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input \rgf_c1bus_wb[0]_i_4_1 ;
  input \rgf_c1bus_wb[1]_i_2_1 ;
  input \rgf_c1bus_wb_reg[8]_1 ;
  input \sr[6]_i_9_0 ;
  input \sr[6]_i_6_2 ;
  input \rgf_c1bus_wb_reg[8]_2 ;
  input \sr[6]_i_9_1 ;
  input \sr[6]_i_6_3 ;
  input \rgf_c1bus_wb_reg[1]_1 ;
  input \rgf_c1bus_wb_reg[13]_6 ;
  input \rgf_c0bus_wb[12]_i_2_0 ;
  input \rgf_c0bus_wb[13]_i_4_0 ;
  input \rgf_c0bus_wb[15]_i_4_1 ;
  input \rgf_c0bus_wb[15]_i_4_2 ;
  input [0:0]\sr[6]_i_5_0 ;
  input [0:0]SR;
  input [1:0]irq_lev;
     output [15:0]ir0;
     output [15:0]ir1;
  output fdatx_5_sn_1;
  output fdatx_14_sn_1;
  output fdat_0_sn_1;
  output fdat_12_sn_1;
  output fdat_5_sn_1;
  input bdatw_12_sn_1;
  input bdatw_11_sn_1;
  input bdatw_10_sn_1;
  input bdatw_9_sn_1;
  input bdatw_8_sn_1;
  input bdatw_6_sn_1;
  input bdatw_5_sn_1;
  input bbus_o_14_sn_1;
  input bbus_o_13_sn_1;
  input bbus_o_7_sn_1;
  input bbus_o_6_sn_1;
  input bbus_o_3_sn_1;
  input bbus_o_2_sn_1;
  input bbus_o_1_sn_1;
  input bbus_o_0_sn_1;
  input ccmd_4_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]DI;
  wire [0:0]E;
  wire [2:0]O;
  wire [15:0]Q;
  wire [0:0]S;
  wire [0:0]SR;
  wire [15:0]a0bus_0;
  wire [3:0]a0bus_sel_0;
  wire [3:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [0:0]a1bus_b02;
  wire [3:0]a1bus_sel_0;
  wire [4:0]a1bus_sel_cr;
  wire [15:0]a1bus_sr;
  wire [15:0]abus_o;
  wire [3:0]alu_sr_flag0;
  wire [0:0]alu_sr_flag1;
  wire [1:0]b0bus_sel_0;
  wire [4:0]b0bus_sel_cr;
  wire [15:0]b0bus_sr;
  wire [4:0]b1bus_b02;
  wire [5:0]b1bus_sel_cr;
  wire [14:0]b1bus_sr;
  wire [14:0]badr;
  wire [3:0]\badr[10]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_1 ;
  wire [2:0]\badr[14]_INST_0_i_2 ;
  wire [1:0]\badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_109_n_0 ;
  wire \badr[15]_INST_0_i_110_n_0 ;
  wire \badr[15]_INST_0_i_111_n_0 ;
  wire \badr[15]_INST_0_i_112_n_0 ;
  wire \badr[15]_INST_0_i_114_0 ;
  wire \badr[15]_INST_0_i_139_n_0 ;
  wire \badr[15]_INST_0_i_140_n_0 ;
  wire \badr[15]_INST_0_i_142_n_0 ;
  wire \badr[15]_INST_0_i_143_n_0 ;
  wire \badr[15]_INST_0_i_144_n_0 ;
  wire \badr[15]_INST_0_i_146_n_0 ;
  wire \badr[15]_INST_0_i_147_n_0 ;
  wire \badr[15]_INST_0_i_148_n_0 ;
  wire \badr[15]_INST_0_i_149_n_0 ;
  wire \badr[15]_INST_0_i_150_n_0 ;
  wire \badr[15]_INST_0_i_151_n_0 ;
  wire \badr[15]_INST_0_i_152_n_0 ;
  wire \badr[15]_INST_0_i_153_n_0 ;
  wire \badr[15]_INST_0_i_154_n_0 ;
  wire \badr[15]_INST_0_i_155_n_0 ;
  wire \badr[15]_INST_0_i_156_n_0 ;
  wire \badr[15]_INST_0_i_157_n_0 ;
  wire \badr[15]_INST_0_i_158_n_0 ;
  wire \badr[15]_INST_0_i_159_n_0 ;
  wire \badr[15]_INST_0_i_160_n_0 ;
  wire \badr[15]_INST_0_i_161_n_0 ;
  wire \badr[15]_INST_0_i_162_n_0 ;
  wire \badr[15]_INST_0_i_163_n_0 ;
  wire \badr[15]_INST_0_i_164_n_0 ;
  wire \badr[15]_INST_0_i_165_n_0 ;
  wire \badr[15]_INST_0_i_166_n_0 ;
  wire \badr[15]_INST_0_i_167_n_0 ;
  wire \badr[15]_INST_0_i_168_n_0 ;
  wire \badr[15]_INST_0_i_169_n_0 ;
  wire \badr[15]_INST_0_i_170_n_0 ;
  wire \badr[15]_INST_0_i_171_n_0 ;
  wire \badr[15]_INST_0_i_173_n_0 ;
  wire \badr[15]_INST_0_i_174_n_0 ;
  wire \badr[15]_INST_0_i_175_n_0 ;
  wire \badr[15]_INST_0_i_176_n_0 ;
  wire \badr[15]_INST_0_i_177_n_0 ;
  wire \badr[15]_INST_0_i_178_n_0 ;
  wire \badr[15]_INST_0_i_179_n_0 ;
  wire \badr[15]_INST_0_i_180_n_0 ;
  wire \badr[15]_INST_0_i_181_n_0 ;
  wire \badr[15]_INST_0_i_182_n_0 ;
  wire \badr[15]_INST_0_i_183_n_0 ;
  wire \badr[15]_INST_0_i_184_n_0 ;
  wire \badr[15]_INST_0_i_187_n_0 ;
  wire \badr[15]_INST_0_i_188_n_0 ;
  wire \badr[15]_INST_0_i_189_n_0 ;
  wire \badr[15]_INST_0_i_190_n_0 ;
  wire \badr[15]_INST_0_i_191_n_0 ;
  wire \badr[15]_INST_0_i_192_n_0 ;
  wire \badr[15]_INST_0_i_193_n_0 ;
  wire \badr[15]_INST_0_i_194_n_0 ;
  wire \badr[15]_INST_0_i_195_n_0 ;
  wire \badr[15]_INST_0_i_196_n_0 ;
  wire \badr[15]_INST_0_i_197_n_0 ;
  wire \badr[15]_INST_0_i_198_n_0 ;
  wire \badr[15]_INST_0_i_199_n_0 ;
  wire [0:0]\badr[15]_INST_0_i_1_0 ;
  wire [0:0]\badr[15]_INST_0_i_1_1 ;
  wire \badr[15]_INST_0_i_2 ;
  wire \badr[15]_INST_0_i_200_n_0 ;
  wire \badr[15]_INST_0_i_201_n_0 ;
  wire \badr[15]_INST_0_i_202_n_0 ;
  wire \badr[15]_INST_0_i_203_n_0 ;
  wire \badr[15]_INST_0_i_204_n_0 ;
  wire \badr[15]_INST_0_i_205_n_0 ;
  wire \badr[15]_INST_0_i_206_n_0 ;
  wire \badr[15]_INST_0_i_207_n_0 ;
  wire \badr[15]_INST_0_i_208_n_0 ;
  wire \badr[15]_INST_0_i_209_n_0 ;
  wire \badr[15]_INST_0_i_224_n_0 ;
  wire \badr[15]_INST_0_i_225_n_0 ;
  wire \badr[15]_INST_0_i_226_n_0 ;
  wire \badr[15]_INST_0_i_227_n_0 ;
  wire \badr[15]_INST_0_i_229_n_0 ;
  wire \badr[15]_INST_0_i_230_n_0 ;
  wire \badr[15]_INST_0_i_231_n_0 ;
  wire \badr[15]_INST_0_i_232_n_0 ;
  wire \badr[15]_INST_0_i_233_n_0 ;
  wire \badr[15]_INST_0_i_234_n_0 ;
  wire \badr[15]_INST_0_i_235_n_0 ;
  wire \badr[15]_INST_0_i_236_n_0 ;
  wire \badr[15]_INST_0_i_237_n_0 ;
  wire \badr[15]_INST_0_i_238_n_0 ;
  wire \badr[15]_INST_0_i_239_n_0 ;
  wire \badr[15]_INST_0_i_240_n_0 ;
  wire \badr[15]_INST_0_i_241_n_0 ;
  wire \badr[15]_INST_0_i_242_n_0 ;
  wire \badr[15]_INST_0_i_243_n_0 ;
  wire \badr[15]_INST_0_i_244_n_0 ;
  wire \badr[15]_INST_0_i_245_n_0 ;
  wire \badr[15]_INST_0_i_246_n_0 ;
  wire \badr[15]_INST_0_i_247_n_0 ;
  wire \badr[15]_INST_0_i_248_n_0 ;
  wire \badr[15]_INST_0_i_249_n_0 ;
  wire \badr[15]_INST_0_i_250_n_0 ;
  wire \badr[15]_INST_0_i_251_n_0 ;
  wire \badr[15]_INST_0_i_252_n_0 ;
  wire \badr[15]_INST_0_i_253_n_0 ;
  wire \badr[15]_INST_0_i_254_n_0 ;
  wire \badr[15]_INST_0_i_255_n_0 ;
  wire \badr[15]_INST_0_i_256_n_0 ;
  wire \badr[15]_INST_0_i_257_n_0 ;
  wire \badr[15]_INST_0_i_258_n_0 ;
  wire \badr[15]_INST_0_i_259_n_0 ;
  wire \badr[15]_INST_0_i_25_0 ;
  wire \badr[15]_INST_0_i_25_n_0 ;
  wire \badr[15]_INST_0_i_260_n_0 ;
  wire \badr[15]_INST_0_i_261_n_0 ;
  wire \badr[15]_INST_0_i_262_n_0 ;
  wire \badr[15]_INST_0_i_263_n_0 ;
  wire \badr[15]_INST_0_i_264_n_0 ;
  wire \badr[15]_INST_0_i_265_n_0 ;
  wire \badr[15]_INST_0_i_266_n_0 ;
  wire \badr[15]_INST_0_i_267_n_0 ;
  wire \badr[15]_INST_0_i_268_n_0 ;
  wire \badr[15]_INST_0_i_269_n_0 ;
  wire \badr[15]_INST_0_i_26_n_0 ;
  wire \badr[15]_INST_0_i_270_n_0 ;
  wire \badr[15]_INST_0_i_271_n_0 ;
  wire \badr[15]_INST_0_i_272_n_0 ;
  wire \badr[15]_INST_0_i_273_n_0 ;
  wire \badr[15]_INST_0_i_274_n_0 ;
  wire \badr[15]_INST_0_i_275_n_0 ;
  wire \badr[15]_INST_0_i_276_n_0 ;
  wire \badr[15]_INST_0_i_277_n_0 ;
  wire \badr[15]_INST_0_i_278_n_0 ;
  wire \badr[15]_INST_0_i_279_n_0 ;
  wire \badr[15]_INST_0_i_280_n_0 ;
  wire \badr[15]_INST_0_i_281_n_0 ;
  wire \badr[15]_INST_0_i_282_n_0 ;
  wire \badr[15]_INST_0_i_283_n_0 ;
  wire \badr[15]_INST_0_i_284_n_0 ;
  wire \badr[15]_INST_0_i_285_n_0 ;
  wire \badr[15]_INST_0_i_286_n_0 ;
  wire \badr[15]_INST_0_i_287_n_0 ;
  wire \badr[15]_INST_0_i_288_n_0 ;
  wire \badr[15]_INST_0_i_289_n_0 ;
  wire \badr[15]_INST_0_i_28_0 ;
  wire \badr[15]_INST_0_i_290_n_0 ;
  wire \badr[15]_INST_0_i_291_n_0 ;
  wire \badr[15]_INST_0_i_292_n_0 ;
  wire \badr[15]_INST_0_i_293_n_0 ;
  wire \badr[15]_INST_0_i_294_n_0 ;
  wire \badr[15]_INST_0_i_296_n_0 ;
  wire \badr[15]_INST_0_i_297_n_0 ;
  wire \badr[15]_INST_0_i_298_n_0 ;
  wire \badr[15]_INST_0_i_299_n_0 ;
  wire [3:0]\badr[15]_INST_0_i_2_0 ;
  wire [0:0]\badr[15]_INST_0_i_2_1 ;
  wire [1:0]\badr[15]_INST_0_i_2_2 ;
  wire \badr[15]_INST_0_i_300_n_0 ;
  wire \badr[15]_INST_0_i_301_n_0 ;
  wire \badr[15]_INST_0_i_302_n_0 ;
  wire \badr[15]_INST_0_i_303_n_0 ;
  wire \badr[15]_INST_0_i_304_n_0 ;
  wire \badr[15]_INST_0_i_305_n_0 ;
  wire \badr[15]_INST_0_i_306_n_0 ;
  wire \badr[15]_INST_0_i_307_n_0 ;
  wire \badr[15]_INST_0_i_308_n_0 ;
  wire \badr[15]_INST_0_i_309_n_0 ;
  wire \badr[15]_INST_0_i_310_n_0 ;
  wire \badr[15]_INST_0_i_311_n_0 ;
  wire \badr[15]_INST_0_i_312_n_0 ;
  wire \badr[15]_INST_0_i_313_n_0 ;
  wire \badr[15]_INST_0_i_314_n_0 ;
  wire \badr[15]_INST_0_i_315_n_0 ;
  wire \badr[15]_INST_0_i_316_n_0 ;
  wire \badr[15]_INST_0_i_317_n_0 ;
  wire \badr[15]_INST_0_i_318_n_0 ;
  wire \badr[15]_INST_0_i_319_n_0 ;
  wire \badr[15]_INST_0_i_320_n_0 ;
  wire \badr[15]_INST_0_i_321_n_0 ;
  wire \badr[15]_INST_0_i_322_n_0 ;
  wire \badr[15]_INST_0_i_323_n_0 ;
  wire \badr[15]_INST_0_i_324_n_0 ;
  wire \badr[15]_INST_0_i_325_n_0 ;
  wire \badr[15]_INST_0_i_326_n_0 ;
  wire \badr[15]_INST_0_i_327_n_0 ;
  wire \badr[15]_INST_0_i_39_n_0 ;
  wire \badr[15]_INST_0_i_41_n_0 ;
  wire \badr[15]_INST_0_i_42_n_0 ;
  wire \badr[15]_INST_0_i_70_n_0 ;
  wire \badr[15]_INST_0_i_71_n_0 ;
  wire \badr[15]_INST_0_i_72_n_0 ;
  wire \badr[15]_INST_0_i_73_n_0 ;
  wire \badr[15]_INST_0_i_74_n_0 ;
  wire \badr[15]_INST_0_i_75_n_0 ;
  wire \badr[15]_INST_0_i_76_n_0 ;
  wire \badr[15]_INST_0_i_77_n_0 ;
  wire \badr[15]_INST_0_i_78_n_0 ;
  wire \badr[15]_INST_0_i_79_n_0 ;
  wire \badr[15]_INST_0_i_80_n_0 ;
  wire \badr[15]_INST_0_i_81_n_0 ;
  wire \badr[15]_INST_0_i_82_n_0 ;
  wire \badr[15]_INST_0_i_83_n_0 ;
  wire \badr[15]_INST_0_i_84_n_0 ;
  wire \badr[15]_INST_0_i_85_n_0 ;
  wire \badr[15]_INST_0_i_86_n_0 ;
  wire \badr[15]_INST_0_i_87_n_0 ;
  wire \badr[15]_INST_0_i_88_n_0 ;
  wire \badr[15]_INST_0_i_89_n_0 ;
  wire \badr[15]_INST_0_i_90_n_0 ;
  wire \badr[1]_INST_0_i_2 ;
  wire [2:0]\badr[2]_INST_0_i_2 ;
  wire [1:0]\badr[4]_INST_0_i_1 ;
  wire [3:0]\badr[6]_INST_0_i_2 ;
  wire \badrx[15]_INST_0_i_2_n_0 ;
  wire \badrx[15]_INST_0_i_3_n_0 ;
  wire \badrx[15]_INST_0_i_5_n_0 ;
  wire \badrx[15]_INST_0_i_6_n_0 ;
  wire \badrx[15]_INST_0_i_7_n_0 ;
  wire [0:0]bank_sel;
  wire [14:0]bbus_o;
  wire \bbus_o[0]_0 ;
  wire \bbus_o[0]_INST_0_i_1_0 ;
  wire \bbus_o[0]_INST_0_i_2_n_0 ;
  wire \bbus_o[0]_INST_0_i_3_n_0 ;
  wire \bbus_o[0]_INST_0_i_8_n_0 ;
  wire \bbus_o[1]_0 ;
  wire \bbus_o[1]_INST_0_i_1_0 ;
  wire \bbus_o[1]_INST_0_i_1_1 ;
  wire \bbus_o[1]_INST_0_i_1_2 ;
  wire \bbus_o[1]_INST_0_i_1_n_0 ;
  wire \bbus_o[1]_INST_0_i_2_n_0 ;
  wire \bbus_o[1]_INST_0_i_3_n_0 ;
  wire \bbus_o[2]_0 ;
  wire \bbus_o[2]_INST_0_i_1_0 ;
  wire \bbus_o[2]_INST_0_i_1_n_0 ;
  wire \bbus_o[2]_INST_0_i_2_n_0 ;
  wire \bbus_o[2]_INST_0_i_3_n_0 ;
  wire \bbus_o[2]_INST_0_i_8_n_0 ;
  wire \bbus_o[3]_0 ;
  wire \bbus_o[3]_INST_0_i_1_0 ;
  wire \bbus_o[3]_INST_0_i_1_n_0 ;
  wire \bbus_o[3]_INST_0_i_2_n_0 ;
  wire \bbus_o[3]_INST_0_i_3_n_0 ;
  wire \bbus_o[3]_INST_0_i_8_n_0 ;
  wire \bbus_o[4]_INST_0_i_2_n_0 ;
  wire \bbus_o[4]_INST_0_i_3_n_0 ;
  wire \bbus_o[4]_INST_0_i_45_n_0 ;
  wire \bbus_o[4]_INST_0_i_48_n_0 ;
  wire \bbus_o[4]_INST_0_i_49_0 ;
  wire \bbus_o[4]_INST_0_i_49_n_0 ;
  wire \bbus_o[4]_INST_0_i_50_n_0 ;
  wire \bbus_o[4]_INST_0_i_51_n_0 ;
  wire \bbus_o[4]_INST_0_i_52_n_0 ;
  wire \bbus_o[4]_INST_0_i_53_n_0 ;
  wire \bbus_o[4]_INST_0_i_54_n_0 ;
  wire \bbus_o[4]_INST_0_i_55_n_0 ;
  wire \bbus_o[4]_INST_0_i_56_n_0 ;
  wire \bbus_o[4]_INST_0_i_57_n_0 ;
  wire \bbus_o[4]_INST_0_i_58_n_0 ;
  wire \bbus_o[4]_INST_0_i_59_n_0 ;
  wire \bbus_o[4]_INST_0_i_60_n_0 ;
  wire \bbus_o[4]_INST_0_i_61_n_0 ;
  wire \bbus_o[4]_INST_0_i_62_n_0 ;
  wire \bbus_o[4]_INST_0_i_8_n_0 ;
  wire \bbus_o[5]_INST_0_i_8_n_0 ;
  wire \bbus_o[6]_INST_0_i_8_n_0 ;
  wire \bbus_o[7]_INST_0_i_8_n_0 ;
  wire bbus_o_0_sn_1;
  wire bbus_o_13_sn_1;
  wire bbus_o_14_sn_1;
  wire bbus_o_1_sn_1;
  wire bbus_o_2_sn_1;
  wire bbus_o_3_sn_1;
  wire bbus_o_6_sn_1;
  wire bbus_o_7_sn_1;
  wire \bcmd[0]_INST_0_i_10_n_0 ;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_13_n_0 ;
  wire \bcmd[0]_INST_0_i_14_n_0 ;
  wire \bcmd[0]_INST_0_i_15_n_0 ;
  wire \bcmd[0]_INST_0_i_16_n_0 ;
  wire \bcmd[0]_INST_0_i_17_n_0 ;
  wire \bcmd[0]_INST_0_i_18_n_0 ;
  wire \bcmd[0]_INST_0_i_19_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_20_n_0 ;
  wire \bcmd[0]_INST_0_i_21_n_0 ;
  wire \bcmd[0]_INST_0_i_22_n_0 ;
  wire \bcmd[0]_INST_0_i_23_n_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_3_n_0 ;
  wire \bcmd[0]_INST_0_i_4_n_0 ;
  wire \bcmd[0]_INST_0_i_5_n_0 ;
  wire \bcmd[0]_INST_0_i_6_n_0 ;
  wire \bcmd[0]_INST_0_i_7_n_0 ;
  wire \bcmd[0]_INST_0_i_8_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1] ;
  wire \bcmd[1]_0 ;
  wire \bcmd[1]_INST_0_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_11_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_14_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_17_n_0 ;
  wire \bcmd[1]_INST_0_i_18_n_0 ;
  wire \bcmd[1]_INST_0_i_19_n_0 ;
  wire \bcmd[1]_INST_0_i_2_n_0 ;
  wire \bcmd[1]_INST_0_i_3_n_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_6_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_8_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2]_INST_0_0 ;
  wire \bcmd[2]_INST_0_i_11_n_0 ;
  wire \bcmd[2]_INST_0_i_2_n_0 ;
  wire \bcmd[2]_INST_0_i_3_n_0 ;
  wire \bcmd[2]_INST_0_i_4_n_0 ;
  wire \bcmd[2]_INST_0_i_5_n_0 ;
  wire \bcmd[2]_INST_0_i_7_n_0 ;
  wire \bcmd[2]_INST_0_i_8_n_0 ;
  wire \bcmd[2]_INST_0_i_9_n_0 ;
  wire [4:0]bdatr;
  wire [15:0]\bdatr[15] ;
  wire [13:0]bdatw;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_INST_0_i_16_n_0 ;
  wire \bdatw[10]_INST_0_i_17_n_0 ;
  wire \bdatw[10]_INST_0_i_18_n_0 ;
  wire \bdatw[10]_INST_0_i_29_n_0 ;
  wire \bdatw[10]_INST_0_i_3_n_0 ;
  wire \bdatw[10]_INST_0_i_40_n_0 ;
  wire \bdatw[10]_INST_0_i_45_n_0 ;
  wire \bdatw[10]_INST_0_i_70_n_0 ;
  wire \bdatw[11]_0 ;
  wire \bdatw[11]_INST_0_i_16_0 ;
  wire \bdatw[11]_INST_0_i_16_n_0 ;
  wire \bdatw[11]_INST_0_i_17_n_0 ;
  wire \bdatw[11]_INST_0_i_28_n_0 ;
  wire \bdatw[11]_INST_0_i_29_n_0 ;
  wire \bdatw[11]_INST_0_i_3_n_0 ;
  wire \bdatw[11]_INST_0_i_40_n_0 ;
  wire \bdatw[11]_INST_0_i_41_n_0 ;
  wire \bdatw[11]_INST_0_i_58_n_0 ;
  wire \bdatw[12]_0 ;
  wire \bdatw[12]_INST_0_i_17_n_0 ;
  wire \bdatw[12]_INST_0_i_38_n_0 ;
  wire \bdatw[12]_INST_0_i_39_n_0 ;
  wire \bdatw[12]_INST_0_i_3_n_0 ;
  wire \bdatw[12]_INST_0_i_56_n_0 ;
  wire \bdatw[13]_INST_0_i_17_n_0 ;
  wire \bdatw[13]_INST_0_i_28_n_0 ;
  wire \bdatw[13]_INST_0_i_29_n_0 ;
  wire \bdatw[13]_INST_0_i_58_n_0 ;
  wire \bdatw[14]_INST_0_i_105_n_0 ;
  wire \bdatw[14]_INST_0_i_106_n_0 ;
  wire \bdatw[14]_INST_0_i_107_n_0 ;
  wire \bdatw[14]_INST_0_i_108_n_0 ;
  wire \bdatw[14]_INST_0_i_109_n_0 ;
  wire \bdatw[14]_INST_0_i_110_n_0 ;
  wire \bdatw[14]_INST_0_i_111_n_0 ;
  wire \bdatw[14]_INST_0_i_17_n_0 ;
  wire \bdatw[14]_INST_0_i_18_n_0 ;
  wire \bdatw[14]_INST_0_i_29_n_0 ;
  wire \bdatw[14]_INST_0_i_30_n_0 ;
  wire \bdatw[14]_INST_0_i_77_n_0 ;
  wire \bdatw[14]_INST_0_i_89_n_0 ;
  wire \bdatw[14]_INST_0_i_90_n_0 ;
  wire \bdatw[15] ;
  wire \bdatw[15]_0 ;
  wire \bdatw[15]_1 ;
  wire \bdatw[15]_2 ;
  wire \bdatw[15]_INST_0_i_100_n_0 ;
  wire \bdatw[15]_INST_0_i_101_n_0 ;
  wire \bdatw[15]_INST_0_i_103_n_0 ;
  wire \bdatw[15]_INST_0_i_104_n_0 ;
  wire \bdatw[15]_INST_0_i_105_n_0 ;
  wire \bdatw[15]_INST_0_i_106_n_0 ;
  wire \bdatw[15]_INST_0_i_107_n_0 ;
  wire \bdatw[15]_INST_0_i_108_n_0 ;
  wire \bdatw[15]_INST_0_i_109_n_0 ;
  wire \bdatw[15]_INST_0_i_117_n_0 ;
  wire \bdatw[15]_INST_0_i_129_n_0 ;
  wire \bdatw[15]_INST_0_i_12_n_0 ;
  wire \bdatw[15]_INST_0_i_13_n_0 ;
  wire \bdatw[15]_INST_0_i_140_n_0 ;
  wire \bdatw[15]_INST_0_i_141_n_0 ;
  wire \bdatw[15]_INST_0_i_142_n_0 ;
  wire \bdatw[15]_INST_0_i_143_n_0 ;
  wire \bdatw[15]_INST_0_i_144_n_0 ;
  wire \bdatw[15]_INST_0_i_145_n_0 ;
  wire \bdatw[15]_INST_0_i_146_n_0 ;
  wire \bdatw[15]_INST_0_i_147_n_0 ;
  wire \bdatw[15]_INST_0_i_148_n_0 ;
  wire \bdatw[15]_INST_0_i_149_n_0 ;
  wire \bdatw[15]_INST_0_i_150_n_0 ;
  wire \bdatw[15]_INST_0_i_151_n_0 ;
  wire \bdatw[15]_INST_0_i_152_n_0 ;
  wire \bdatw[15]_INST_0_i_153_n_0 ;
  wire \bdatw[15]_INST_0_i_154_n_0 ;
  wire \bdatw[15]_INST_0_i_155_n_0 ;
  wire \bdatw[15]_INST_0_i_156_n_0 ;
  wire \bdatw[15]_INST_0_i_157_n_0 ;
  wire \bdatw[15]_INST_0_i_158_n_0 ;
  wire \bdatw[15]_INST_0_i_159_n_0 ;
  wire \bdatw[15]_INST_0_i_160_n_0 ;
  wire \bdatw[15]_INST_0_i_161_n_0 ;
  wire \bdatw[15]_INST_0_i_162_n_0 ;
  wire \bdatw[15]_INST_0_i_163_n_0 ;
  wire \bdatw[15]_INST_0_i_164_n_0 ;
  wire \bdatw[15]_INST_0_i_165_n_0 ;
  wire \bdatw[15]_INST_0_i_166_n_0 ;
  wire \bdatw[15]_INST_0_i_167_n_0 ;
  wire \bdatw[15]_INST_0_i_168_n_0 ;
  wire \bdatw[15]_INST_0_i_171_n_0 ;
  wire \bdatw[15]_INST_0_i_172_n_0 ;
  wire \bdatw[15]_INST_0_i_173_n_0 ;
  wire \bdatw[15]_INST_0_i_177_n_0 ;
  wire \bdatw[15]_INST_0_i_178_n_0 ;
  wire \bdatw[15]_INST_0_i_179_n_0 ;
  wire \bdatw[15]_INST_0_i_180_n_0 ;
  wire \bdatw[15]_INST_0_i_181_n_0 ;
  wire \bdatw[15]_INST_0_i_182_n_0 ;
  wire \bdatw[15]_INST_0_i_183_n_0 ;
  wire \bdatw[15]_INST_0_i_184_n_0 ;
  wire \bdatw[15]_INST_0_i_185_n_0 ;
  wire \bdatw[15]_INST_0_i_186_n_0 ;
  wire \bdatw[15]_INST_0_i_187_n_0 ;
  wire \bdatw[15]_INST_0_i_188_n_0 ;
  wire \bdatw[15]_INST_0_i_189_n_0 ;
  wire \bdatw[15]_INST_0_i_190_n_0 ;
  wire \bdatw[15]_INST_0_i_191_n_0 ;
  wire \bdatw[15]_INST_0_i_192_n_0 ;
  wire \bdatw[15]_INST_0_i_193_n_0 ;
  wire \bdatw[15]_INST_0_i_194_n_0 ;
  wire \bdatw[15]_INST_0_i_195_n_0 ;
  wire \bdatw[15]_INST_0_i_196_n_0 ;
  wire \bdatw[15]_INST_0_i_197_n_0 ;
  wire \bdatw[15]_INST_0_i_198_n_0 ;
  wire \bdatw[15]_INST_0_i_199_n_0 ;
  wire \bdatw[15]_INST_0_i_19_n_0 ;
  wire \bdatw[15]_INST_0_i_202_n_0 ;
  wire \bdatw[15]_INST_0_i_203_n_0 ;
  wire \bdatw[15]_INST_0_i_204_n_0 ;
  wire \bdatw[15]_INST_0_i_205_n_0 ;
  wire \bdatw[15]_INST_0_i_206_n_0 ;
  wire \bdatw[15]_INST_0_i_207_n_0 ;
  wire \bdatw[15]_INST_0_i_208_n_0 ;
  wire \bdatw[15]_INST_0_i_209_n_0 ;
  wire \bdatw[15]_INST_0_i_222_n_0 ;
  wire \bdatw[15]_INST_0_i_223_n_0 ;
  wire \bdatw[15]_INST_0_i_224_n_0 ;
  wire \bdatw[15]_INST_0_i_225_n_0 ;
  wire \bdatw[15]_INST_0_i_226_n_0 ;
  wire \bdatw[15]_INST_0_i_227_n_0 ;
  wire \bdatw[15]_INST_0_i_228_n_0 ;
  wire \bdatw[15]_INST_0_i_229_n_0 ;
  wire \bdatw[15]_INST_0_i_231_n_0 ;
  wire \bdatw[15]_INST_0_i_232_n_0 ;
  wire \bdatw[15]_INST_0_i_233_n_0 ;
  wire \bdatw[15]_INST_0_i_234_n_0 ;
  wire \bdatw[15]_INST_0_i_235_n_0 ;
  wire \bdatw[15]_INST_0_i_236_n_0 ;
  wire \bdatw[15]_INST_0_i_237_n_0 ;
  wire \bdatw[15]_INST_0_i_238_n_0 ;
  wire \bdatw[15]_INST_0_i_239_n_0 ;
  wire \bdatw[15]_INST_0_i_240_n_0 ;
  wire \bdatw[15]_INST_0_i_241_n_0 ;
  wire \bdatw[15]_INST_0_i_242_n_0 ;
  wire \bdatw[15]_INST_0_i_243_n_0 ;
  wire \bdatw[15]_INST_0_i_244_n_0 ;
  wire \bdatw[15]_INST_0_i_245_n_0 ;
  wire \bdatw[15]_INST_0_i_246_n_0 ;
  wire \bdatw[15]_INST_0_i_247_n_0 ;
  wire \bdatw[15]_INST_0_i_248_n_0 ;
  wire \bdatw[15]_INST_0_i_249_n_0 ;
  wire \bdatw[15]_INST_0_i_250_n_0 ;
  wire \bdatw[15]_INST_0_i_251_n_0 ;
  wire \bdatw[15]_INST_0_i_252_n_0 ;
  wire \bdatw[15]_INST_0_i_253_n_0 ;
  wire \bdatw[15]_INST_0_i_254_n_0 ;
  wire \bdatw[15]_INST_0_i_255_n_0 ;
  wire \bdatw[15]_INST_0_i_256_n_0 ;
  wire \bdatw[15]_INST_0_i_257_n_0 ;
  wire \bdatw[15]_INST_0_i_258_n_0 ;
  wire \bdatw[15]_INST_0_i_259_n_0 ;
  wire \bdatw[15]_INST_0_i_260_n_0 ;
  wire \bdatw[15]_INST_0_i_261_n_0 ;
  wire \bdatw[15]_INST_0_i_262_n_0 ;
  wire \bdatw[15]_INST_0_i_263_n_0 ;
  wire \bdatw[15]_INST_0_i_264_n_0 ;
  wire \bdatw[15]_INST_0_i_40_n_0 ;
  wire \bdatw[15]_INST_0_i_41_n_0 ;
  wire \bdatw[15]_INST_0_i_57_n_0 ;
  wire \bdatw[15]_INST_0_i_58_n_0 ;
  wire \bdatw[15]_INST_0_i_59_n_0 ;
  wire \bdatw[15]_INST_0_i_60_n_0 ;
  wire \bdatw[15]_INST_0_i_61_n_0 ;
  wire \bdatw[15]_INST_0_i_62_n_0 ;
  wire \bdatw[15]_INST_0_i_63_n_0 ;
  wire \bdatw[15]_INST_0_i_64_n_0 ;
  wire \bdatw[15]_INST_0_i_65_n_0 ;
  wire \bdatw[15]_INST_0_i_66_n_0 ;
  wire \bdatw[15]_INST_0_i_67_0 ;
  wire \bdatw[15]_INST_0_i_67_n_0 ;
  wire \bdatw[15]_INST_0_i_71_n_0 ;
  wire \bdatw[15]_INST_0_i_99_n_0 ;
  wire \bdatw[8]_0 ;
  wire \bdatw[8]_INST_0_i_16_0 ;
  wire \bdatw[8]_INST_0_i_16_1 ;
  wire \bdatw[8]_INST_0_i_16_2 ;
  wire \bdatw[8]_INST_0_i_17_n_0 ;
  wire \bdatw[8]_INST_0_i_28_n_0 ;
  wire \bdatw[8]_INST_0_i_39_n_0 ;
  wire \bdatw[8]_INST_0_i_3_n_0 ;
  wire \bdatw[8]_INST_0_i_40_n_0 ;
  wire \bdatw[8]_INST_0_i_57_n_0 ;
  wire \bdatw[9]_0 ;
  wire \bdatw[9]_INST_0_i_16_0 ;
  wire \bdatw[9]_INST_0_i_16_n_0 ;
  wire \bdatw[9]_INST_0_i_17_n_0 ;
  wire \bdatw[9]_INST_0_i_39_n_0 ;
  wire \bdatw[9]_INST_0_i_3_n_0 ;
  wire \bdatw[9]_INST_0_i_44_n_0 ;
  wire \bdatw[9]_INST_0_i_69_n_0 ;
  wire bdatw_10_sn_1;
  wire bdatw_11_sn_1;
  wire bdatw_12_sn_1;
  wire bdatw_5_sn_1;
  wire bdatw_6_sn_1;
  wire bdatw_8_sn_1;
  wire bdatw_9_sn_1;
  wire brdy;
  wire [9:0]cbus_i;
  wire [15:0]\cbus_i[15] ;
  wire [4:0]ccmd;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_15_n_0 ;
  wire \ccmd[0]_INST_0_i_16_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_19_n_0 ;
  wire \ccmd[0]_INST_0_i_1_0 ;
  wire \ccmd[0]_INST_0_i_1_1 ;
  wire \ccmd[0]_INST_0_i_1_2 ;
  wire \ccmd[0]_INST_0_i_1_n_0 ;
  wire \ccmd[0]_INST_0_i_21_n_0 ;
  wire \ccmd[0]_INST_0_i_22_n_0 ;
  wire \ccmd[0]_INST_0_i_23_n_0 ;
  wire \ccmd[0]_INST_0_i_24_n_0 ;
  wire \ccmd[0]_INST_0_i_25_n_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_6_n_0 ;
  wire \ccmd[0]_INST_0_i_7_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1]_INST_0_i_10_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_12_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_15_n_0 ;
  wire \ccmd[1]_INST_0_i_16_n_0 ;
  wire \ccmd[1]_INST_0_i_17_n_0 ;
  wire \ccmd[1]_INST_0_i_18_n_0 ;
  wire \ccmd[1]_INST_0_i_19_n_0 ;
  wire \ccmd[1]_INST_0_i_1_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_6_n_0 ;
  wire \ccmd[1]_INST_0_i_7_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_10_n_0 ;
  wire \ccmd[2]_INST_0_i_11_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_13_n_0 ;
  wire \ccmd[2]_INST_0_i_14_n_0 ;
  wire \ccmd[2]_INST_0_i_16_n_0 ;
  wire \ccmd[2]_INST_0_i_17_n_0 ;
  wire \ccmd[2]_INST_0_i_18_n_0 ;
  wire \ccmd[2]_INST_0_i_19_n_0 ;
  wire \ccmd[2]_INST_0_i_1_n_0 ;
  wire \ccmd[2]_INST_0_i_20_n_0 ;
  wire \ccmd[2]_INST_0_i_2_0 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_3_0 ;
  wire \ccmd[2]_INST_0_i_3_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[2]_INST_0_i_7_n_0 ;
  wire \ccmd[2]_INST_0_i_8_n_0 ;
  wire \ccmd[2]_INST_0_i_9_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_12_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_14_n_0 ;
  wire \ccmd[3]_INST_0_i_15_n_0 ;
  wire \ccmd[3]_INST_0_i_17_n_0 ;
  wire \ccmd[3]_INST_0_i_18_n_0 ;
  wire \ccmd[3]_INST_0_i_1_n_0 ;
  wire \ccmd[3]_INST_0_i_20_n_0 ;
  wire \ccmd[3]_INST_0_i_21_n_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_8_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire \ccmd[4]_INST_0_i_11_n_0 ;
  wire \ccmd[4]_INST_0_i_12_n_0 ;
  wire \ccmd[4]_INST_0_i_13_n_0 ;
  wire \ccmd[4]_INST_0_i_14_n_0 ;
  wire \ccmd[4]_INST_0_i_15_n_0 ;
  wire \ccmd[4]_INST_0_i_16_n_0 ;
  wire \ccmd[4]_INST_0_i_17_n_0 ;
  wire \ccmd[4]_INST_0_i_18_n_0 ;
  wire \ccmd[4]_INST_0_i_19_n_0 ;
  wire \ccmd[4]_INST_0_i_20_n_0 ;
  wire \ccmd[4]_INST_0_i_2_n_0 ;
  wire \ccmd[4]_INST_0_i_3_n_0 ;
  wire \ccmd[4]_INST_0_i_4_n_0 ;
  wire \ccmd[4]_INST_0_i_5_n_0 ;
  wire \ccmd[4]_INST_0_i_6_n_0 ;
  wire \ccmd[4]_INST_0_i_7_n_0 ;
  wire \ccmd[4]_INST_0_i_8_n_0 ;
  wire \ccmd[4]_INST_0_i_9_n_0 ;
  wire ccmd_4_sn_1;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take0_fl_reg_0;
  wire ctl_bcc_take1_fl;
  wire ctl_bcc_take1_fl_reg_0;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_16;
  wire ctl_fetch0_fl_i_16_0;
  wire ctl_fetch0_fl_i_8;
  wire ctl_fetch0_fl_reg_0;
  wire ctl_fetch0_fl_reg_1;
  wire ctl_fetch0_fl_reg_2;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch1_fl_i_16;
  wire ctl_fetch1_fl_i_20_n_0;
  wire ctl_fetch1_fl_i_36_n_0;
  wire ctl_fetch1_fl_reg_i_6;
  wire ctl_fetch_ext_fl;
  wire ctl_fetch_ext_fl_i_1_n_0;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire ctl_sp_dec0;
  wire ctl_sr_ldie0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  (* DONT_TOUCH *) wire [15:0]eir;
  wire \eir_fl[15]_i_1_n_0 ;
  wire \eir_fl[1]_i_1_n_0 ;
  wire \eir_fl[2]_i_1_n_0 ;
  wire \eir_fl[3]_i_1_n_0 ;
  wire \eir_fl[4]_i_1_n_0 ;
  wire \eir_fl[5]_i_1_n_0 ;
  wire \eir_fl[6]_i_1_n_0 ;
  wire \eir_fl[6]_i_2_n_0 ;
  wire \eir_fl_reg_n_0_[0] ;
  wire \eir_fl_reg_n_0_[10] ;
  wire \eir_fl_reg_n_0_[11] ;
  wire \eir_fl_reg_n_0_[12] ;
  wire \eir_fl_reg_n_0_[13] ;
  wire \eir_fl_reg_n_0_[14] ;
  wire \eir_fl_reg_n_0_[15] ;
  wire \eir_fl_reg_n_0_[1] ;
  wire \eir_fl_reg_n_0_[2] ;
  wire \eir_fl_reg_n_0_[3] ;
  wire \eir_fl_reg_n_0_[4] ;
  wire \eir_fl_reg_n_0_[5] ;
  wire \eir_fl_reg_n_0_[6] ;
  wire \eir_fl_reg_n_0_[7] ;
  wire \eir_fl_reg_n_0_[8] ;
  wire \eir_fl_reg_n_0_[9] ;
  wire [12:0]fadr;
  wire \fadr[15]_INST_0_i_11_n_0 ;
  wire \fadr[15]_INST_0_i_13_n_0 ;
  wire \fadr[15]_INST_0_i_16_n_0 ;
  wire \fadr[15]_INST_0_i_18_n_0 ;
  wire [0:0]\fadr[3] ;
  wire fadr_1_fl;
  wire [1:0]fch_irq_lev;
  wire fch_irq_lev0;
  wire \fch_irq_lev[0]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_2_0 ;
  wire \fch_irq_lev[1]_i_3_n_0 ;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev[1]_i_5_n_0 ;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire fch_irq_req_fl_reg_0;
  (* DONT_TOUCH *) wire fch_issu1;
  wire fch_issu1_fl;
  wire fch_issu1_inferred_i_100_n_0;
  wire fch_issu1_inferred_i_101_n_0;
  wire fch_issu1_inferred_i_102_n_0;
  wire fch_issu1_inferred_i_103_n_0;
  wire fch_issu1_inferred_i_104_n_0;
  wire fch_issu1_inferred_i_105_n_0;
  wire fch_issu1_inferred_i_106_n_0;
  wire fch_issu1_inferred_i_107_n_0;
  wire fch_issu1_inferred_i_108_n_0;
  wire fch_issu1_inferred_i_109_n_0;
  wire fch_issu1_inferred_i_110_n_0;
  wire fch_issu1_inferred_i_111_n_0;
  wire fch_issu1_inferred_i_113_n_0;
  wire fch_issu1_inferred_i_114_n_0;
  wire fch_issu1_inferred_i_115_n_0;
  wire fch_issu1_inferred_i_116_n_0;
  wire fch_issu1_inferred_i_117_n_0;
  wire fch_issu1_inferred_i_118_n_0;
  wire fch_issu1_inferred_i_119_n_0;
  wire fch_issu1_inferred_i_120_n_0;
  wire fch_issu1_inferred_i_121_n_0;
  wire fch_issu1_inferred_i_122_n_0;
  wire fch_issu1_inferred_i_123_n_0;
  wire fch_issu1_inferred_i_124_n_0;
  wire fch_issu1_inferred_i_125_n_0;
  wire fch_issu1_inferred_i_126_n_0;
  wire fch_issu1_inferred_i_127_n_0;
  wire fch_issu1_inferred_i_128_n_0;
  wire fch_issu1_inferred_i_129_n_0;
  wire fch_issu1_inferred_i_130_n_0;
  wire fch_issu1_inferred_i_131_n_0;
  wire fch_issu1_inferred_i_132_n_0;
  wire fch_issu1_inferred_i_133_n_0;
  wire fch_issu1_inferred_i_134_n_0;
  wire fch_issu1_inferred_i_135_n_0;
  wire fch_issu1_inferred_i_136_n_0;
  wire fch_issu1_inferred_i_137_n_0;
  wire fch_issu1_inferred_i_138_n_0;
  wire fch_issu1_inferred_i_139_n_0;
  wire fch_issu1_inferred_i_140_n_0;
  wire fch_issu1_inferred_i_141_n_0;
  wire fch_issu1_inferred_i_142_n_0;
  wire fch_issu1_inferred_i_143_n_0;
  wire fch_issu1_inferred_i_145_n_0;
  wire fch_issu1_inferred_i_146_n_0;
  wire fch_issu1_inferred_i_147_n_0;
  wire fch_issu1_inferred_i_148_n_0;
  wire fch_issu1_inferred_i_149_n_0;
  wire fch_issu1_inferred_i_14_n_0;
  wire fch_issu1_inferred_i_150_n_0;
  wire fch_issu1_inferred_i_151_n_0;
  wire fch_issu1_inferred_i_152_n_0;
  wire fch_issu1_inferred_i_153_n_0;
  wire fch_issu1_inferred_i_154_n_0;
  wire fch_issu1_inferred_i_155_n_0;
  wire fch_issu1_inferred_i_156_n_0;
  wire fch_issu1_inferred_i_157_n_0;
  wire fch_issu1_inferred_i_158_n_0;
  wire fch_issu1_inferred_i_159_n_0;
  wire fch_issu1_inferred_i_15_n_0;
  wire fch_issu1_inferred_i_160_n_0;
  wire fch_issu1_inferred_i_161_n_0;
  wire fch_issu1_inferred_i_162_n_0;
  wire fch_issu1_inferred_i_163_n_0;
  wire fch_issu1_inferred_i_164_n_0;
  wire fch_issu1_inferred_i_165_n_0;
  wire fch_issu1_inferred_i_167_n_0;
  wire fch_issu1_inferred_i_168_n_0;
  wire fch_issu1_inferred_i_169_n_0;
  wire fch_issu1_inferred_i_16_n_0;
  wire fch_issu1_inferred_i_170_n_0;
  wire fch_issu1_inferred_i_171_n_0;
  wire fch_issu1_inferred_i_172_n_0;
  wire fch_issu1_inferred_i_173_n_0;
  wire fch_issu1_inferred_i_174_n_0;
  wire fch_issu1_inferred_i_175_n_0;
  wire fch_issu1_inferred_i_176_n_0;
  wire fch_issu1_inferred_i_177_n_0;
  wire fch_issu1_inferred_i_178_n_0;
  wire fch_issu1_inferred_i_179_n_0;
  wire fch_issu1_inferred_i_17_n_0;
  wire fch_issu1_inferred_i_180_n_0;
  wire fch_issu1_inferred_i_181_n_0;
  wire fch_issu1_inferred_i_182_n_0;
  wire fch_issu1_inferred_i_183_n_0;
  wire fch_issu1_inferred_i_184_n_0;
  wire fch_issu1_inferred_i_185_n_0;
  wire fch_issu1_inferred_i_186_n_0;
  wire fch_issu1_inferred_i_187_n_0;
  wire fch_issu1_inferred_i_188_n_0;
  wire fch_issu1_inferred_i_189_n_0;
  wire fch_issu1_inferred_i_190_n_0;
  wire fch_issu1_inferred_i_191_n_0;
  wire fch_issu1_inferred_i_192_n_0;
  wire fch_issu1_inferred_i_193_n_0;
  wire fch_issu1_inferred_i_194_n_0;
  wire fch_issu1_inferred_i_195_n_0;
  wire fch_issu1_inferred_i_196_n_0;
  wire fch_issu1_inferred_i_197_n_0;
  wire fch_issu1_inferred_i_198_n_0;
  wire fch_issu1_inferred_i_25_n_0;
  wire fch_issu1_inferred_i_26_n_0;
  wire fch_issu1_inferred_i_27_n_0;
  wire fch_issu1_inferred_i_36_n_0;
  wire fch_issu1_inferred_i_37_n_0;
  wire fch_issu1_inferred_i_39_n_0;
  wire fch_issu1_inferred_i_43_n_0;
  wire fch_issu1_inferred_i_44_n_0;
  wire fch_issu1_inferred_i_45_n_0;
  wire fch_issu1_inferred_i_46_n_0;
  wire fch_issu1_inferred_i_47_n_0;
  wire fch_issu1_inferred_i_49_0;
  wire fch_issu1_inferred_i_49_n_0;
  wire fch_issu1_inferred_i_51_n_0;
  wire fch_issu1_inferred_i_52_n_0;
  wire fch_issu1_inferred_i_53_n_0;
  wire fch_issu1_inferred_i_54_n_0;
  wire fch_issu1_inferred_i_55_n_0;
  wire fch_issu1_inferred_i_56_n_0;
  wire fch_issu1_inferred_i_57_n_0;
  wire fch_issu1_inferred_i_58_n_0;
  wire fch_issu1_inferred_i_62_n_0;
  wire fch_issu1_inferred_i_63_n_0;
  wire fch_issu1_inferred_i_64_n_0;
  wire fch_issu1_inferred_i_65_n_0;
  wire fch_issu1_inferred_i_66_n_0;
  wire fch_issu1_inferred_i_67_n_0;
  wire fch_issu1_inferred_i_69_n_0;
  wire fch_issu1_inferred_i_71_n_0;
  wire fch_issu1_inferred_i_72_n_0;
  wire fch_issu1_inferred_i_73_n_0;
  wire fch_issu1_inferred_i_76_n_0;
  wire fch_issu1_inferred_i_77_n_0;
  wire fch_issu1_inferred_i_78_n_0;
  wire fch_issu1_inferred_i_81_n_0;
  wire fch_issu1_inferred_i_82_n_0;
  wire fch_issu1_inferred_i_83_n_0;
  wire fch_issu1_inferred_i_84_n_0;
  wire fch_issu1_inferred_i_85_n_0;
  wire fch_issu1_inferred_i_86_n_0;
  wire fch_issu1_inferred_i_87_n_0;
  wire fch_issu1_inferred_i_88_n_0;
  wire fch_issu1_inferred_i_89_n_0;
  wire fch_issu1_inferred_i_90_n_0;
  wire fch_issu1_inferred_i_91_n_0;
  wire fch_issu1_inferred_i_92_n_0;
  wire fch_issu1_inferred_i_93_n_0;
  wire fch_issu1_inferred_i_94_n_0;
  wire fch_issu1_inferred_i_95_n_0;
  wire fch_issu1_inferred_i_96_n_0;
  wire fch_issu1_inferred_i_97_n_0;
  wire fch_issu1_inferred_i_99_n_0;
  wire fch_issu1_ir;
  wire fch_leir_nir_reg;
  wire fch_leir_nir_reg_0;
  wire fch_leir_nir_reg_1;
  wire fch_leir_nir_reg_2;
  wire fch_leir_nir_reg_3;
  wire fch_leir_nir_reg_4;
  wire fch_leir_nir_reg_5;
  wire fch_leir_nir_reg_6;
  wire fch_leir_nir_reg_7;
  wire fch_memacc1;
  wire fch_nir_lir;
  wire [12:0]fch_pc;
  wire fch_pc_nx2_carry__0_n_0;
  wire fch_pc_nx2_carry__0_n_1;
  wire fch_pc_nx2_carry__0_n_2;
  wire fch_pc_nx2_carry__0_n_3;
  wire fch_pc_nx2_carry__1_n_0;
  wire fch_pc_nx2_carry__1_n_1;
  wire fch_pc_nx2_carry__1_n_2;
  wire fch_pc_nx2_carry__1_n_3;
  wire fch_pc_nx2_carry__2_n_1;
  wire fch_pc_nx2_carry__2_n_2;
  wire fch_pc_nx2_carry__2_n_3;
  wire fch_pc_nx2_carry_n_0;
  wire fch_pc_nx2_carry_n_1;
  wire fch_pc_nx2_carry_n_2;
  wire fch_pc_nx2_carry_n_3;
  wire fch_pc_nx4_carry__0_n_0;
  wire fch_pc_nx4_carry__0_n_1;
  wire fch_pc_nx4_carry__0_n_2;
  wire fch_pc_nx4_carry__0_n_3;
  wire fch_pc_nx4_carry__0_n_4;
  wire fch_pc_nx4_carry__0_n_5;
  wire fch_pc_nx4_carry__0_n_6;
  wire fch_pc_nx4_carry__0_n_7;
  wire fch_pc_nx4_carry__1_n_0;
  wire fch_pc_nx4_carry__1_n_1;
  wire fch_pc_nx4_carry__1_n_2;
  wire fch_pc_nx4_carry__1_n_3;
  wire fch_pc_nx4_carry__1_n_4;
  wire fch_pc_nx4_carry__1_n_5;
  wire fch_pc_nx4_carry__1_n_6;
  wire fch_pc_nx4_carry__1_n_7;
  wire fch_pc_nx4_carry__2_n_2;
  wire fch_pc_nx4_carry__2_n_3;
  wire fch_pc_nx4_carry_n_0;
  wire fch_pc_nx4_carry_n_1;
  wire fch_pc_nx4_carry_n_2;
  wire fch_pc_nx4_carry_n_3;
  wire fch_pc_nx4_carry_n_4;
  wire fch_pc_nx4_carry_n_5;
  wire fch_pc_nx4_carry_n_6;
  wire fch_pc_nx4_carry_n_7;
  wire fch_term;
  wire fch_term_fl;
  wire fch_wrbufn1;
  wire fctl_n_133;
  wire fctl_n_150;
  wire fctl_n_151;
  wire fctl_n_152;
  wire fctl_n_153;
  wire fctl_n_154;
  wire fctl_n_155;
  wire fctl_n_156;
  wire fctl_n_157;
  wire fctl_n_158;
  wire fctl_n_67;
  wire fctl_n_85;
  wire fctl_n_86;
  wire fctl_n_87;
  wire fctl_n_88;
  wire fctl_n_89;
  wire fctl_n_91;
  wire fctl_n_94;
  wire fctl_n_95;
  wire fctl_n_96;
  wire [15:0]fdat;
  wire fdat_0_sn_1;
  wire fdat_12_sn_1;
  wire fdat_5_sn_1;
  wire [15:0]fdatx;
  wire fdatx_14_sn_1;
  wire fdatx_5_sn_1;
  wire [1:0]\grn[15]_i_3__5 ;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[15] ;
  wire [2:0]\grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \i_/bbus_o[0]_INST_0_i_18 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_20 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_20_0 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_21 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_21_0 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_22 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_22_0 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_23 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_23_0 ;
  wire [4:0]\i_/bdatw[12]_INST_0_i_64 ;
  wire [15:0]\i_/rgf_c1bus_wb[4]_i_86 ;
  wire [15:0]\i_/rgf_c1bus_wb[4]_i_87 ;
  wire [14:0]\i_/rgf_c1bus_wb[4]_i_96 ;
  (* DONT_TOUCH *) wire [15:0]ir0;
  wire [15:0]ir0_fl;
  wire [0:0]ir0_id;
  wire [21:20]ir0_id_fl;
  wire \ir0_id_fl[21]_i_4_n_0 ;
  (* DONT_TOUCH *) wire [15:0]ir1;
  wire [15:0]ir1_fl;
  wire [21:20]ir1_id_fl;
  wire \ir1_id_fl_reg[20]_0 ;
  wire \ir1_id_fl_reg[21]_0 ;
  wire ir1_inferred_i_17_n_0;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire [24:12]lir_id_0;
  wire [15:0]nir;
  wire [24:12]nir_id;
  wire \nir_id[12]_i_2_n_0 ;
  wire \nir_id[12]_i_3_n_0 ;
  wire \nir_id[12]_i_4_n_0 ;
  wire \nir_id[13]_i_2_n_0 ;
  wire \nir_id[13]_i_3_n_0 ;
  wire \nir_id[13]_i_4_n_0 ;
  wire \nir_id[13]_i_5_n_0 ;
  wire \nir_id[13]_i_6_n_0 ;
  wire \nir_id[14]_i_10_n_0 ;
  wire \nir_id[14]_i_11_n_0 ;
  wire \nir_id[14]_i_12_n_0 ;
  wire \nir_id[14]_i_13_n_0 ;
  wire \nir_id[14]_i_2_n_0 ;
  wire \nir_id[14]_i_3_n_0 ;
  wire \nir_id[14]_i_4_n_0 ;
  wire \nir_id[14]_i_5_n_0 ;
  wire \nir_id[14]_i_6_n_0 ;
  wire \nir_id[14]_i_7_n_0 ;
  wire \nir_id[14]_i_8_n_0 ;
  wire \nir_id[14]_i_9_n_0 ;
  wire \nir_id[16]_i_2_n_0 ;
  wire \nir_id[16]_i_3_n_0 ;
  wire \nir_id[16]_i_4_n_0 ;
  wire \nir_id[17]_i_2_n_0 ;
  wire \nir_id[17]_i_3_n_0 ;
  wire \nir_id[17]_i_4_n_0 ;
  wire \nir_id[17]_i_5_n_0 ;
  wire \nir_id[17]_i_6_n_0 ;
  wire \nir_id[17]_i_7_n_0 ;
  wire \nir_id[18]_i_2_n_0 ;
  wire \nir_id[18]_i_3_n_0 ;
  wire \nir_id[18]_i_4_n_0 ;
  wire \nir_id[18]_i_5_n_0 ;
  wire \nir_id[18]_i_6_n_0 ;
  wire \nir_id[18]_i_7_n_0 ;
  wire \nir_id[18]_i_8_n_0 ;
  wire \nir_id[19]_i_2_n_0 ;
  wire \nir_id[19]_i_3_n_0 ;
  wire \nir_id[19]_i_4_n_0 ;
  wire \nir_id[19]_i_5_n_0 ;
  wire \nir_id[19]_i_6_n_0 ;
  wire \nir_id[19]_i_7_n_0 ;
  wire \nir_id[24]_i_10_n_0 ;
  wire \nir_id[24]_i_11_n_0 ;
  wire \nir_id[24]_i_12_n_0 ;
  wire \nir_id[24]_i_13_n_0 ;
  wire \nir_id[24]_i_5_n_0 ;
  wire \nir_id[24]_i_6_n_0 ;
  wire \nir_id[24]_i_7_n_0 ;
  wire \nir_id[24]_i_8_n_0 ;
  wire [1:0]\nir_id_reg[21]_0 ;
  wire \nir_id_reg[24]_0 ;
  wire [0:0]p_0_in;
  wire [4:0]p_0_in2_in;
  wire p_0_in_1;
  wire [0:0]p_1_in;
  wire [4:0]p_1_in3_in;
  wire p_2_in;
  wire [12:0]p_2_in_0;
  wire [15:0]\pc0_reg[15]_0 ;
  wire [15:0]\pc0_reg[15]_1 ;
  wire pc10_carry__0_n_0;
  wire pc10_carry__0_n_1;
  wire pc10_carry__0_n_2;
  wire pc10_carry__0_n_3;
  wire pc10_carry__0_n_4;
  wire pc10_carry__0_n_5;
  wire pc10_carry__0_n_6;
  wire pc10_carry__0_n_7;
  wire pc10_carry__1_n_0;
  wire pc10_carry__1_n_1;
  wire pc10_carry__1_n_2;
  wire pc10_carry__1_n_3;
  wire pc10_carry__1_n_4;
  wire pc10_carry__1_n_5;
  wire pc10_carry__1_n_6;
  wire pc10_carry__1_n_7;
  wire pc10_carry__2_n_1;
  wire pc10_carry__2_n_2;
  wire pc10_carry__2_n_3;
  wire pc10_carry__2_n_4;
  wire pc10_carry__2_n_5;
  wire pc10_carry__2_n_6;
  wire pc10_carry__2_n_7;
  wire pc10_carry_n_0;
  wire pc10_carry_n_1;
  wire pc10_carry_n_2;
  wire pc10_carry_n_3;
  wire pc10_carry_n_4;
  wire pc10_carry_n_5;
  wire pc10_carry_n_6;
  wire pc10_carry_n_7;
  wire [15:0]\pc1_reg[15]_0 ;
  wire [2:0]\pc1_reg[15]_1 ;
  wire \pc[14]_i_5_n_0 ;
  wire \pc_reg[13] ;
  wire \pc_reg[14] ;
  wire [2:0]\pc_reg[15] ;
  wire [15:0]\pc_reg[15]_0 ;
  wire \pc_reg[15]_1 ;
  wire \read_cyc_reg[1] ;
  wire \read_cyc_reg[1]_0 ;
  wire \rgf_c0bus_wb[0]_i_11_n_0 ;
  wire \rgf_c0bus_wb[0]_i_12_n_0 ;
  wire \rgf_c0bus_wb[0]_i_15_n_0 ;
  wire \rgf_c0bus_wb[0]_i_16_n_0 ;
  wire \rgf_c0bus_wb[0]_i_2_0 ;
  wire \rgf_c0bus_wb[0]_i_2_1 ;
  wire \rgf_c0bus_wb[0]_i_2_n_0 ;
  wire \rgf_c0bus_wb[0]_i_5_n_0 ;
  wire \rgf_c0bus_wb[0]_i_6_n_0 ;
  wire \rgf_c0bus_wb[0]_i_7_n_0 ;
  wire \rgf_c0bus_wb[0]_i_8_n_0 ;
  wire \rgf_c0bus_wb[0]_i_9_n_0 ;
  wire \rgf_c0bus_wb[10]_i_11_n_0 ;
  wire \rgf_c0bus_wb[10]_i_12_n_0 ;
  wire \rgf_c0bus_wb[10]_i_13_n_0 ;
  wire \rgf_c0bus_wb[10]_i_15_n_0 ;
  wire \rgf_c0bus_wb[10]_i_16_n_0 ;
  wire \rgf_c0bus_wb[10]_i_23_n_0 ;
  wire \rgf_c0bus_wb[10]_i_25_n_0 ;
  wire \rgf_c0bus_wb[10]_i_26_n_0 ;
  wire \rgf_c0bus_wb[10]_i_3_n_0 ;
  wire \rgf_c0bus_wb[10]_i_4_0 ;
  wire \rgf_c0bus_wb[10]_i_4_1 ;
  wire \rgf_c0bus_wb[10]_i_4_n_0 ;
  wire \rgf_c0bus_wb[10]_i_5_n_0 ;
  wire \rgf_c0bus_wb[11]_i_11_0 ;
  wire \rgf_c0bus_wb[11]_i_12_n_0 ;
  wire \rgf_c0bus_wb[11]_i_14_n_0 ;
  wire \rgf_c0bus_wb[11]_i_15_n_0 ;
  wire \rgf_c0bus_wb[11]_i_16_n_0 ;
  wire \rgf_c0bus_wb[11]_i_17_n_0 ;
  wire \rgf_c0bus_wb[11]_i_18_n_0 ;
  wire \rgf_c0bus_wb[11]_i_19_n_0 ;
  wire \rgf_c0bus_wb[11]_i_27_n_0 ;
  wire \rgf_c0bus_wb[11]_i_2_n_0 ;
  wire \rgf_c0bus_wb[11]_i_3_0 ;
  wire \rgf_c0bus_wb[11]_i_4_0 ;
  wire \rgf_c0bus_wb[11]_i_4_n_0 ;
  wire \rgf_c0bus_wb[11]_i_5_0 ;
  wire \rgf_c0bus_wb[11]_i_5_n_0 ;
  wire \rgf_c0bus_wb[11]_i_6_n_0 ;
  wire \rgf_c0bus_wb[11]_i_7_n_0 ;
  wire \rgf_c0bus_wb[12]_i_10_n_0 ;
  wire \rgf_c0bus_wb[12]_i_11_n_0 ;
  wire \rgf_c0bus_wb[12]_i_12_n_0 ;
  wire \rgf_c0bus_wb[12]_i_13_n_0 ;
  wire \rgf_c0bus_wb[12]_i_15_n_0 ;
  wire \rgf_c0bus_wb[12]_i_2_0 ;
  wire \rgf_c0bus_wb[12]_i_2_n_0 ;
  wire \rgf_c0bus_wb[12]_i_3_0 ;
  wire \rgf_c0bus_wb[12]_i_3_1 ;
  wire \rgf_c0bus_wb[12]_i_3_n_0 ;
  wire \rgf_c0bus_wb[12]_i_4_n_0 ;
  wire \rgf_c0bus_wb[12]_i_5_n_0 ;
  wire \rgf_c0bus_wb[12]_i_6_n_0 ;
  wire \rgf_c0bus_wb[12]_i_7_n_0 ;
  wire \rgf_c0bus_wb[12]_i_9_n_0 ;
  wire \rgf_c0bus_wb[13]_i_10_0 ;
  wire \rgf_c0bus_wb[13]_i_11_n_0 ;
  wire \rgf_c0bus_wb[13]_i_12_n_0 ;
  wire \rgf_c0bus_wb[13]_i_13_n_0 ;
  wire \rgf_c0bus_wb[13]_i_16_n_0 ;
  wire \rgf_c0bus_wb[13]_i_17_n_0 ;
  wire \rgf_c0bus_wb[13]_i_18_n_0 ;
  wire \rgf_c0bus_wb[13]_i_25_n_0 ;
  wire \rgf_c0bus_wb[13]_i_2_0 ;
  wire \rgf_c0bus_wb[13]_i_2_1 ;
  wire \rgf_c0bus_wb[13]_i_2_2 ;
  wire \rgf_c0bus_wb[13]_i_2_n_0 ;
  wire \rgf_c0bus_wb[13]_i_4_0 ;
  wire \rgf_c0bus_wb[13]_i_4_n_0 ;
  wire \rgf_c0bus_wb[13]_i_5_n_0 ;
  wire \rgf_c0bus_wb[13]_i_6_n_0 ;
  wire \rgf_c0bus_wb[13]_i_7_n_0 ;
  wire \rgf_c0bus_wb[13]_i_8_n_0 ;
  wire \rgf_c0bus_wb[13]_i_9_n_0 ;
  wire \rgf_c0bus_wb[14]_i_10_n_0 ;
  wire \rgf_c0bus_wb[14]_i_11_n_0 ;
  wire \rgf_c0bus_wb[14]_i_13_n_0 ;
  wire \rgf_c0bus_wb[14]_i_14_n_0 ;
  wire \rgf_c0bus_wb[14]_i_15_n_0 ;
  wire \rgf_c0bus_wb[14]_i_16_n_0 ;
  wire \rgf_c0bus_wb[14]_i_17_n_0 ;
  wire \rgf_c0bus_wb[14]_i_2_n_0 ;
  wire \rgf_c0bus_wb[14]_i_4_n_0 ;
  wire \rgf_c0bus_wb[14]_i_5_0 ;
  wire \rgf_c0bus_wb[14]_i_5_n_0 ;
  wire \rgf_c0bus_wb[14]_i_7_n_0 ;
  wire \rgf_c0bus_wb[14]_i_8_n_0 ;
  wire \rgf_c0bus_wb[14]_i_9_n_0 ;
  wire \rgf_c0bus_wb[15]_i_10_n_0 ;
  wire \rgf_c0bus_wb[15]_i_11_n_0 ;
  wire \rgf_c0bus_wb[15]_i_12_n_0 ;
  wire \rgf_c0bus_wb[15]_i_13_n_0 ;
  wire \rgf_c0bus_wb[15]_i_14_n_0 ;
  wire \rgf_c0bus_wb[15]_i_15_n_0 ;
  wire \rgf_c0bus_wb[15]_i_16_n_0 ;
  wire \rgf_c0bus_wb[15]_i_17_n_0 ;
  wire \rgf_c0bus_wb[15]_i_19_n_0 ;
  wire \rgf_c0bus_wb[15]_i_20_n_0 ;
  wire \rgf_c0bus_wb[15]_i_22_n_0 ;
  wire \rgf_c0bus_wb[15]_i_24_n_0 ;
  wire \rgf_c0bus_wb[15]_i_2_n_0 ;
  wire \rgf_c0bus_wb[15]_i_4_0 ;
  wire \rgf_c0bus_wb[15]_i_4_1 ;
  wire \rgf_c0bus_wb[15]_i_4_2 ;
  wire \rgf_c0bus_wb[15]_i_4_n_0 ;
  wire \rgf_c0bus_wb[15]_i_7_0 ;
  wire \rgf_c0bus_wb[15]_i_7_n_0 ;
  wire \rgf_c0bus_wb[15]_i_8_0 ;
  wire \rgf_c0bus_wb[15]_i_8_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10_n_0 ;
  wire \rgf_c0bus_wb[1]_i_11_n_0 ;
  wire \rgf_c0bus_wb[1]_i_13_n_0 ;
  wire \rgf_c0bus_wb[1]_i_14_n_0 ;
  wire \rgf_c0bus_wb[1]_i_15_n_0 ;
  wire \rgf_c0bus_wb[1]_i_2_n_0 ;
  wire \rgf_c0bus_wb[1]_i_3_0 ;
  wire \rgf_c0bus_wb[1]_i_3_n_0 ;
  wire \rgf_c0bus_wb[1]_i_4_n_0 ;
  wire \rgf_c0bus_wb[1]_i_5_n_0 ;
  wire \rgf_c0bus_wb[1]_i_7_n_0 ;
  wire \rgf_c0bus_wb[1]_i_8_n_0 ;
  wire \rgf_c0bus_wb[1]_i_9_n_0 ;
  wire \rgf_c0bus_wb[2]_i_10_n_0 ;
  wire \rgf_c0bus_wb[2]_i_11_n_0 ;
  wire \rgf_c0bus_wb[2]_i_12_n_0 ;
  wire \rgf_c0bus_wb[2]_i_13_n_0 ;
  wire \rgf_c0bus_wb[2]_i_15_n_0 ;
  wire \rgf_c0bus_wb[2]_i_16_n_0 ;
  wire \rgf_c0bus_wb[2]_i_17_n_0 ;
  wire \rgf_c0bus_wb[2]_i_2_0 ;
  wire \rgf_c0bus_wb[2]_i_2_n_0 ;
  wire \rgf_c0bus_wb[2]_i_3_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4_n_0 ;
  wire \rgf_c0bus_wb[2]_i_6_n_0 ;
  wire \rgf_c0bus_wb[2]_i_8_n_0 ;
  wire \rgf_c0bus_wb[2]_i_9_n_0 ;
  wire \rgf_c0bus_wb[3]_i_10_n_0 ;
  wire \rgf_c0bus_wb[3]_i_11_n_0 ;
  wire \rgf_c0bus_wb[3]_i_12_n_0 ;
  wire \rgf_c0bus_wb[3]_i_13_n_0 ;
  wire \rgf_c0bus_wb[3]_i_14_n_0 ;
  wire \rgf_c0bus_wb[3]_i_15_n_0 ;
  wire \rgf_c0bus_wb[3]_i_16_n_0 ;
  wire \rgf_c0bus_wb[3]_i_17_n_0 ;
  wire \rgf_c0bus_wb[3]_i_18_n_0 ;
  wire \rgf_c0bus_wb[3]_i_2_n_0 ;
  wire \rgf_c0bus_wb[3]_i_4_n_0 ;
  wire \rgf_c0bus_wb[3]_i_5_n_0 ;
  wire \rgf_c0bus_wb[3]_i_6_n_0 ;
  wire \rgf_c0bus_wb[3]_i_7_n_0 ;
  wire \rgf_c0bus_wb[4]_i_10_n_0 ;
  wire \rgf_c0bus_wb[4]_i_13_n_0 ;
  wire \rgf_c0bus_wb[4]_i_14_n_0 ;
  wire \rgf_c0bus_wb[4]_i_15_n_0 ;
  wire \rgf_c0bus_wb[4]_i_16_n_0 ;
  wire \rgf_c0bus_wb[4]_i_17_n_0 ;
  wire \rgf_c0bus_wb[4]_i_20_n_0 ;
  wire \rgf_c0bus_wb[4]_i_2_0 ;
  wire \rgf_c0bus_wb[4]_i_2_1 ;
  wire \rgf_c0bus_wb[4]_i_2_n_0 ;
  wire \rgf_c0bus_wb[4]_i_3_0 ;
  wire \rgf_c0bus_wb[4]_i_3_1 ;
  wire \rgf_c0bus_wb[4]_i_3_n_0 ;
  wire \rgf_c0bus_wb[4]_i_4_n_0 ;
  wire \rgf_c0bus_wb[4]_i_5_0 ;
  wire \rgf_c0bus_wb[4]_i_5_n_0 ;
  wire \rgf_c0bus_wb[4]_i_6_0 ;
  wire \rgf_c0bus_wb[4]_i_6_1 ;
  wire \rgf_c0bus_wb[4]_i_6_n_0 ;
  wire \rgf_c0bus_wb[4]_i_9_n_0 ;
  wire \rgf_c0bus_wb[5]_i_10_n_0 ;
  wire \rgf_c0bus_wb[5]_i_11_n_0 ;
  wire \rgf_c0bus_wb[5]_i_12_n_0 ;
  wire \rgf_c0bus_wb[5]_i_13_n_0 ;
  wire \rgf_c0bus_wb[5]_i_15_n_0 ;
  wire \rgf_c0bus_wb[5]_i_16_n_0 ;
  wire \rgf_c0bus_wb[5]_i_17_n_0 ;
  wire \rgf_c0bus_wb[5]_i_2_0 ;
  wire \rgf_c0bus_wb[5]_i_2_1 ;
  wire \rgf_c0bus_wb[5]_i_2_n_0 ;
  wire \rgf_c0bus_wb[5]_i_3_0 ;
  wire \rgf_c0bus_wb[5]_i_3_1 ;
  wire \rgf_c0bus_wb[5]_i_3_2 ;
  wire \rgf_c0bus_wb[5]_i_3_n_0 ;
  wire \rgf_c0bus_wb[5]_i_4_n_0 ;
  wire \rgf_c0bus_wb[5]_i_5_n_0 ;
  wire \rgf_c0bus_wb[5]_i_6_n_0 ;
  wire \rgf_c0bus_wb[5]_i_8_n_0 ;
  wire \rgf_c0bus_wb[5]_i_9_n_0 ;
  wire \rgf_c0bus_wb[6]_i_10_n_0 ;
  wire \rgf_c0bus_wb[6]_i_11_n_0 ;
  wire \rgf_c0bus_wb[6]_i_13_n_0 ;
  wire \rgf_c0bus_wb[6]_i_15_n_0 ;
  wire \rgf_c0bus_wb[6]_i_16_n_0 ;
  wire \rgf_c0bus_wb[6]_i_2_n_0 ;
  wire \rgf_c0bus_wb[6]_i_3_n_0 ;
  wire \rgf_c0bus_wb[6]_i_4_n_0 ;
  wire \rgf_c0bus_wb[6]_i_7_n_0 ;
  wire \rgf_c0bus_wb[6]_i_8_n_0 ;
  wire \rgf_c0bus_wb[6]_i_9_n_0 ;
  wire \rgf_c0bus_wb[7]_i_13_n_0 ;
  wire \rgf_c0bus_wb[7]_i_14_n_0 ;
  wire \rgf_c0bus_wb[7]_i_2_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3_n_0 ;
  wire \rgf_c0bus_wb[7]_i_4_n_0 ;
  wire \rgf_c0bus_wb[7]_i_5_n_0 ;
  wire \rgf_c0bus_wb[7]_i_9_n_0 ;
  wire \rgf_c0bus_wb[8]_i_10_n_0 ;
  wire \rgf_c0bus_wb[8]_i_11_n_0 ;
  wire \rgf_c0bus_wb[8]_i_13_n_0 ;
  wire \rgf_c0bus_wb[8]_i_15_n_0 ;
  wire \rgf_c0bus_wb[8]_i_16_n_0 ;
  wire \rgf_c0bus_wb[8]_i_18_n_0 ;
  wire \rgf_c0bus_wb[8]_i_2_n_0 ;
  wire \rgf_c0bus_wb[8]_i_3_n_0 ;
  wire \rgf_c0bus_wb[8]_i_4_n_0 ;
  wire \rgf_c0bus_wb[8]_i_5_n_0 ;
  wire \rgf_c0bus_wb[9]_i_10_n_0 ;
  wire \rgf_c0bus_wb[9]_i_11_n_0 ;
  wire \rgf_c0bus_wb[9]_i_12_n_0 ;
  wire \rgf_c0bus_wb[9]_i_13_n_0 ;
  wire \rgf_c0bus_wb[9]_i_14_n_0 ;
  wire \rgf_c0bus_wb[9]_i_15_n_0 ;
  wire \rgf_c0bus_wb[9]_i_16_n_0 ;
  wire \rgf_c0bus_wb[9]_i_18_n_0 ;
  wire \rgf_c0bus_wb[9]_i_2_n_0 ;
  wire \rgf_c0bus_wb[9]_i_3_0 ;
  wire \rgf_c0bus_wb[9]_i_3_1 ;
  wire \rgf_c0bus_wb[9]_i_3_n_0 ;
  wire \rgf_c0bus_wb[9]_i_4_n_0 ;
  wire \rgf_c0bus_wb[9]_i_5_n_0 ;
  wire \rgf_c0bus_wb[9]_i_9_n_0 ;
  wire \rgf_c0bus_wb_reg[0] ;
  wire \rgf_c0bus_wb_reg[0]_i_4_n_0 ;
  wire \rgf_c0bus_wb_reg[10] ;
  wire \rgf_c0bus_wb_reg[10]_0 ;
  wire \rgf_c0bus_wb_reg[10]_1 ;
  wire \rgf_c0bus_wb_reg[10]_2 ;
  wire \rgf_c0bus_wb_reg[10]_3 ;
  wire \rgf_c0bus_wb_reg[10]_i_17_0 ;
  wire \rgf_c0bus_wb_reg[10]_i_17_1 ;
  wire \rgf_c0bus_wb_reg[10]_i_17_2 ;
  wire \rgf_c0bus_wb_reg[10]_i_17_n_0 ;
  wire \rgf_c0bus_wb_reg[11] ;
  wire [3:0]\rgf_c0bus_wb_reg[11]_0 ;
  wire \rgf_c0bus_wb_reg[11]_1 ;
  wire \rgf_c0bus_wb_reg[11]_2 ;
  wire \rgf_c0bus_wb_reg[11]_3 ;
  wire \rgf_c0bus_wb_reg[12] ;
  wire \rgf_c0bus_wb_reg[12]_0 ;
  wire \rgf_c0bus_wb_reg[13] ;
  wire \rgf_c0bus_wb_reg[13]_0 ;
  wire \rgf_c0bus_wb_reg[13]_1 ;
  wire \rgf_c0bus_wb_reg[14] ;
  wire \rgf_c0bus_wb_reg[14]_0 ;
  wire [3:0]\rgf_c0bus_wb_reg[15] ;
  wire \rgf_c0bus_wb_reg[15]_0 ;
  wire \rgf_c0bus_wb_reg[15]_i_3_n_0 ;
  wire \rgf_c0bus_wb_reg[1] ;
  wire \rgf_c0bus_wb_reg[1]_0 ;
  wire \rgf_c0bus_wb_reg[2] ;
  wire \rgf_c0bus_wb_reg[2]_0 ;
  wire \rgf_c0bus_wb_reg[2]_1 ;
  wire [3:0]\rgf_c0bus_wb_reg[3] ;
  wire \rgf_c0bus_wb_reg[3]_0 ;
  wire \rgf_c0bus_wb_reg[4] ;
  wire \rgf_c0bus_wb_reg[4]_0 ;
  wire \rgf_c0bus_wb_reg[4]_1 ;
  wire \rgf_c0bus_wb_reg[4]_2 ;
  wire \rgf_c0bus_wb_reg[5] ;
  wire \rgf_c0bus_wb_reg[5]_0 ;
  wire \rgf_c0bus_wb_reg[5]_1 ;
  wire \rgf_c0bus_wb_reg[6] ;
  wire \rgf_c0bus_wb_reg[6]_0 ;
  wire \rgf_c0bus_wb_reg[6]_1 ;
  wire \rgf_c0bus_wb_reg[7] ;
  wire [3:0]\rgf_c0bus_wb_reg[7]_0 ;
  wire \rgf_c0bus_wb_reg[7]_1 ;
  wire \rgf_c0bus_wb_reg[7]_2 ;
  wire \rgf_c0bus_wb_reg[7]_3 ;
  wire \rgf_c0bus_wb_reg[7]_i_11_n_0 ;
  wire \rgf_c0bus_wb_reg[8] ;
  wire \rgf_c0bus_wb_reg[8]_0 ;
  wire \rgf_c0bus_wb_reg[8]_1 ;
  wire \rgf_c0bus_wb_reg[8]_2 ;
  wire \rgf_c0bus_wb_reg[8]_3 ;
  wire \rgf_c0bus_wb_reg[8]_4 ;
  wire \rgf_c0bus_wb_reg[9] ;
  wire \rgf_c0bus_wb_reg[9]_0 ;
  wire \rgf_c0bus_wb_reg[9]_1 ;
  wire \rgf_c0bus_wb_reg[9]_2 ;
  wire \rgf_c1bus_wb[0]_i_10_n_0 ;
  wire \rgf_c1bus_wb[0]_i_11_n_0 ;
  wire \rgf_c1bus_wb[0]_i_13_n_0 ;
  wire \rgf_c1bus_wb[0]_i_14_n_0 ;
  wire \rgf_c1bus_wb[0]_i_15_n_0 ;
  wire \rgf_c1bus_wb[0]_i_16_0 ;
  wire \rgf_c1bus_wb[0]_i_16_n_0 ;
  wire \rgf_c1bus_wb[0]_i_17_n_0 ;
  wire \rgf_c1bus_wb[0]_i_18_n_0 ;
  wire \rgf_c1bus_wb[0]_i_19_n_0 ;
  wire \rgf_c1bus_wb[0]_i_20_n_0 ;
  wire \rgf_c1bus_wb[0]_i_21_n_0 ;
  wire \rgf_c1bus_wb[0]_i_22_n_0 ;
  wire \rgf_c1bus_wb[0]_i_23_n_0 ;
  wire \rgf_c1bus_wb[0]_i_24_n_0 ;
  wire \rgf_c1bus_wb[0]_i_25_n_0 ;
  wire \rgf_c1bus_wb[0]_i_26_n_0 ;
  wire \rgf_c1bus_wb[0]_i_27_n_0 ;
  wire \rgf_c1bus_wb[0]_i_2_n_0 ;
  wire \rgf_c1bus_wb[0]_i_3_n_0 ;
  wire \rgf_c1bus_wb[0]_i_4_0 ;
  wire \rgf_c1bus_wb[0]_i_4_1 ;
  wire \rgf_c1bus_wb[0]_i_4_n_0 ;
  wire \rgf_c1bus_wb[0]_i_6_n_0 ;
  wire \rgf_c1bus_wb[0]_i_7_n_0 ;
  wire \rgf_c1bus_wb[0]_i_9_n_0 ;
  wire \rgf_c1bus_wb[10]_i_12_n_0 ;
  wire \rgf_c1bus_wb[10]_i_13_n_0 ;
  wire \rgf_c1bus_wb[10]_i_14_n_0 ;
  wire \rgf_c1bus_wb[10]_i_16_n_0 ;
  wire \rgf_c1bus_wb[10]_i_17_n_0 ;
  wire \rgf_c1bus_wb[10]_i_18_n_0 ;
  wire \rgf_c1bus_wb[10]_i_3_n_0 ;
  wire \rgf_c1bus_wb[10]_i_4_n_0 ;
  wire \rgf_c1bus_wb[10]_i_5_n_0 ;
  wire \rgf_c1bus_wb[10]_i_9_n_0 ;
  wire \rgf_c1bus_wb[11]_i_11_n_0 ;
  wire \rgf_c1bus_wb[11]_i_15_n_0 ;
  wire \rgf_c1bus_wb[11]_i_16_n_0 ;
  wire \rgf_c1bus_wb[11]_i_17_n_0 ;
  wire \rgf_c1bus_wb[11]_i_18_n_0 ;
  wire \rgf_c1bus_wb[11]_i_19_n_0 ;
  wire \rgf_c1bus_wb[11]_i_20_n_0 ;
  wire \rgf_c1bus_wb[11]_i_21_n_0 ;
  wire \rgf_c1bus_wb[11]_i_22_n_0 ;
  wire \rgf_c1bus_wb[11]_i_2_n_0 ;
  wire \rgf_c1bus_wb[11]_i_3_0 ;
  wire \rgf_c1bus_wb[11]_i_3_n_0 ;
  wire \rgf_c1bus_wb[11]_i_4_n_0 ;
  wire \rgf_c1bus_wb[11]_i_5_n_0 ;
  wire \rgf_c1bus_wb[11]_i_6_0 ;
  wire \rgf_c1bus_wb[11]_i_6_n_0 ;
  wire \rgf_c1bus_wb[11]_i_8_n_0 ;
  wire \rgf_c1bus_wb[12]_i_10_n_0 ;
  wire \rgf_c1bus_wb[12]_i_12_n_0 ;
  wire \rgf_c1bus_wb[12]_i_13_n_0 ;
  wire \rgf_c1bus_wb[12]_i_14_n_0 ;
  wire \rgf_c1bus_wb[12]_i_22_n_0 ;
  wire \rgf_c1bus_wb[12]_i_23_n_0 ;
  wire \rgf_c1bus_wb[12]_i_24_n_0 ;
  wire \rgf_c1bus_wb[12]_i_25_n_0 ;
  wire \rgf_c1bus_wb[12]_i_2_n_0 ;
  wire \rgf_c1bus_wb[12]_i_3_n_0 ;
  wire \rgf_c1bus_wb[12]_i_4_n_0 ;
  wire \rgf_c1bus_wb[12]_i_5_n_0 ;
  wire \rgf_c1bus_wb[12]_i_6_n_0 ;
  wire \rgf_c1bus_wb[12]_i_8_n_0 ;
  wire \rgf_c1bus_wb[12]_i_9_n_0 ;
  wire \rgf_c1bus_wb[13]_i_11_n_0 ;
  wire \rgf_c1bus_wb[13]_i_12_n_0 ;
  wire \rgf_c1bus_wb[13]_i_13_n_0 ;
  wire \rgf_c1bus_wb[13]_i_14_n_0 ;
  wire \rgf_c1bus_wb[13]_i_15_n_0 ;
  wire \rgf_c1bus_wb[13]_i_17_n_0 ;
  wire \rgf_c1bus_wb[13]_i_23_n_0 ;
  wire \rgf_c1bus_wb[13]_i_2_0 ;
  wire \rgf_c1bus_wb[13]_i_2_n_0 ;
  wire \rgf_c1bus_wb[13]_i_3_n_0 ;
  wire \rgf_c1bus_wb[13]_i_5_0 ;
  wire \rgf_c1bus_wb[13]_i_5_n_0 ;
  wire \rgf_c1bus_wb[13]_i_7_n_0 ;
  wire \rgf_c1bus_wb[14]_i_11_n_0 ;
  wire \rgf_c1bus_wb[14]_i_12_n_0 ;
  wire \rgf_c1bus_wb[14]_i_13_n_0 ;
  wire \rgf_c1bus_wb[14]_i_14_n_0 ;
  wire \rgf_c1bus_wb[14]_i_15_n_0 ;
  wire \rgf_c1bus_wb[14]_i_19_n_0 ;
  wire \rgf_c1bus_wb[14]_i_21_n_0 ;
  wire \rgf_c1bus_wb[14]_i_22_n_0 ;
  wire \rgf_c1bus_wb[14]_i_23_n_0 ;
  wire \rgf_c1bus_wb[14]_i_24_n_0 ;
  wire \rgf_c1bus_wb[14]_i_25_n_0 ;
  wire \rgf_c1bus_wb[14]_i_26_n_0 ;
  wire \rgf_c1bus_wb[14]_i_27_n_0 ;
  wire \rgf_c1bus_wb[14]_i_28_0 ;
  wire \rgf_c1bus_wb[14]_i_28_1 ;
  wire \rgf_c1bus_wb[14]_i_28_2 ;
  wire \rgf_c1bus_wb[14]_i_34_n_0 ;
  wire \rgf_c1bus_wb[14]_i_35_n_0 ;
  wire \rgf_c1bus_wb[14]_i_36_n_0 ;
  wire \rgf_c1bus_wb[14]_i_37_n_0 ;
  wire \rgf_c1bus_wb[14]_i_38_n_0 ;
  wire \rgf_c1bus_wb[14]_i_39_n_0 ;
  wire \rgf_c1bus_wb[14]_i_3_0 ;
  wire \rgf_c1bus_wb[14]_i_3_1 ;
  wire \rgf_c1bus_wb[14]_i_3_n_0 ;
  wire \rgf_c1bus_wb[14]_i_40_n_0 ;
  wire \rgf_c1bus_wb[14]_i_41_n_0 ;
  wire \rgf_c1bus_wb[14]_i_42_n_0 ;
  wire \rgf_c1bus_wb[14]_i_43_n_0 ;
  wire \rgf_c1bus_wb[14]_i_44_n_0 ;
  wire \rgf_c1bus_wb[14]_i_45_n_0 ;
  wire \rgf_c1bus_wb[14]_i_46_n_0 ;
  wire \rgf_c1bus_wb[14]_i_47_n_0 ;
  wire \rgf_c1bus_wb[14]_i_48_n_0 ;
  wire \rgf_c1bus_wb[14]_i_49_n_0 ;
  wire \rgf_c1bus_wb[14]_i_4_n_0 ;
  wire \rgf_c1bus_wb[14]_i_50_n_0 ;
  wire \rgf_c1bus_wb[14]_i_51_n_0 ;
  wire \rgf_c1bus_wb[14]_i_52_n_0 ;
  wire \rgf_c1bus_wb[14]_i_53_0 ;
  wire \rgf_c1bus_wb[14]_i_53_n_0 ;
  wire \rgf_c1bus_wb[14]_i_54_n_0 ;
  wire \rgf_c1bus_wb[14]_i_55_n_0 ;
  wire \rgf_c1bus_wb[14]_i_56_n_0 ;
  wire \rgf_c1bus_wb[14]_i_57_n_0 ;
  wire \rgf_c1bus_wb[14]_i_58_n_0 ;
  wire \rgf_c1bus_wb[14]_i_59_n_0 ;
  wire \rgf_c1bus_wb[14]_i_5_n_0 ;
  wire \rgf_c1bus_wb[14]_i_60_n_0 ;
  wire \rgf_c1bus_wb[14]_i_61_n_0 ;
  wire \rgf_c1bus_wb[14]_i_62_n_0 ;
  wire \rgf_c1bus_wb[14]_i_63_n_0 ;
  wire \rgf_c1bus_wb[14]_i_64_n_0 ;
  wire \rgf_c1bus_wb[14]_i_65_n_0 ;
  wire \rgf_c1bus_wb[14]_i_66_n_0 ;
  wire \rgf_c1bus_wb[14]_i_67_n_0 ;
  wire \rgf_c1bus_wb[14]_i_68_n_0 ;
  wire \rgf_c1bus_wb[14]_i_6_n_0 ;
  wire \rgf_c1bus_wb[14]_i_7_n_0 ;
  wire \rgf_c1bus_wb[14]_i_8_n_0 ;
  wire \rgf_c1bus_wb[14]_i_9_n_0 ;
  wire \rgf_c1bus_wb[15]_i_10_0 ;
  wire \rgf_c1bus_wb[15]_i_10_n_0 ;
  wire \rgf_c1bus_wb[15]_i_11_n_0 ;
  wire \rgf_c1bus_wb[15]_i_12_n_0 ;
  wire \rgf_c1bus_wb[15]_i_13_n_0 ;
  wire \rgf_c1bus_wb[15]_i_14_0 ;
  wire \rgf_c1bus_wb[15]_i_14_1 ;
  wire \rgf_c1bus_wb[15]_i_16_n_0 ;
  wire \rgf_c1bus_wb[15]_i_17_n_0 ;
  wire \rgf_c1bus_wb[15]_i_19_n_0 ;
  wire \rgf_c1bus_wb[15]_i_23_n_0 ;
  wire \rgf_c1bus_wb[15]_i_24_n_0 ;
  wire \rgf_c1bus_wb[15]_i_3_n_0 ;
  wire \rgf_c1bus_wb[15]_i_4_0 ;
  wire \rgf_c1bus_wb[15]_i_4_n_0 ;
  wire \rgf_c1bus_wb[15]_i_5_n_0 ;
  wire \rgf_c1bus_wb[15]_i_7_n_0 ;
  wire \rgf_c1bus_wb[15]_i_9_n_0 ;
  wire \rgf_c1bus_wb[1]_i_10_n_0 ;
  wire \rgf_c1bus_wb[1]_i_12_n_0 ;
  wire \rgf_c1bus_wb[1]_i_15_n_0 ;
  wire \rgf_c1bus_wb[1]_i_17_n_0 ;
  wire \rgf_c1bus_wb[1]_i_18_n_0 ;
  wire \rgf_c1bus_wb[1]_i_19_n_0 ;
  wire \rgf_c1bus_wb[1]_i_2_0 ;
  wire \rgf_c1bus_wb[1]_i_2_1 ;
  wire \rgf_c1bus_wb[1]_i_2_n_0 ;
  wire \rgf_c1bus_wb[1]_i_3_n_0 ;
  wire \rgf_c1bus_wb[1]_i_5_n_0 ;
  wire \rgf_c1bus_wb[1]_i_6_n_0 ;
  wire \rgf_c1bus_wb[1]_i_7_n_0 ;
  wire \rgf_c1bus_wb[1]_i_8_n_0 ;
  wire \rgf_c1bus_wb[1]_i_9_n_0 ;
  wire \rgf_c1bus_wb[2]_i_10_n_0 ;
  wire \rgf_c1bus_wb[2]_i_11_n_0 ;
  wire \rgf_c1bus_wb[2]_i_12_n_0 ;
  wire \rgf_c1bus_wb[2]_i_14_n_0 ;
  wire \rgf_c1bus_wb[2]_i_15_n_0 ;
  wire \rgf_c1bus_wb[2]_i_16_n_0 ;
  wire \rgf_c1bus_wb[2]_i_17_n_0 ;
  wire \rgf_c1bus_wb[2]_i_2_n_0 ;
  wire \rgf_c1bus_wb[2]_i_3_n_0 ;
  wire \rgf_c1bus_wb[2]_i_5_n_0 ;
  wire \rgf_c1bus_wb[2]_i_7_n_0 ;
  wire \rgf_c1bus_wb[2]_i_8_n_0 ;
  wire \rgf_c1bus_wb[2]_i_9_n_0 ;
  wire \rgf_c1bus_wb[3]_i_10_n_0 ;
  wire \rgf_c1bus_wb[3]_i_11_n_0 ;
  wire \rgf_c1bus_wb[3]_i_12_n_0 ;
  wire \rgf_c1bus_wb[3]_i_13_n_0 ;
  wire \rgf_c1bus_wb[3]_i_3_n_0 ;
  wire \rgf_c1bus_wb[3]_i_4_n_0 ;
  wire \rgf_c1bus_wb[3]_i_5_n_0 ;
  wire \rgf_c1bus_wb[3]_i_7_n_0 ;
  wire \rgf_c1bus_wb[3]_i_8_n_0 ;
  wire \rgf_c1bus_wb[3]_i_9_n_0 ;
  wire \rgf_c1bus_wb[4]_i_10_n_0 ;
  wire \rgf_c1bus_wb[4]_i_11_0 ;
  wire \rgf_c1bus_wb[4]_i_11_1 ;
  wire \rgf_c1bus_wb[4]_i_11_2 ;
  wire \rgf_c1bus_wb[4]_i_11_n_0 ;
  wire \rgf_c1bus_wb[4]_i_13_n_0 ;
  wire \rgf_c1bus_wb[4]_i_14_n_0 ;
  wire \rgf_c1bus_wb[4]_i_15_n_0 ;
  wire \rgf_c1bus_wb[4]_i_16_n_0 ;
  wire \rgf_c1bus_wb[4]_i_22_n_0 ;
  wire \rgf_c1bus_wb[4]_i_2_n_0 ;
  wire \rgf_c1bus_wb[4]_i_4_0 ;
  wire \rgf_c1bus_wb[4]_i_4_1 ;
  wire \rgf_c1bus_wb[4]_i_4_2 ;
  wire \rgf_c1bus_wb[4]_i_4_3 ;
  wire \rgf_c1bus_wb[4]_i_4_n_0 ;
  wire \rgf_c1bus_wb[4]_i_5_n_0 ;
  wire \rgf_c1bus_wb[5]_i_10_n_0 ;
  wire \rgf_c1bus_wb[5]_i_12_n_0 ;
  wire \rgf_c1bus_wb[5]_i_2_n_0 ;
  wire \rgf_c1bus_wb[5]_i_3_n_0 ;
  wire \rgf_c1bus_wb[5]_i_5_n_0 ;
  wire \rgf_c1bus_wb[5]_i_6_n_0 ;
  wire \rgf_c1bus_wb[5]_i_7_n_0 ;
  wire \rgf_c1bus_wb[5]_i_8_n_0 ;
  wire \rgf_c1bus_wb[5]_i_9_0 ;
  wire \rgf_c1bus_wb[5]_i_9_1 ;
  wire \rgf_c1bus_wb[5]_i_9_2 ;
  wire \rgf_c1bus_wb[6]_i_10_n_0 ;
  wire \rgf_c1bus_wb[6]_i_11_n_0 ;
  wire \rgf_c1bus_wb[6]_i_12_n_0 ;
  wire \rgf_c1bus_wb[6]_i_15_n_0 ;
  wire \rgf_c1bus_wb[6]_i_16_n_0 ;
  wire \rgf_c1bus_wb[6]_i_2_n_0 ;
  wire \rgf_c1bus_wb[6]_i_3_n_0 ;
  wire \rgf_c1bus_wb[6]_i_5_n_0 ;
  wire \rgf_c1bus_wb[6]_i_7_n_0 ;
  wire \rgf_c1bus_wb[6]_i_8_n_0 ;
  wire \rgf_c1bus_wb[6]_i_9_n_0 ;
  wire \rgf_c1bus_wb[7]_i_11_n_0 ;
  wire \rgf_c1bus_wb[7]_i_12_n_0 ;
  wire \rgf_c1bus_wb[7]_i_13_n_0 ;
  wire \rgf_c1bus_wb[7]_i_15_n_0 ;
  wire \rgf_c1bus_wb[7]_i_16_n_0 ;
  wire \rgf_c1bus_wb[7]_i_17_n_0 ;
  wire \rgf_c1bus_wb[7]_i_18_n_0 ;
  wire \rgf_c1bus_wb[7]_i_2_n_0 ;
  wire \rgf_c1bus_wb[7]_i_5_n_0 ;
  wire \rgf_c1bus_wb[7]_i_6_n_0 ;
  wire \rgf_c1bus_wb[7]_i_9_n_0 ;
  wire \rgf_c1bus_wb[8]_i_12_n_0 ;
  wire \rgf_c1bus_wb[8]_i_13_n_0 ;
  wire \rgf_c1bus_wb[8]_i_14_n_0 ;
  wire \rgf_c1bus_wb[8]_i_15_n_0 ;
  wire \rgf_c1bus_wb[8]_i_16_n_0 ;
  wire \rgf_c1bus_wb[8]_i_2_n_0 ;
  wire \rgf_c1bus_wb[8]_i_3_n_0 ;
  wire \rgf_c1bus_wb[8]_i_5_n_0 ;
  wire \rgf_c1bus_wb[8]_i_6_n_0 ;
  wire \rgf_c1bus_wb[8]_i_7_n_0 ;
  wire \rgf_c1bus_wb[8]_i_9_n_0 ;
  wire \rgf_c1bus_wb[9]_i_10_n_0 ;
  wire \rgf_c1bus_wb[9]_i_11_n_0 ;
  wire \rgf_c1bus_wb[9]_i_12_n_0 ;
  wire \rgf_c1bus_wb[9]_i_13_n_0 ;
  wire \rgf_c1bus_wb[9]_i_14_n_0 ;
  wire \rgf_c1bus_wb[9]_i_15_n_0 ;
  wire \rgf_c1bus_wb[9]_i_18_n_0 ;
  wire \rgf_c1bus_wb[9]_i_19_n_0 ;
  wire \rgf_c1bus_wb[9]_i_2_n_0 ;
  wire \rgf_c1bus_wb[9]_i_3_0 ;
  wire \rgf_c1bus_wb[9]_i_3_1 ;
  wire \rgf_c1bus_wb[9]_i_3_2 ;
  wire \rgf_c1bus_wb[9]_i_3_n_0 ;
  wire \rgf_c1bus_wb[9]_i_7_n_0 ;
  wire \rgf_c1bus_wb[9]_i_8_n_0 ;
  wire \rgf_c1bus_wb[9]_i_9_n_0 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire \rgf_c1bus_wb_reg[10] ;
  wire \rgf_c1bus_wb_reg[10]_0 ;
  wire [1:0]\rgf_c1bus_wb_reg[11] ;
  wire \rgf_c1bus_wb_reg[11]_0 ;
  wire \rgf_c1bus_wb_reg[11]_i_7_n_0 ;
  wire \rgf_c1bus_wb_reg[12] ;
  wire \rgf_c1bus_wb_reg[12]_0 ;
  wire \rgf_c1bus_wb_reg[12]_1 ;
  wire \rgf_c1bus_wb_reg[12]_i_15_n_0 ;
  wire \rgf_c1bus_wb_reg[13] ;
  wire \rgf_c1bus_wb_reg[13]_0 ;
  wire \rgf_c1bus_wb_reg[13]_1 ;
  wire \rgf_c1bus_wb_reg[13]_2 ;
  wire \rgf_c1bus_wb_reg[13]_3 ;
  wire \rgf_c1bus_wb_reg[13]_4 ;
  wire \rgf_c1bus_wb_reg[13]_5 ;
  wire \rgf_c1bus_wb_reg[13]_6 ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire \rgf_c1bus_wb_reg[14]_0 ;
  wire \rgf_c1bus_wb_reg[14]_1 ;
  wire \rgf_c1bus_wb_reg[14]_2 ;
  wire \rgf_c1bus_wb_reg[14]_3 ;
  wire [1:0]\rgf_c1bus_wb_reg[15] ;
  wire \rgf_c1bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb_reg[15]_1 ;
  wire \rgf_c1bus_wb_reg[1] ;
  wire \rgf_c1bus_wb_reg[1]_0 ;
  wire \rgf_c1bus_wb_reg[1]_1 ;
  wire \rgf_c1bus_wb_reg[2] ;
  wire \rgf_c1bus_wb_reg[2]_0 ;
  wire \rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[3]_0 ;
  wire \rgf_c1bus_wb_reg[3]_1 ;
  wire [2:0]\rgf_c1bus_wb_reg[3]_2 ;
  wire \rgf_c1bus_wb_reg[3]_3 ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[4]_0 ;
  wire \rgf_c1bus_wb_reg[4]_1 ;
  wire \rgf_c1bus_wb_reg[4]_2 ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[5]_0 ;
  wire \rgf_c1bus_wb_reg[6] ;
  wire \rgf_c1bus_wb_reg[6]_0 ;
  wire \rgf_c1bus_wb_reg[6]_1 ;
  wire \rgf_c1bus_wb_reg[6]_2 ;
  wire \rgf_c1bus_wb_reg[6]_3 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire \rgf_c1bus_wb_reg[7]_0 ;
  wire [2:0]\rgf_c1bus_wb_reg[7]_1 ;
  wire \rgf_c1bus_wb_reg[7]_2 ;
  wire \rgf_c1bus_wb_reg[7]_3 ;
  wire \rgf_c1bus_wb_reg[8] ;
  wire \rgf_c1bus_wb_reg[8]_0 ;
  wire \rgf_c1bus_wb_reg[8]_1 ;
  wire \rgf_c1bus_wb_reg[8]_2 ;
  wire \rgf_c1bus_wb_reg[9] ;
  wire \rgf_c1bus_wb_reg[9]_0 ;
  wire \rgf_c1bus_wb_reg[9]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_33_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_5_0 ;
  wire \rgf_selc0_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_28_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_29_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_9_n_0 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[0] ;
  wire \rgf_selc0_rn_wb_reg[0]_0 ;
  wire \rgf_selc0_rn_wb_reg[0]_1 ;
  wire rgf_selc0_stat;
  wire \rgf_selc0_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_wb[1]_i_26_n_0 ;
  wire \rgf_selc0_wb[1]_i_28_n_0 ;
  wire \rgf_selc0_wb[1]_i_29_n_0 ;
  wire \rgf_selc0_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_wb[1]_i_30_n_0 ;
  wire \rgf_selc0_wb[1]_i_31_n_0 ;
  wire \rgf_selc0_wb[1]_i_32_n_0 ;
  wire \rgf_selc0_wb[1]_i_33_n_0 ;
  wire \rgf_selc0_wb[1]_i_34_n_0 ;
  wire \rgf_selc0_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_wb[1]_i_4_0 ;
  wire \rgf_selc0_wb[1]_i_4_1 ;
  wire \rgf_selc0_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_1 ;
  wire \rgf_selc1_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb_reg[0] ;
  wire \rgf_selc1_rn_wb_reg[2] ;
  wire rgf_selc1_stat;
  wire [15:0]rgf_selc1_stat_reg;
  wire [15:0]rgf_selc1_stat_reg_0;
  wire [15:0]rgf_selc1_stat_reg_1;
  wire [15:0]rgf_selc1_stat_reg_10;
  wire [15:0]rgf_selc1_stat_reg_11;
  wire [15:0]rgf_selc1_stat_reg_12;
  wire [15:0]rgf_selc1_stat_reg_13;
  wire [15:0]rgf_selc1_stat_reg_14;
  wire [15:0]rgf_selc1_stat_reg_15;
  wire [15:0]rgf_selc1_stat_reg_16;
  wire [15:0]rgf_selc1_stat_reg_17;
  wire [15:0]rgf_selc1_stat_reg_18;
  wire [15:0]rgf_selc1_stat_reg_19;
  wire [15:0]rgf_selc1_stat_reg_2;
  wire [15:0]rgf_selc1_stat_reg_20;
  wire [15:0]rgf_selc1_stat_reg_21;
  wire [15:0]rgf_selc1_stat_reg_22;
  wire [15:0]rgf_selc1_stat_reg_23;
  wire [15:0]rgf_selc1_stat_reg_24;
  wire [15:0]rgf_selc1_stat_reg_25;
  wire [15:0]rgf_selc1_stat_reg_26;
  wire [15:0]rgf_selc1_stat_reg_27;
  wire [15:0]rgf_selc1_stat_reg_28;
  wire [15:0]rgf_selc1_stat_reg_29;
  wire [15:0]rgf_selc1_stat_reg_3;
  wire [15:0]rgf_selc1_stat_reg_30;
  wire [15:0]rgf_selc1_stat_reg_31;
  wire [15:0]rgf_selc1_stat_reg_4;
  wire [15:0]rgf_selc1_stat_reg_5;
  wire [15:0]rgf_selc1_stat_reg_6;
  wire [15:0]rgf_selc1_stat_reg_7;
  wire [15:0]rgf_selc1_stat_reg_8;
  wire [15:0]rgf_selc1_stat_reg_9;
  wire \rgf_selc1_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_wb[1]_i_26_n_0 ;
  wire \rgf_selc1_wb[1]_i_29_n_0 ;
  wire \rgf_selc1_wb[1]_i_30_n_0 ;
  wire \rgf_selc1_wb[1]_i_31_n_0 ;
  wire \rgf_selc1_wb[1]_i_32_n_0 ;
  wire \rgf_selc1_wb[1]_i_33_n_0 ;
  wire \rgf_selc1_wb[1]_i_34_n_0 ;
  wire \rgf_selc1_wb[1]_i_35_n_0 ;
  wire \rgf_selc1_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_wb[1]_i_5_0 ;
  wire \rgf_selc1_wb[1]_i_5_1 ;
  wire \rgf_selc1_wb[1]_i_5_2 ;
  wire \rgf_selc1_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_wb_reg[0] ;
  wire [2:0]\rgf_selc1_wb_reg[1] ;
  wire \rgf_selc1_wb_reg[1]_0 ;
  wire \rgf_selc1_wb_reg[1]_i_21_n_0 ;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_fl;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_10;
  wire rst_n_fl_reg_11;
  wire rst_n_fl_reg_12;
  wire rst_n_fl_reg_2;
  wire rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire rst_n_fl_reg_5;
  wire rst_n_fl_reg_6;
  wire rst_n_fl_reg_7;
  wire rst_n_fl_reg_8;
  wire rst_n_fl_reg_9;
  wire \sp[0]_i_2_n_0 ;
  wire \sp[15]_i_10_n_0 ;
  wire \sp[15]_i_11_n_0 ;
  wire \sp[15]_i_13_n_0 ;
  wire \sp[15]_i_14_n_0 ;
  wire \sp[15]_i_15_n_0 ;
  wire \sp[15]_i_16_n_0 ;
  wire \sp[15]_i_17_n_0 ;
  wire \sp[15]_i_18_n_0 ;
  wire \sp[15]_i_19_n_0 ;
  wire \sp[15]_i_2 ;
  wire \sp[15]_i_20_n_0 ;
  wire \sp[15]_i_21_n_0 ;
  wire \sp[15]_i_22_n_0 ;
  wire \sp[15]_i_23_n_0 ;
  wire \sp[15]_i_24_n_0 ;
  wire \sp[15]_i_8_0 ;
  wire \sp[15]_i_9_n_0 ;
  wire [0:0]\sp_reg[0] ;
  wire [0:0]\sp_reg[0]_0 ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire [15:0]\sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[13]_i_11_n_0 ;
  wire \sr[13]_i_12_n_0 ;
  wire \sr[13]_i_13_n_0 ;
  wire \sr[13]_i_14_n_0 ;
  wire \sr[13]_i_15_n_0 ;
  wire [2:0]\sr[13]_i_5 ;
  wire [1:0]\sr[13]_i_5_0 ;
  wire \sr[13]_i_6_n_0 ;
  wire \sr[13]_i_7_n_0 ;
  wire \sr[13]_i_8_n_0 ;
  wire \sr[15]_i_2 ;
  wire \sr[15]_i_9_n_0 ;
  wire \sr[3]_i_3 ;
  wire \sr[3]_i_7_n_0 ;
  wire \sr[4]_i_100_0 ;
  wire \sr[4]_i_100_1 ;
  wire \sr[4]_i_100_2 ;
  wire \sr[4]_i_100_n_0 ;
  wire \sr[4]_i_101_n_0 ;
  wire \sr[4]_i_102_0 ;
  wire \sr[4]_i_102_1 ;
  wire \sr[4]_i_102_2 ;
  wire \sr[4]_i_102_3 ;
  wire \sr[4]_i_102_n_0 ;
  wire \sr[4]_i_103_n_0 ;
  wire \sr[4]_i_104_n_0 ;
  wire \sr[4]_i_106_n_0 ;
  wire \sr[4]_i_107_n_0 ;
  wire \sr[4]_i_108_n_0 ;
  wire \sr[4]_i_109_n_0 ;
  wire \sr[4]_i_10_0 ;
  wire \sr[4]_i_10_1 ;
  wire \sr[4]_i_10_2 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_110_n_0 ;
  wire \sr[4]_i_111_0 ;
  wire \sr[4]_i_111_n_0 ;
  wire \sr[4]_i_112_n_0 ;
  wire \sr[4]_i_113_n_0 ;
  wire \sr[4]_i_114_n_0 ;
  wire \sr[4]_i_116_n_0 ;
  wire \sr[4]_i_117_n_0 ;
  wire \sr[4]_i_118_n_0 ;
  wire \sr[4]_i_119_n_0 ;
  wire \sr[4]_i_11_0 ;
  wire \sr[4]_i_11_n_0 ;
  wire \sr[4]_i_120_n_0 ;
  wire \sr[4]_i_121_n_0 ;
  wire \sr[4]_i_124_n_0 ;
  wire \sr[4]_i_125_n_0 ;
  wire \sr[4]_i_126_n_0 ;
  wire \sr[4]_i_127_0 ;
  wire \sr[4]_i_127_1 ;
  wire \sr[4]_i_127_n_0 ;
  wire \sr[4]_i_128 ;
  wire \sr[4]_i_128_0 ;
  wire \sr[4]_i_129_n_0 ;
  wire \sr[4]_i_12_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_134_n_0 ;
  wire \sr[4]_i_136_n_0 ;
  wire \sr[4]_i_137_n_0 ;
  wire \sr[4]_i_139_n_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_140_n_0 ;
  wire \sr[4]_i_141_n_0 ;
  wire \sr[4]_i_143_n_0 ;
  wire \sr[4]_i_144_n_0 ;
  wire \sr[4]_i_145_n_0 ;
  wire \sr[4]_i_147_n_0 ;
  wire \sr[4]_i_149_n_0 ;
  wire \sr[4]_i_14_n_0 ;
  wire \sr[4]_i_150_n_0 ;
  wire \sr[4]_i_151_n_0 ;
  wire \sr[4]_i_153_n_0 ;
  wire \sr[4]_i_157_n_0 ;
  wire \sr[4]_i_158_n_0 ;
  wire \sr[4]_i_15_0 ;
  wire \sr[4]_i_15_n_0 ;
  wire \sr[4]_i_163_n_0 ;
  wire \sr[4]_i_168_n_0 ;
  wire \sr[4]_i_16_0 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_170_n_0 ;
  wire \sr[4]_i_171_n_0 ;
  wire \sr[4]_i_172_n_0 ;
  wire \sr[4]_i_174_n_0 ;
  wire \sr[4]_i_177_n_0 ;
  wire \sr[4]_i_178_n_0 ;
  wire \sr[4]_i_17_0 ;
  wire \sr[4]_i_17_1 ;
  wire \sr[4]_i_17_n_0 ;
  wire \sr[4]_i_185_n_0 ;
  wire \sr[4]_i_18_0 ;
  wire \sr[4]_i_18_1 ;
  wire \sr[4]_i_18_2 ;
  wire \sr[4]_i_18_3 ;
  wire \sr[4]_i_18_n_0 ;
  wire \sr[4]_i_19_n_0 ;
  wire \sr[4]_i_201_n_0 ;
  wire \sr[4]_i_204_n_0 ;
  wire \sr[4]_i_20_0 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_221_n_0 ;
  wire \sr[4]_i_222_n_0 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_25_0 ;
  wire \sr[4]_i_25_n_0 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_0 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_28_0 ;
  wire \sr[4]_i_28_1 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_29_0 ;
  wire \sr[4]_i_29_1 ;
  wire \sr[4]_i_29_2 ;
  wire \sr[4]_i_29_3 ;
  wire \sr[4]_i_29_n_0 ;
  wire \sr[4]_i_30_0 ;
  wire \sr[4]_i_30_1 ;
  wire \sr[4]_i_30_n_0 ;
  wire \sr[4]_i_31_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_33_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_35_0 ;
  wire \sr[4]_i_35_1 ;
  wire \sr[4]_i_35_n_0 ;
  wire \sr[4]_i_36_0 ;
  wire \sr[4]_i_36_1 ;
  wire \sr[4]_i_36_2 ;
  wire \sr[4]_i_36_n_0 ;
  wire \sr[4]_i_37_0 ;
  wire \sr[4]_i_37_n_0 ;
  wire \sr[4]_i_38_n_0 ;
  wire \sr[4]_i_39_0 ;
  wire \sr[4]_i_39_n_0 ;
  wire \sr[4]_i_3_0 ;
  wire \sr[4]_i_40_n_0 ;
  wire \sr[4]_i_41_0 ;
  wire \sr[4]_i_41_n_0 ;
  wire \sr[4]_i_42_n_0 ;
  wire \sr[4]_i_43_0 ;
  wire \sr[4]_i_43_1 ;
  wire \sr[4]_i_43_2 ;
  wire \sr[4]_i_43_n_0 ;
  wire \sr[4]_i_44_0 ;
  wire \sr[4]_i_44_n_0 ;
  wire \sr[4]_i_45_0 ;
  wire \sr[4]_i_45_n_0 ;
  wire \sr[4]_i_46_0 ;
  wire \sr[4]_i_46_1 ;
  wire \sr[4]_i_46_2 ;
  wire \sr[4]_i_46_n_0 ;
  wire \sr[4]_i_48_n_0 ;
  wire \sr[4]_i_49_n_0 ;
  wire \sr[4]_i_50_n_0 ;
  wire \sr[4]_i_51_n_0 ;
  wire \sr[4]_i_52_0 ;
  wire \sr[4]_i_52_n_0 ;
  wire \sr[4]_i_53_0 ;
  wire \sr[4]_i_53_1 ;
  wire \sr[4]_i_53_n_0 ;
  wire \sr[4]_i_54_0 ;
  wire \sr[4]_i_54_1 ;
  wire \sr[4]_i_54_n_0 ;
  wire \sr[4]_i_55_0 ;
  wire \sr[4]_i_55_1 ;
  wire \sr[4]_i_55_2 ;
  wire \sr[4]_i_55_n_0 ;
  wire \sr[4]_i_56_n_0 ;
  wire \sr[4]_i_58_0 ;
  wire \sr[4]_i_58_n_0 ;
  wire \sr[4]_i_59_n_0 ;
  wire \sr[4]_i_60_0 ;
  wire \sr[4]_i_60_1 ;
  wire \sr[4]_i_60_2 ;
  wire \sr[4]_i_60_n_0 ;
  wire \sr[4]_i_61_n_0 ;
  wire \sr[4]_i_62_n_0 ;
  wire \sr[4]_i_63_0 ;
  wire \sr[4]_i_63_1 ;
  wire \sr[4]_i_63_n_0 ;
  wire \sr[4]_i_64_0 ;
  wire \sr[4]_i_64_1 ;
  wire \sr[4]_i_64_n_0 ;
  wire \sr[4]_i_65_0 ;
  wire \sr[4]_i_65_n_0 ;
  wire \sr[4]_i_66_0 ;
  wire \sr[4]_i_66_n_0 ;
  wire \sr[4]_i_67_0 ;
  wire \sr[4]_i_67_n_0 ;
  wire \sr[4]_i_68_0 ;
  wire \sr[4]_i_68_1 ;
  wire \sr[4]_i_68_n_0 ;
  wire \sr[4]_i_69_0 ;
  wire \sr[4]_i_69_n_0 ;
  wire \sr[4]_i_6_0 ;
  wire \sr[4]_i_70_0 ;
  wire \sr[4]_i_70_n_0 ;
  wire \sr[4]_i_71_0 ;
  wire \sr[4]_i_71_n_0 ;
  wire \sr[4]_i_72_0 ;
  wire \sr[4]_i_72_n_0 ;
  wire \sr[4]_i_73_n_0 ;
  wire \sr[4]_i_74_n_0 ;
  wire \sr[4]_i_75_n_0 ;
  wire \sr[4]_i_76_n_0 ;
  wire \sr[4]_i_77_n_0 ;
  wire \sr[4]_i_78_n_0 ;
  wire \sr[4]_i_79_n_0 ;
  wire \sr[4]_i_81_n_0 ;
  wire \sr[4]_i_82_n_0 ;
  wire \sr[4]_i_83_n_0 ;
  wire \sr[4]_i_84_n_0 ;
  wire \sr[4]_i_85_n_0 ;
  wire \sr[4]_i_86_n_0 ;
  wire \sr[4]_i_87_n_0 ;
  wire \sr[4]_i_88_n_0 ;
  wire \sr[4]_i_90_n_0 ;
  wire \sr[4]_i_91 ;
  wire \sr[4]_i_92_n_0 ;
  wire \sr[4]_i_93_n_0 ;
  wire \sr[4]_i_95_n_0 ;
  wire \sr[4]_i_96_n_0 ;
  wire \sr[4]_i_97_n_0 ;
  wire \sr[4]_i_98_0 ;
  wire \sr[4]_i_98_1 ;
  wire \sr[4]_i_98_n_0 ;
  wire \sr[4]_i_99_n_0 ;
  wire \sr[4]_i_9_0 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_10_n_0 ;
  wire \sr[5]_i_7_n_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[5]_i_9_n_0 ;
  wire \sr[6]_i_10_n_0 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_14_n_0 ;
  wire \sr[6]_i_15_n_0 ;
  wire \sr[6]_i_16 ;
  wire \sr[6]_i_16_0 ;
  wire \sr[6]_i_16_1 ;
  wire \sr[6]_i_18_n_0 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_5 ;
  wire [0:0]\sr[6]_i_5_0 ;
  wire \sr[6]_i_6_0 ;
  wire \sr[6]_i_6_1 ;
  wire \sr[6]_i_6_2 ;
  wire \sr[6]_i_6_3 ;
  wire \sr[6]_i_6_n_0 ;
  wire \sr[6]_i_7_n_0 ;
  wire \sr[6]_i_8_n_0 ;
  wire \sr[6]_i_9_0 ;
  wire \sr[6]_i_9_1 ;
  wire \sr[6]_i_9_n_0 ;
  wire \sr_reg[0] ;
  wire \sr_reg[0]_0 ;
  wire \sr_reg[0]_1 ;
  wire \sr_reg[0]_10 ;
  wire \sr_reg[0]_11 ;
  wire \sr_reg[0]_12 ;
  wire \sr_reg[0]_13 ;
  wire \sr_reg[0]_14 ;
  wire \sr_reg[0]_15 ;
  wire \sr_reg[0]_16 ;
  wire \sr_reg[0]_17 ;
  wire \sr_reg[0]_18 ;
  wire \sr_reg[0]_19 ;
  wire \sr_reg[0]_2 ;
  wire \sr_reg[0]_20 ;
  wire \sr_reg[0]_21 ;
  wire \sr_reg[0]_22 ;
  wire \sr_reg[0]_23 ;
  wire \sr_reg[0]_24 ;
  wire \sr_reg[0]_25 ;
  wire \sr_reg[0]_26 ;
  wire \sr_reg[0]_27 ;
  wire \sr_reg[0]_28 ;
  wire \sr_reg[0]_29 ;
  wire \sr_reg[0]_3 ;
  wire \sr_reg[0]_30 ;
  wire \sr_reg[0]_31 ;
  wire \sr_reg[0]_32 ;
  wire \sr_reg[0]_33 ;
  wire \sr_reg[0]_34 ;
  wire \sr_reg[0]_35 ;
  wire [0:0]\sr_reg[0]_36 ;
  wire [0:0]\sr_reg[0]_37 ;
  wire [0:0]\sr_reg[0]_38 ;
  wire [0:0]\sr_reg[0]_39 ;
  wire \sr_reg[0]_4 ;
  wire [0:0]\sr_reg[0]_40 ;
  wire [0:0]\sr_reg[0]_41 ;
  wire [0:0]\sr_reg[0]_42 ;
  wire [0:0]\sr_reg[0]_43 ;
  wire [0:0]\sr_reg[0]_44 ;
  wire [0:0]\sr_reg[0]_45 ;
  wire [0:0]\sr_reg[0]_46 ;
  wire [0:0]\sr_reg[0]_47 ;
  wire [0:0]\sr_reg[0]_48 ;
  wire [0:0]\sr_reg[0]_49 ;
  wire \sr_reg[0]_5 ;
  wire [0:0]\sr_reg[0]_50 ;
  wire [0:0]\sr_reg[0]_51 ;
  wire [0:0]\sr_reg[0]_52 ;
  wire [0:0]\sr_reg[0]_53 ;
  wire [0:0]\sr_reg[0]_54 ;
  wire [0:0]\sr_reg[0]_55 ;
  wire [0:0]\sr_reg[0]_56 ;
  wire [0:0]\sr_reg[0]_57 ;
  wire [0:0]\sr_reg[0]_58 ;
  wire [0:0]\sr_reg[0]_59 ;
  wire \sr_reg[0]_6 ;
  wire \sr_reg[0]_7 ;
  wire \sr_reg[0]_8 ;
  wire \sr_reg[0]_9 ;
  wire [15:0]\sr_reg[15] ;
  wire [15:0]\sr_reg[15]_0 ;
  wire \sr_reg[1] ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[1]_1 ;
  wire \sr_reg[1]_10 ;
  wire \sr_reg[1]_11 ;
  wire \sr_reg[1]_12 ;
  wire \sr_reg[1]_13 ;
  wire [0:0]\sr_reg[1]_14 ;
  wire [0:0]\sr_reg[1]_15 ;
  wire [0:0]\sr_reg[1]_16 ;
  wire [0:0]\sr_reg[1]_17 ;
  wire [0:0]\sr_reg[1]_18 ;
  wire [0:0]\sr_reg[1]_19 ;
  wire \sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_20 ;
  wire [0:0]\sr_reg[1]_21 ;
  wire \sr_reg[1]_3 ;
  wire \sr_reg[1]_4 ;
  wire \sr_reg[1]_5 ;
  wire \sr_reg[1]_6 ;
  wire \sr_reg[1]_7 ;
  wire \sr_reg[1]_8 ;
  wire \sr_reg[1]_9 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire [0:0]\sr_reg[6]_1 ;
  wire \stat[0]_i_10__0_n_0 ;
  wire \stat[0]_i_10__1_n_0 ;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_11__0_n_0 ;
  wire \stat[0]_i_11__1_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12__1_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13__0_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14__0_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15_0 ;
  wire \stat[0]_i_15__0_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16__0_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_17__0_n_0 ;
  wire \stat[0]_i_17_n_0 ;
  wire \stat[0]_i_18__0_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_19__0_n_0 ;
  wire \stat[0]_i_19_n_0 ;
  wire \stat[0]_i_20__0_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21__0_n_0 ;
  wire \stat[0]_i_21_n_0 ;
  wire \stat[0]_i_22__0_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23__0_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24__0_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25__0_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26__0_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_27__0_n_0 ;
  wire \stat[0]_i_27_n_0 ;
  wire \stat[0]_i_28__0_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2__0_n_0 ;
  wire \stat[0]_i_2__1_0 ;
  wire \stat[0]_i_2__1_n_0 ;
  wire \stat[0]_i_30_0 ;
  wire \stat[0]_i_30__0_n_0 ;
  wire \stat[0]_i_30_n_0 ;
  wire \stat[0]_i_31__0_n_0 ;
  wire \stat[0]_i_31_n_0 ;
  wire \stat[0]_i_32__0_n_0 ;
  wire \stat[0]_i_33__0_n_0 ;
  wire \stat[0]_i_33_n_0 ;
  wire \stat[0]_i_34_n_0 ;
  wire \stat[0]_i_3__0_n_0 ;
  wire \stat[0]_i_3__1_n_0 ;
  wire \stat[0]_i_3__2_n_0 ;
  wire \stat[0]_i_4__0_n_0 ;
  wire \stat[0]_i_4__1_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5__0_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7__0_n_0 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8_0 ;
  wire \stat[0]_i_8__0_n_0 ;
  wire \stat[0]_i_8__1_n_0 ;
  wire \stat[0]_i_9__0_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_10__0_n_0 ;
  wire \stat[1]_i_10_n_0 ;
  wire \stat[1]_i_11__0_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_12__0_n_0 ;
  wire \stat[1]_i_12_n_0 ;
  wire \stat[1]_i_13__0_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_14__0_n_0 ;
  wire \stat[1]_i_14_n_0 ;
  wire \stat[1]_i_15_n_0 ;
  wire \stat[1]_i_16_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_2__0_n_0 ;
  wire \stat[1]_i_2__1_n_0 ;
  wire \stat[1]_i_3__0_n_0 ;
  wire \stat[1]_i_3_n_0 ;
  wire \stat[1]_i_4__0_n_0 ;
  wire \stat[1]_i_4__1_n_0 ;
  wire \stat[1]_i_5__0_n_0 ;
  wire \stat[1]_i_5_n_0 ;
  wire \stat[1]_i_6__0_n_0 ;
  wire \stat[1]_i_6_n_0 ;
  wire \stat[1]_i_7__0_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[1]_i_9__0_n_0 ;
  wire \stat[1]_i_9_n_0 ;
  wire \stat[2]_i_10__0_n_0 ;
  wire \stat[2]_i_10_n_0 ;
  wire \stat[2]_i_11_n_0 ;
  wire \stat[2]_i_12__0_n_0 ;
  wire \stat[2]_i_12_n_0 ;
  wire \stat[2]_i_13__0_n_0 ;
  wire \stat[2]_i_13_n_0 ;
  wire \stat[2]_i_14_n_0 ;
  wire \stat[2]_i_15_n_0 ;
  wire \stat[2]_i_2__1 ;
  wire \stat[2]_i_4 ;
  wire \stat[2]_i_4__0_n_0 ;
  wire \stat[2]_i_5__1_n_0 ;
  wire \stat[2]_i_5_n_0 ;
  wire \stat[2]_i_9__0_n_0 ;
  wire \stat[2]_i_9_n_0 ;
  wire \stat_reg[0] ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_12 ;
  wire \stat_reg[0]_13 ;
  wire \stat_reg[0]_14 ;
  wire [0:0]\stat_reg[0]_15 ;
  wire \stat_reg[0]_16 ;
  wire \stat_reg[0]_17 ;
  wire \stat_reg[0]_18 ;
  wire \stat_reg[0]_19 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_20 ;
  wire \stat_reg[0]_21 ;
  wire \stat_reg[0]_22 ;
  wire \stat_reg[0]_23 ;
  wire \stat_reg[0]_24 ;
  wire \stat_reg[0]_25 ;
  wire \stat_reg[0]_26 ;
  wire \stat_reg[0]_27 ;
  wire \stat_reg[0]_28 ;
  wire \stat_reg[0]_29 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_30 ;
  wire \stat_reg[0]_31 ;
  wire \stat_reg[0]_32 ;
  wire \stat_reg[0]_33 ;
  wire \stat_reg[0]_34 ;
  wire \stat_reg[0]_35 ;
  wire \stat_reg[0]_36 ;
  wire \stat_reg[0]_37 ;
  wire \stat_reg[0]_38 ;
  wire \stat_reg[0]_39 ;
  wire [2:0]\stat_reg[0]_4 ;
  wire \stat_reg[0]_40 ;
  wire \stat_reg[0]_41 ;
  wire \stat_reg[0]_42 ;
  wire \stat_reg[0]_43 ;
  wire \stat_reg[0]_44 ;
  wire \stat_reg[0]_45 ;
  wire \stat_reg[0]_46 ;
  wire \stat_reg[0]_47 ;
  wire \stat_reg[0]_48 ;
  wire \stat_reg[0]_49 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_50 ;
  wire \stat_reg[0]_51 ;
  wire \stat_reg[0]_52 ;
  wire \stat_reg[0]_53 ;
  wire \stat_reg[0]_54 ;
  wire \stat_reg[0]_55 ;
  wire [1:0]\stat_reg[0]_56 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire [2:0]\stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire [2:0]\stat_reg[2] ;
  wire [1:0]\stat_reg[2]_0 ;
  wire [2:0]\stat_reg[2]_1 ;
  wire \stat_reg[2]_10 ;
  wire \stat_reg[2]_11 ;
  wire [1:0]\stat_reg[2]_12 ;
  wire \stat_reg[2]_13 ;
  wire \stat_reg[2]_14 ;
  wire \stat_reg[2]_15 ;
  wire \stat_reg[2]_16 ;
  wire \stat_reg[2]_17 ;
  wire \stat_reg[2]_18 ;
  wire [0:0]\stat_reg[2]_19 ;
  wire [1:0]\stat_reg[2]_2 ;
  wire \stat_reg[2]_20 ;
  wire \stat_reg[2]_21 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire \stat_reg[2]_7 ;
  wire \stat_reg[2]_8 ;
  wire \stat_reg[2]_9 ;
  wire tout__1_carry__0;
  wire [3:0]tout__1_carry__0_i_1_0;
  wire [1:0]tout__1_carry__0_i_3__0_0;
  wire [3:0]tout__1_carry__1_i_1_0;
  wire tout__1_carry_i_11_0;
  wire tout__1_carry_i_11_n_0;
  wire tout__1_carry_i_12_n_0;
  wire tout__1_carry_i_13_n_0;
  wire tout__1_carry_i_14_n_0;
  wire tout__1_carry_i_15_n_0;
  wire tout__1_carry_i_16_n_0;
  wire tout__1_carry_i_17_n_0;
  wire tout__1_carry_i_18_n_0;
  wire tout__1_carry_i_19_n_0;
  wire [3:0]tout__1_carry_i_1_0;
  wire [3:0]tout__1_carry_i_1__0_0;
  wire tout__1_carry_i_20_n_0;
  wire tout__1_carry_i_21_n_0;
  wire tout__1_carry_i_22_0;
  wire tout__1_carry_i_22_n_0;
  wire tout__1_carry_i_23_n_0;
  wire tout__1_carry_i_24_n_0;
  wire tout__1_carry_i_25_0;
  wire tout__1_carry_i_25_n_0;
  wire tout__1_carry_i_26_n_0;
  wire tout__1_carry_i_27_n_0;
  wire tout__1_carry_i_28_n_0;
  wire tout__1_carry_i_29_n_0;
  wire tout__1_carry_i_30_n_0;
  wire tout__1_carry_i_31_n_0;
  wire tout__1_carry_i_32_n_0;
  wire tout__1_carry_i_33_n_0;
  wire tout__1_carry_i_34_n_0;
  wire tout__1_carry_i_36_n_0;
  wire tout__1_carry_i_37_n_0;
  wire tout__1_carry_i_9_n_0;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[0]_1 ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[15] ;
  wire [15:0]\tr_reg[15]_0 ;
  wire [15:0]\tr_reg[15]_1 ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[4]_0 ;
  wire \tr_reg[4]_1 ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[0]),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[10]),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[11]),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[12]),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[13]),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[14]),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[15]),
        .O(abus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[1]),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[2]),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[3]),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[4]),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[5]),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[6]),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[7]),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[8]),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(a0bus_0[9]),
        .O(abus_o[9]));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[0]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[0]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[0]),
        .O(\stat_reg[1]_5 [0]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[0]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [0]),
        .O(a1bus_sr[0]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [0]),
        .I5(\iv_reg[15]_0 [0]),
        .O(\tr_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[10]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[10]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[10]),
        .O(badr[9]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[10]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [10]),
        .O(a1bus_sr[10]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [10]),
        .I5(\iv_reg[15]_0 [10]),
        .O(\tr_reg[10] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[11]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[11]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[11]),
        .O(badr[10]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[11]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [11]),
        .O(a1bus_sr[11]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [11]),
        .I5(\iv_reg[15]_0 [11]),
        .O(\tr_reg[11] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[12]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[12]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[12]),
        .O(badr[11]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[12]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [12]),
        .O(a1bus_sr[12]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [12]),
        .I5(\iv_reg[15]_0 [12]),
        .O(\tr_reg[12] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[13]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[13]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[13]),
        .O(badr[12]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[13]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [13]),
        .O(a1bus_sr[13]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [13]),
        .I5(\iv_reg[15]_0 [13]),
        .O(\tr_reg[13] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[14]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[14]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[14]),
        .O(badr[13]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[14]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [14]),
        .O(a1bus_sr[14]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [14]),
        .I5(\iv_reg[15]_0 [14]),
        .O(\tr_reg[14] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[15]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[15]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[15]),
        .O(badr[14]));
  LUT6 #(
    .INIT(64'h5554555554545454)) 
    \badr[15]_INST_0_i_107 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\badr[15]_INST_0_i_187_n_0 ),
        .I2(\badr[15]_INST_0_i_188_n_0 ),
        .I3(\badr[15]_INST_0_i_189_n_0 ),
        .I4(\badr[15]_INST_0_i_190_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0]_0 ),
        .O(\stat_reg[2]_18 ));
  LUT6 #(
    .INIT(64'hFFFFAAFBAAAAAAAA)) 
    \badr[15]_INST_0_i_108 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_192_n_0 ),
        .I2(\badr[15]_INST_0_i_193_n_0 ),
        .I3(\badr[15]_INST_0_i_111_n_0 ),
        .I4(\badr[15]_INST_0_i_194_n_0 ),
        .I5(ctl_fetch0_fl_reg_0),
        .O(ctl_sela0_rn[0]));
  LUT6 #(
    .INIT(64'h0000557F557F557F)) 
    \badr[15]_INST_0_i_109 
       (.I0(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I2(\badr[15]_INST_0_i_195_n_0 ),
        .I3(\badr[15]_INST_0_i_196_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .O(\badr[15]_INST_0_i_109_n_0 ));
  LUT6 #(
    .INIT(64'h00FCFFFFAAAAFFFF)) 
    \badr[15]_INST_0_i_110 
       (.I0(\badr[15]_INST_0_i_197_n_0 ),
        .I1(\badr[15]_INST_0_i_198_n_0 ),
        .I2(ir0[10]),
        .I3(\badr[15]_INST_0_i_199_n_0 ),
        .I4(ir0[12]),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_110_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \badr[15]_INST_0_i_111 
       (.I0(ir0[15]),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .O(\badr[15]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'h4440FFFF44404440)) 
    \badr[15]_INST_0_i_112 
       (.I0(\badr[15]_INST_0_i_200_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[11]),
        .I3(\bcmd[2]_INST_0_i_9_n_0 ),
        .I4(\fadr[15]_INST_0_i_11_n_0 ),
        .I5(\badr[15]_INST_0_i_201_n_0 ),
        .O(\badr[15]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'h8A888A8A8A888A88)) 
    \badr[15]_INST_0_i_113 
       (.I0(\stat_reg[0]_50 ),
        .I1(\badr[15]_INST_0_i_202_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I3(\badr[15]_INST_0_i_203_n_0 ),
        .I4(\badr[15]_INST_0_i_204_n_0 ),
        .I5(\badr[15]_INST_0_i_205_n_0 ),
        .O(ctl_sela0));
  LUT6 #(
    .INIT(64'h5455545454555455)) 
    \badr[15]_INST_0_i_114 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\badr[15]_INST_0_i_206_n_0 ),
        .I2(\badr[15]_INST_0_i_207_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_10_n_0 ),
        .I4(\badr[15]_INST_0_i_208_n_0 ),
        .I5(\badr[15]_INST_0_i_209_n_0 ),
        .O(\stat_reg[2]_20 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \badr[15]_INST_0_i_117 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\stat_reg[2]_18 ),
        .O(a0bus_sel_0[0]));
  LUT5 #(
    .INIT(32'h80000000)) 
    \badr[15]_INST_0_i_118 
       (.I0(ctl_sela0_rn[1]),
        .I1(\stat_reg[2]_20 ),
        .I2(ctl_sela0),
        .I3(ctl_sela0_rn[0]),
        .I4(\stat_reg[2]_18 ),
        .O(a0bus_sel_0[3]));
  LUT6 #(
    .INIT(64'hFFFF4044FFFFFFFF)) 
    \badr[15]_INST_0_i_139 
       (.I0(\badr[15]_INST_0_i_78_n_0 ),
        .I1(\badr[15]_INST_0_i_77_n_0 ),
        .I2(\badr[15]_INST_0_i_76_n_0 ),
        .I3(\badr[15]_INST_0_i_224_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(ctl_sela1),
        .O(\badr[15]_INST_0_i_139_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[15]_INST_0_i_14 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\badr[15]_INST_0_i_26_n_0 ),
        .O(a1bus_sel_cr[3]));
  LUT6 #(
    .INIT(64'h55454444FFFFFFFF)) 
    \badr[15]_INST_0_i_140 
       (.I0(\badr[15]_INST_0_i_84_n_0 ),
        .I1(\bcmd[2]_INST_0_i_7_n_0 ),
        .I2(\bcmd[2]_INST_0_i_5_n_0 ),
        .I3(\badr[15]_INST_0_i_225_n_0 ),
        .I4(\stat[1]_i_6__0_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_53_0 ),
        .O(\badr[15]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'h0000000045440000)) 
    \badr[15]_INST_0_i_141 
       (.I0(\badr[15]_INST_0_i_139_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(\badr[15]_INST_0_i_83_n_0 ),
        .I3(\badr[15]_INST_0_i_140_n_0 ),
        .I4(\badr[15]_INST_0_i_26_n_0 ),
        .I5(\stat_reg[2]_16 ),
        .O(a1bus_sel_0[0]));
  LUT6 #(
    .INIT(64'hFFFDFFDEFFFF9FFC)) 
    \badr[15]_INST_0_i_142 
       (.I0(ir1[7]),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_142_n_0 ));
  LUT5 #(
    .INIT(32'h0000F08F)) 
    \badr[15]_INST_0_i_143 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_143_n_0 ));
  LUT6 #(
    .INIT(64'h0C00EFFF000033FF)) 
    \badr[15]_INST_0_i_144 
       (.I0(ir1[7]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(ir1[8]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_144_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_146 
       (.I0(ir1[13]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_146_n_0 ));
  LUT5 #(
    .INIT(32'hFFBAEEBA)) 
    \badr[15]_INST_0_i_147 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[15]),
        .I2(\sr_reg[15]_0 [6]),
        .I3(ir1[12]),
        .I4(\sr_reg[15]_0 [7]),
        .O(\badr[15]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'h0000E0EFEFEFEFEF)) 
    \badr[15]_INST_0_i_148 
       (.I0(\badrx[15]_INST_0_i_5_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(rst_n_fl_reg_9),
        .I3(\rgf_selc1_wb[0]_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_143_n_0 ),
        .I5(ir1[10]),
        .O(\badr[15]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBAAAAAAAA)) 
    \badr[15]_INST_0_i_149 
       (.I0(\badr[15]_INST_0_i_226_n_0 ),
        .I1(\bcmd[0]_INST_0_i_7_n_0 ),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_227_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_34_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_16_0 ),
        .O(\badr[15]_INST_0_i_149_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \badr[15]_INST_0_i_15 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\badr[15]_INST_0_i_26_n_0 ),
        .O(a1bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'hAAAB)) 
    \badr[15]_INST_0_i_150 
       (.I0(\badr[15]_INST_0_i_229_n_0 ),
        .I1(\badr[15]_INST_0_i_230_n_0 ),
        .I2(ir1[13]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_150_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F2FF00FF)) 
    \badr[15]_INST_0_i_151 
       (.I0(\badr[15]_INST_0_i_231_n_0 ),
        .I1(\badr[15]_INST_0_i_232_n_0 ),
        .I2(\badr[15]_INST_0_i_233_n_0 ),
        .I3(\badrx[15]_INST_0_i_5_n_0 ),
        .I4(\badr[15]_INST_0_i_234_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\badr[15]_INST_0_i_151_n_0 ));
  LUT5 #(
    .INIT(32'hFF1FFFFF)) 
    \badr[15]_INST_0_i_152 
       (.I0(ir1[14]),
        .I1(\sr_reg[15]_0 [7]),
        .I2(ir1[13]),
        .I3(ir1[15]),
        .I4(ir1[12]),
        .O(\badr[15]_INST_0_i_152_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_153 
       (.I0(ir1[6]),
        .I1(ir1[11]),
        .I2(ir1[15]),
        .I3(ir1[14]),
        .O(\badr[15]_INST_0_i_153_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_154 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .O(\badr[15]_INST_0_i_154_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_155 
       (.I0(ir1[10]),
        .I1(ir1[5]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[4]),
        .I5(ir1[2]),
        .O(\badr[15]_INST_0_i_155_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_156 
       (.I0(ir1[2]),
        .I1(ir1[6]),
        .O(\badr[15]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFF7DFFFDFF)) 
    \badr[15]_INST_0_i_157 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .I4(ir1[2]),
        .I5(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .O(\badr[15]_INST_0_i_157_n_0 ));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \badr[15]_INST_0_i_158 
       (.I0(\badr[15]_INST_0_i_28_0 ),
        .I1(\bdatw[9]_INST_0_i_69_n_0 ),
        .I2(\badr[15]_INST_0_i_236_n_0 ),
        .I3(\bdatw[15]_INST_0_i_186_n_0 ),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\badr[15]_INST_0_i_158_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_159 
       (.I0(ir1[11]),
        .I1(ir1[14]),
        .O(\badr[15]_INST_0_i_159_n_0 ));
  LUT5 #(
    .INIT(32'h00000200)) 
    \badr[15]_INST_0_i_160 
       (.I0(fch_irq_req),
        .I1(ir1[3]),
        .I2(ir1[2]),
        .I3(ir1[0]),
        .I4(ir1[1]),
        .O(\badr[15]_INST_0_i_160_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF1BFFFFFFFF)) 
    \badr[15]_INST_0_i_161 
       (.I0(ir1[8]),
        .I1(ir1[5]),
        .I2(ir1[2]),
        .I3(ir1[11]),
        .I4(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_6_n_0 ),
        .O(\badr[15]_INST_0_i_161_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0DCD050)) 
    \badr[15]_INST_0_i_162 
       (.I0(\badr[15]_INST_0_i_237_n_0 ),
        .I1(\badr[15]_INST_0_i_238_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[2]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_162_n_0 ));
  LUT5 #(
    .INIT(32'h01000000)) 
    \badr[15]_INST_0_i_163 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I4(ir1[9]),
        .O(\badr[15]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'h00040000FFFFFFFF)) 
    \badr[15]_INST_0_i_164 
       (.I0(\badr[15]_INST_0_i_239_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .I4(\badr[15]_INST_0_i_240_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_6_n_0 ),
        .O(\badr[15]_INST_0_i_164_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFEEEEFFFFFFFF)) 
    \badr[15]_INST_0_i_165 
       (.I0(\badr[15]_INST_0_i_241_n_0 ),
        .I1(\badr[15]_INST_0_i_242_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(\stat[2]_i_10__0_n_0 ),
        .I5(\badrx[15]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'hF8FFFAFFFAFFFAFF)) 
    \badr[15]_INST_0_i_166 
       (.I0(\bcmd[2]_INST_0_i_4_n_0 ),
        .I1(\stat[2]_i_10__0_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[0]),
        .I4(ir1[3]),
        .I5(\badr[15]_INST_0_i_243_n_0 ),
        .O(\badr[15]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFFFFFF)) 
    \badr[15]_INST_0_i_167 
       (.I0(\bcmd[0]_INST_0_i_7_n_0 ),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(\bdatw[15]_INST_0_i_186_n_0 ),
        .I3(ir1[13]),
        .I4(ir1[12]),
        .I5(\bdatw[9]_INST_0_i_69_n_0 ),
        .O(\badr[15]_INST_0_i_167_n_0 ));
  LUT5 #(
    .INIT(32'h8F8F0F8F)) 
    \badr[15]_INST_0_i_168 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[15]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .O(\badr[15]_INST_0_i_168_n_0 ));
  LUT6 #(
    .INIT(64'hFFBF0000FFFFFFFF)) 
    \badr[15]_INST_0_i_169 
       (.I0(ir1[11]),
        .I1(\badr[15]_INST_0_i_244_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I3(\bdatw[15]_INST_0_i_189_n_0 ),
        .I4(\badr[15]_INST_0_i_237_n_0 ),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEEAEAFEAEAAAA)) 
    \badr[15]_INST_0_i_170 
       (.I0(\badr[15]_INST_0_i_245_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[6]),
        .I3(ir1[3]),
        .I4(\badr[15]_INST_0_i_238_n_0 ),
        .I5(\badr[15]_INST_0_i_163_n_0 ),
        .O(\badr[15]_INST_0_i_170_n_0 ));
  LUT6 #(
    .INIT(64'h454545FF45454545)) 
    \badr[15]_INST_0_i_171 
       (.I0(\badr[15]_INST_0_i_246_n_0 ),
        .I1(\badr[15]_INST_0_i_247_n_0 ),
        .I2(ir1[9]),
        .I3(\badr[15]_INST_0_i_248_n_0 ),
        .I4(\badr[15]_INST_0_i_249_n_0 ),
        .I5(\badr[15]_INST_0_i_250_n_0 ),
        .O(\badr[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'h0400000004040000)) 
    \badr[15]_INST_0_i_173 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[9]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\badr[15]_INST_0_i_159_n_0 ),
        .I4(ir1[15]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_173_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF7FFFFFFFFFF)) 
    \badr[15]_INST_0_i_174 
       (.I0(\rgf_c1bus_wb[14]_i_53_0 ),
        .I1(\stat[2]_i_5__1_n_0 ),
        .I2(ir1[3]),
        .I3(ir1[1]),
        .I4(ir1[2]),
        .I5(\stat[1]_i_11__0_n_0 ),
        .O(\badr[15]_INST_0_i_174_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_175 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(\stat[2]_i_10__0_n_0 ),
        .I5(ir1[6]),
        .O(\badr[15]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'hEEE0FFFFEEEEFFFF)) 
    \badr[15]_INST_0_i_176 
       (.I0(ir1[6]),
        .I1(\bcmd[2]_INST_0_i_4_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .I3(\stat[2]_i_11_n_0 ),
        .I4(ir1[1]),
        .I5(fctl_n_96),
        .O(\badr[15]_INST_0_i_176_n_0 ));
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \badr[15]_INST_0_i_177 
       (.I0(\rgf_selc1_wb_reg[1]_0 ),
        .I1(\bdatw[9]_INST_0_i_69_n_0 ),
        .I2(\badr[15]_INST_0_i_236_n_0 ),
        .I3(\bdatw[15]_INST_0_i_186_n_0 ),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\badr[15]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'hDDDF0000FDFFFDFF)) 
    \badr[15]_INST_0_i_178 
       (.I0(ir1[9]),
        .I1(\bdatw[15]_INST_0_i_188_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[1]),
        .I4(\badr[15]_INST_0_i_237_n_0 ),
        .I5(ir1[4]),
        .O(\badr[15]_INST_0_i_178_n_0 ));
  LUT5 #(
    .INIT(32'h00A80020)) 
    \badr[15]_INST_0_i_179 
       (.I0(rst_n_fl_reg_9),
        .I1(ir1[8]),
        .I2(ir1[4]),
        .I3(ir1[9]),
        .I4(ir1[1]),
        .O(\badr[15]_INST_0_i_179_n_0 ));
  LUT6 #(
    .INIT(64'h0808000808000000)) 
    \badr[15]_INST_0_i_180 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I2(\badr[15]_INST_0_i_251_n_0 ),
        .I3(ir1[6]),
        .I4(ir1[1]),
        .I5(ir1[4]),
        .O(\badr[15]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'h0103030305030303)) 
    \badr[15]_INST_0_i_181 
       (.I0(ir1[1]),
        .I1(ir1[4]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'h0C008C8CCCC08C8C)) 
    \badr[15]_INST_0_i_182 
       (.I0(\rgf_selc1_rn_wb[1]_i_11_n_0 ),
        .I1(\badr[15]_INST_0_i_252_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[4]),
        .I4(ir1[9]),
        .I5(\badr[15]_INST_0_i_253_n_0 ),
        .O(\badr[15]_INST_0_i_182_n_0 ));
  LUT6 #(
    .INIT(64'h20000000000000A0)) 
    \badr[15]_INST_0_i_183 
       (.I0(\badr[15]_INST_0_i_254_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[1]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .I5(ir1[4]),
        .O(\badr[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFEFFFFFFFBFEF)) 
    \badr[15]_INST_0_i_184 
       (.I0(\stat[2]_i_11_n_0 ),
        .I1(ir1[4]),
        .I2(ir1[1]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'h0080008088880080)) 
    \badr[15]_INST_0_i_187 
       (.I0(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(\badr[15]_INST_0_i_255_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I5(ir0[6]),
        .O(\badr[15]_INST_0_i_187_n_0 ));
  LUT6 #(
    .INIT(64'h0A00AA0A0A000300)) 
    \badr[15]_INST_0_i_188 
       (.I0(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .I1(\badr[15]_INST_0_i_256_n_0 ),
        .I2(ir0[3]),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(ir0[2]),
        .O(\badr[15]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'h0004555500040004)) 
    \badr[15]_INST_0_i_189 
       (.I0(\badr[15]_INST_0_i_111_n_0 ),
        .I1(\badr[15]_INST_0_i_257_n_0 ),
        .I2(\badr[15]_INST_0_i_258_n_0 ),
        .I3(\badr[15]_INST_0_i_259_n_0 ),
        .I4(\badr[15]_INST_0_i_260_n_0 ),
        .I5(\badr[15]_INST_0_i_261_n_0 ),
        .O(\badr[15]_INST_0_i_189_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA2AAAAAAA)) 
    \badr[15]_INST_0_i_190 
       (.I0(\badr[15]_INST_0_i_262_n_0 ),
        .I1(\badr[15]_INST_0_i_263_n_0 ),
        .I2(\ccmd[0]_INST_0_i_11_n_0 ),
        .I3(\bdatw[11]_INST_0_i_17_n_0 ),
        .I4(\stat[1]_i_9__0_n_0 ),
        .I5(\badr[15]_INST_0_i_264_n_0 ),
        .O(\badr[15]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'h0010555500100010)) 
    \badr[15]_INST_0_i_191 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I3(\fadr[15]_INST_0_i_11_n_0 ),
        .I4(\badr[15]_INST_0_i_265_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .O(\badr[15]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'h00010101FFFFFFFF)) 
    \badr[15]_INST_0_i_192 
       (.I0(\badr[15]_INST_0_i_266_n_0 ),
        .I1(\badr[15]_INST_0_i_267_n_0 ),
        .I2(\badr[15]_INST_0_i_268_n_0 ),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_269_n_0 ),
        .I5(\badr[15]_INST_0_i_261_n_0 ),
        .O(\badr[15]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'h8880888088808888)) 
    \badr[15]_INST_0_i_193 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(\badr[15]_INST_0_i_270_n_0 ),
        .I3(\badr[15]_INST_0_i_271_n_0 ),
        .I4(ir0[10]),
        .I5(\badr[15]_INST_0_i_272_n_0 ),
        .O(\badr[15]_INST_0_i_193_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFBAFFBAFFBA)) 
    \badr[15]_INST_0_i_194 
       (.I0(\rgf_selc0_rn_wb[0]_i_16_n_0 ),
        .I1(\badr[15]_INST_0_i_273_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_15_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_201_n_0 ),
        .I5(\sr[13]_i_6_n_0 ),
        .O(\badr[15]_INST_0_i_194_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_195 
       (.I0(ir0[2]),
        .I1(ir0[6]),
        .O(\badr[15]_INST_0_i_195_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA00002000)) 
    \badr[15]_INST_0_i_196 
       (.I0(ir0[11]),
        .I1(\badr[15]_INST_0_i_274_n_0 ),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .I4(\bcmd[1]_INST_0_i_13_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .O(\badr[15]_INST_0_i_196_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7F7F700)) 
    \badr[15]_INST_0_i_197 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(crdy),
        .I2(\badr[15]_INST_0_i_275_n_0 ),
        .I3(\ccmd[4]_INST_0_i_20_n_0 ),
        .I4(\badr[15]_INST_0_i_276_n_0 ),
        .I5(\badr[15]_INST_0_i_277_n_0 ),
        .O(\badr[15]_INST_0_i_197_n_0 ));
  LUT6 #(
    .INIT(64'h0D082F7F0B0F4F0F)) 
    \badr[15]_INST_0_i_198 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[7]),
        .I4(ir0[2]),
        .I5(ir0[8]),
        .O(\badr[15]_INST_0_i_198_n_0 ));
  LUT6 #(
    .INIT(64'h11F111F1FFFF11F1)) 
    \badr[15]_INST_0_i_199 
       (.I0(\badr[15]_INST_0_i_278_n_0 ),
        .I1(\badr[15]_INST_0_i_274_n_0 ),
        .I2(\badr[15]_INST_0_i_279_n_0 ),
        .I3(\badr[15]_INST_0_i_280_n_0 ),
        .I4(ir0[5]),
        .I5(\badr[15]_INST_0_i_281_n_0 ),
        .O(\badr[15]_INST_0_i_199_n_0 ));
  LUT4 #(
    .INIT(16'h80FF)) 
    \badr[15]_INST_0_i_200 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[15]),
        .O(\badr[15]_INST_0_i_200_n_0 ));
  LUT5 #(
    .INIT(32'h00000200)) 
    \badr[15]_INST_0_i_201 
       (.I0(fch_irq_req),
        .I1(ir0[2]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ir0[3]),
        .O(\badr[15]_INST_0_i_201_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4440)) 
    \badr[15]_INST_0_i_202 
       (.I0(\fadr[15]_INST_0_i_11_n_0 ),
        .I1(\badr[15]_INST_0_i_282_n_0 ),
        .I2(crdy),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\badr[15]_INST_0_i_283_n_0 ),
        .O(\badr[15]_INST_0_i_202_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAABAFAFAAABA)) 
    \badr[15]_INST_0_i_203 
       (.I0(\badr[15]_INST_0_i_284_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[11]),
        .I3(\badr[15]_INST_0_i_281_n_0 ),
        .I4(\badr[15]_INST_0_i_285_n_0 ),
        .I5(\ccmd[3]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h000000000DCDFFFF)) 
    \badr[15]_INST_0_i_204 
       (.I0(\badr[15]_INST_0_i_286_n_0 ),
        .I1(\ccmd[4]_INST_0_i_12_n_0 ),
        .I2(\badr[15]_INST_0_i_287_n_0 ),
        .I3(crdy),
        .I4(ir0[8]),
        .I5(\badr[15]_INST_0_i_288_n_0 ),
        .O(\badr[15]_INST_0_i_204_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_205 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .O(\badr[15]_INST_0_i_205_n_0 ));
  LUT6 #(
    .INIT(64'h4444444444455545)) 
    \badr[15]_INST_0_i_206 
       (.I0(\ccmd[2]_INST_0_i_2_0 ),
        .I1(\badr[15]_INST_0_i_289_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[14]),
        .I4(\badr[15]_INST_0_i_290_n_0 ),
        .I5(\badr[15]_INST_0_i_291_n_0 ),
        .O(\badr[15]_INST_0_i_206_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \badr[15]_INST_0_i_207 
       (.I0(ir0[6]),
        .I1(\bcmd[0]_INST_0_i_20_n_0 ),
        .I2(ir0[2]),
        .I3(ir0[0]),
        .I4(\ccmd[0]_INST_0_i_11_n_0 ),
        .I5(\badr[15]_INST_0_i_292_n_0 ),
        .O(\badr[15]_INST_0_i_207_n_0 ));
  LUT6 #(
    .INIT(64'hF100FFFFF100F100)) 
    \badr[15]_INST_0_i_208 
       (.I0(\badr[15]_INST_0_i_293_n_0 ),
        .I1(\badr[15]_INST_0_i_294_n_0 ),
        .I2(\badr[15]_INST_0_i_114_0 ),
        .I3(\badr[15]_INST_0_i_296_n_0 ),
        .I4(\badr[15]_INST_0_i_297_n_0 ),
        .I5(\sr[13]_i_6_n_0 ),
        .O(\badr[15]_INST_0_i_208_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4555FFFF)) 
    \badr[15]_INST_0_i_209 
       (.I0(\badr[15]_INST_0_i_298_n_0 ),
        .I1(\badr[15]_INST_0_i_204_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[12]),
        .I4(ir0[13]),
        .I5(\badr[15]_INST_0_i_299_n_0 ),
        .O(\badr[15]_INST_0_i_209_n_0 ));
  LUT5 #(
    .INIT(32'h08000000)) 
    \badr[15]_INST_0_i_210 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(\stat_reg[2]_18 ),
        .O(a0bus_sel_0[1]));
  LUT5 #(
    .INIT(32'h00000800)) 
    \badr[15]_INST_0_i_211 
       (.I0(\stat_reg[2]_20 ),
        .I1(ctl_sela0),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(\stat_reg[2]_18 ),
        .O(a0bus_sel_0[2]));
  LUT6 #(
    .INIT(64'hFF00FF01FFFFFF01)) 
    \badr[15]_INST_0_i_224 
       (.I0(\badr[15]_INST_0_i_300_n_0 ),
        .I1(\badr[15]_INST_0_i_175_n_0 ),
        .I2(ir1[14]),
        .I3(\badr[15]_INST_0_i_301_n_0 ),
        .I4(ir1[12]),
        .I5(\badr[15]_INST_0_i_25_0 ),
        .O(\badr[15]_INST_0_i_224_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF02)) 
    \badr[15]_INST_0_i_225 
       (.I0(\badr[15]_INST_0_i_169_n_0 ),
        .I1(\badr[15]_INST_0_i_302_n_0 ),
        .I2(\badr[15]_INST_0_i_245_n_0 ),
        .I3(ir1[11]),
        .I4(\badr[15]_INST_0_i_303_n_0 ),
        .I5(\badr[15]_INST_0_i_304_n_0 ),
        .O(\badr[15]_INST_0_i_225_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_226 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .O(\badr[15]_INST_0_i_226_n_0 ));
  LUT4 #(
    .INIT(16'hB0FB)) 
    \badr[15]_INST_0_i_227 
       (.I0(ir1[1]),
        .I1(ir1[2]),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .O(\badr[15]_INST_0_i_227_n_0 ));
  LUT5 #(
    .INIT(32'h000022BA)) 
    \badr[15]_INST_0_i_229 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .I2(\sr_reg[15]_0 [6]),
        .I3(ir1[12]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_229_n_0 ));
  LUT6 #(
    .INIT(64'h4404000411045504)) 
    \badr[15]_INST_0_i_230 
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(\sr_reg[15]_0 [4]),
        .I3(ir1[14]),
        .I4(\sr_reg[15]_0 [7]),
        .I5(\sr_reg[15]_0 [5]),
        .O(\badr[15]_INST_0_i_230_n_0 ));
  LUT5 #(
    .INIT(32'hC4CFCFC4)) 
    \badr[15]_INST_0_i_231 
       (.I0(ir1[7]),
        .I1(ir1[10]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .O(\badr[15]_INST_0_i_231_n_0 ));
  LUT6 #(
    .INIT(64'h000003000000AB03)) 
    \badr[15]_INST_0_i_232 
       (.I0(ir1[3]),
        .I1(ir1[6]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[7]),
        .I4(ir1[4]),
        .I5(ir1[5]),
        .O(\badr[15]_INST_0_i_232_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_233 
       (.I0(ir1[6]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_233_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFEFFFEFFFFFFF)) 
    \badr[15]_INST_0_i_234 
       (.I0(ir1[3]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_234_n_0 ));
  LUT5 #(
    .INIT(32'h00083F3F)) 
    \badr[15]_INST_0_i_235 
       (.I0(ir1[7]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\badr[15]_INST_0_i_235_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_236 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .O(\badr[15]_INST_0_i_236_n_0 ));
  LUT5 #(
    .INIT(32'hFF2AFFFF)) 
    \badr[15]_INST_0_i_237 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .O(\badr[15]_INST_0_i_237_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_238 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .O(\badr[15]_INST_0_i_238_n_0 ));
  LUT6 #(
    .INIT(64'h000B0008000F0000)) 
    \badr[15]_INST_0_i_239 
       (.I0(ir1[2]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[5]),
        .I5(ir1[7]),
        .O(\badr[15]_INST_0_i_239_n_0 ));
  LUT6 #(
    .INIT(64'hAA20AA20AA20AAAA)) 
    \badr[15]_INST_0_i_24 
       (.I0(\read_cyc_reg[1] ),
        .I1(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .I2(\badr[15]_INST_0_i_70_n_0 ),
        .I3(\badr[15]_INST_0_i_71_n_0 ),
        .I4(\badr[15]_INST_0_i_72_n_0 ),
        .I5(\badr[15]_INST_0_i_73_n_0 ),
        .O(ctl_sela1));
  LUT5 #(
    .INIT(32'h757F7777)) 
    \badr[15]_INST_0_i_240 
       (.I0(ir1[9]),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[2]),
        .I4(ir1[8]),
        .O(\badr[15]_INST_0_i_240_n_0 ));
  LUT6 #(
    .INIT(64'h00005D5D005D5D5D)) 
    \badr[15]_INST_0_i_241 
       (.I0(ir1[2]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(ir1[5]),
        .I4(ir1[7]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_241_n_0 ));
  LUT5 #(
    .INIT(32'h22002F00)) 
    \badr[15]_INST_0_i_242 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .O(\badr[15]_INST_0_i_242_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \badr[15]_INST_0_i_243 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .O(\badr[15]_INST_0_i_243_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_244 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .O(\badr[15]_INST_0_i_244_n_0 ));
  LUT6 #(
    .INIT(64'h1010100000001000)) 
    \badr[15]_INST_0_i_245 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I3(ir1[3]),
        .I4(ir1[8]),
        .I5(ir1[0]),
        .O(\badr[15]_INST_0_i_245_n_0 ));
  LUT6 #(
    .INIT(64'hAABAFFFFBBBBFFFF)) 
    \badr[15]_INST_0_i_246 
       (.I0(\badr[15]_INST_0_i_305_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[6]),
        .I3(\stat[2]_i_10__0_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_246_n_0 ));
  LUT6 #(
    .INIT(64'h00000000CCCC8088)) 
    \badr[15]_INST_0_i_247 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[0]),
        .I5(\badr[15]_INST_0_i_306_n_0 ),
        .O(\badr[15]_INST_0_i_247_n_0 ));
  LUT6 #(
    .INIT(64'h0100000001030303)) 
    \badr[15]_INST_0_i_248 
       (.I0(ir1[0]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[3]),
        .O(\badr[15]_INST_0_i_248_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0A22FFFFFFFF)) 
    \badr[15]_INST_0_i_249 
       (.I0(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .I3(ir1[7]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\badr[15]_INST_0_i_249_n_0 ));
  LUT6 #(
    .INIT(64'h5555555500545555)) 
    \badr[15]_INST_0_i_25 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\badr[15]_INST_0_i_74_n_0 ),
        .I2(\badr[15]_INST_0_i_75_n_0 ),
        .I3(\badr[15]_INST_0_i_76_n_0 ),
        .I4(\badr[15]_INST_0_i_77_n_0 ),
        .I5(\badr[15]_INST_0_i_78_n_0 ),
        .O(\badr[15]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hEF4FFF0F)) 
    \badr[15]_INST_0_i_250 
       (.I0(ir1[6]),
        .I1(ir1[0]),
        .I2(ir1[9]),
        .I3(ir1[3]),
        .I4(ir1[8]),
        .O(\badr[15]_INST_0_i_250_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[15]_INST_0_i_251 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .O(\badr[15]_INST_0_i_251_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_252 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\badr[15]_INST_0_i_252_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \badr[15]_INST_0_i_253 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .I2(ir1[1]),
        .O(\badr[15]_INST_0_i_253_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_254 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .O(\badr[15]_INST_0_i_254_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_255 
       (.I0(\bcmd[1]_INST_0_i_13_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\badr[15]_INST_0_i_255_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    \badr[15]_INST_0_i_256 
       (.I0(\ccmd[4]_INST_0_i_15_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I4(ir0[15]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\badr[15]_INST_0_i_256_n_0 ));
  LUT6 #(
    .INIT(64'h4070FFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_257 
       (.I0(\badr[15]_INST_0_i_307_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(\badr[15]_INST_0_i_308_n_0 ),
        .I4(ir0[9]),
        .I5(ir0[10]),
        .O(\badr[15]_INST_0_i_257_n_0 ));
  LUT6 #(
    .INIT(64'h55555555555577F7)) 
    \badr[15]_INST_0_i_258 
       (.I0(\bcmd[1]_INST_0_i_6_n_0 ),
        .I1(ir0[4]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_20_n_0 ),
        .I5(\badr[15]_INST_0_i_309_n_0 ),
        .O(\badr[15]_INST_0_i_258_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055155511)) 
    \badr[15]_INST_0_i_259 
       (.I0(ir0[10]),
        .I1(ir0[4]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(\rgf_selc0_rn_wb[1]_i_27_n_0 ),
        .I5(\badr[15]_INST_0_i_310_n_0 ),
        .O(\badr[15]_INST_0_i_259_n_0 ));
  LUT6 #(
    .INIT(64'h5454545544444444)) 
    \badr[15]_INST_0_i_26 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\badr[15]_INST_0_i_79_n_0 ),
        .I2(\badr[15]_INST_0_i_80_n_0 ),
        .I3(\badr[15]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_82_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_53_0 ),
        .O(\badr[15]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000F700F7F7F7F7)) 
    \badr[15]_INST_0_i_260 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(crdy),
        .I2(\badr[15]_INST_0_i_311_n_0 ),
        .I3(\badr[15]_INST_0_i_312_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I5(ir0[10]),
        .O(\badr[15]_INST_0_i_260_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_261 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .O(\badr[15]_INST_0_i_261_n_0 ));
  LUT6 #(
    .INIT(64'hDFFF5F5F5F5F5F5F)) 
    \badr[15]_INST_0_i_262 
       (.I0(ir0[15]),
        .I1(ir0[14]),
        .I2(ir0[9]),
        .I3(ir0[11]),
        .I4(ir0[12]),
        .I5(ir0[13]),
        .O(\badr[15]_INST_0_i_262_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_263 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .O(\badr[15]_INST_0_i_263_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_264 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .O(\badr[15]_INST_0_i_264_n_0 ));
  LUT6 #(
    .INIT(64'hB0BBBBBBFFFFFFFF)) 
    \badr[15]_INST_0_i_265 
       (.I0(ir0[6]),
        .I1(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .I4(ir0[3]),
        .I5(ir0[0]),
        .O(\badr[15]_INST_0_i_265_n_0 ));
  LUT6 #(
    .INIT(64'h4055000000000000)) 
    \badr[15]_INST_0_i_266 
       (.I0(\ccmd[4]_INST_0_i_20_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(crdy),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_266_n_0 ));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    \badr[15]_INST_0_i_267 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .I3(ir0[0]),
        .I4(ir0[6]),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_267_n_0 ));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \badr[15]_INST_0_i_268 
       (.I0(\ccmd[4]_INST_0_i_20_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(crdy),
        .I4(ir0[6]),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_268_n_0 ));
  LUT5 #(
    .INIT(32'h0AAC0CAC)) 
    \badr[15]_INST_0_i_269 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[6]),
        .O(\badr[15]_INST_0_i_269_n_0 ));
  LUT6 #(
    .INIT(64'h5454545544444444)) 
    \badr[15]_INST_0_i_27 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\badr[15]_INST_0_i_83_n_0 ),
        .I2(\badr[15]_INST_0_i_84_n_0 ),
        .I3(\bcmd[2]_INST_0_i_7_n_0 ),
        .I4(\badr[15]_INST_0_i_85_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_53_0 ),
        .O(\stat_reg[2]_15 ));
  LUT6 #(
    .INIT(64'h0055000004400504)) 
    \badr[15]_INST_0_i_270 
       (.I0(\badr[15]_INST_0_i_274_n_0 ),
        .I1(ir0[0]),
        .I2(ir0[4]),
        .I3(ir0[3]),
        .I4(ir0[6]),
        .I5(ir0[5]),
        .O(\badr[15]_INST_0_i_270_n_0 ));
  LUT6 #(
    .INIT(64'h3000FFFFB000B000)) 
    \badr[15]_INST_0_i_271 
       (.I0(\badr[15]_INST_0_i_313_n_0 ),
        .I1(\bcmd[1]_INST_0_i_13_n_0 ),
        .I2(ir0[0]),
        .I3(\badr[15]_INST_0_i_279_n_0 ),
        .I4(\badr[15]_INST_0_i_281_n_0 ),
        .I5(ir0[3]),
        .O(\badr[15]_INST_0_i_271_n_0 ));
  LUT6 #(
    .INIT(64'h22773333303F13B3)) 
    \badr[15]_INST_0_i_272 
       (.I0(ir0[6]),
        .I1(ir0[3]),
        .I2(ir0[7]),
        .I3(ir0[0]),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\badr[15]_INST_0_i_272_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \badr[15]_INST_0_i_273 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .O(\badr[15]_INST_0_i_273_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \badr[15]_INST_0_i_274 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .O(\badr[15]_INST_0_i_274_n_0 ));
  LUT5 #(
    .INIT(32'hCF08CF7F)) 
    \badr[15]_INST_0_i_275 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[2]),
        .I3(ir0[8]),
        .I4(ir0[5]),
        .O(\badr[15]_INST_0_i_275_n_0 ));
  LUT5 #(
    .INIT(32'h707FFFFF)) 
    \badr[15]_INST_0_i_276 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[5]),
        .O(\badr[15]_INST_0_i_276_n_0 ));
  LUT6 #(
    .INIT(64'h8080008080000000)) 
    \badr[15]_INST_0_i_277 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(ir0[2]),
        .O(\badr[15]_INST_0_i_277_n_0 ));
  LUT5 #(
    .INIT(32'hF1B5FFAB)) 
    \badr[15]_INST_0_i_278 
       (.I0(ir0[5]),
        .I1(ir0[2]),
        .I2(ir0[3]),
        .I3(ir0[4]),
        .I4(ir0[6]),
        .O(\badr[15]_INST_0_i_278_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \badr[15]_INST_0_i_279 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .O(\badr[15]_INST_0_i_279_n_0 ));
  LUT6 #(
    .INIT(64'h5554555554545454)) 
    \badr[15]_INST_0_i_28 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\badr[15]_INST_0_i_86_n_0 ),
        .I2(\badr[15]_INST_0_i_87_n_0 ),
        .I3(\badr[15]_INST_0_i_88_n_0 ),
        .I4(\badr[15]_INST_0_i_89_n_0 ),
        .I5(\badr[15]_INST_0_i_90_n_0 ),
        .O(\stat_reg[2]_16 ));
  LUT5 #(
    .INIT(32'hFEFF7EFF)) 
    \badr[15]_INST_0_i_280 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[2]),
        .I4(ir0[3]),
        .O(\badr[15]_INST_0_i_280_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFFFFFF2FFF2FF)) 
    \badr[15]_INST_0_i_281 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(crdy),
        .I5(ir0[8]),
        .O(\badr[15]_INST_0_i_281_n_0 ));
  LUT4 #(
    .INIT(16'h2A02)) 
    \badr[15]_INST_0_i_282 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .O(\badr[15]_INST_0_i_282_n_0 ));
  LUT6 #(
    .INIT(64'h1400110055001500)) 
    \badr[15]_INST_0_i_283 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[15]),
        .I4(ir0[11]),
        .I5(ir0[14]),
        .O(\badr[15]_INST_0_i_283_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \badr[15]_INST_0_i_284 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[11]),
        .I3(ir0[10]),
        .I4(\badr[15]_INST_0_i_314_n_0 ),
        .O(\badr[15]_INST_0_i_284_n_0 ));
  LUT6 #(
    .INIT(64'h1101010100010101)) 
    \badr[15]_INST_0_i_285 
       (.I0(\badr[15]_INST_0_i_315_n_0 ),
        .I1(ir0[10]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_285_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_286 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .O(\badr[15]_INST_0_i_286_n_0 ));
  LUT4 #(
    .INIT(16'h3222)) 
    \badr[15]_INST_0_i_287 
       (.I0(ir0[9]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .O(\badr[15]_INST_0_i_287_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_288 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[8]),
        .I2(crdy),
        .I3(ir0[9]),
        .O(\badr[15]_INST_0_i_288_n_0 ));
  LUT4 #(
    .INIT(16'hFF01)) 
    \badr[15]_INST_0_i_289 
       (.I0(\badr[15]_INST_0_i_316_n_0 ),
        .I1(ir0[13]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\badr[15]_INST_0_i_317_n_0 ),
        .O(\badr[15]_INST_0_i_289_n_0 ));
  LUT6 #(
    .INIT(64'h0008AAAAAAAAAAAA)) 
    \badr[15]_INST_0_i_290 
       (.I0(\badr[15]_INST_0_i_318_n_0 ),
        .I1(\badr[15]_INST_0_i_319_n_0 ),
        .I2(\badr[15]_INST_0_i_320_n_0 ),
        .I3(\badr[15]_INST_0_i_321_n_0 ),
        .I4(ir0[9]),
        .I5(ir0[8]),
        .O(\badr[15]_INST_0_i_290_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1FFF)) 
    \badr[15]_INST_0_i_291 
       (.I0(\sr_reg[15]_0 [7]),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(ir0[15]),
        .O(\badr[15]_INST_0_i_291_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    \badr[15]_INST_0_i_292 
       (.I0(ir0[13]),
        .I1(\badr[15]_INST_0_i_322_n_0 ),
        .I2(\ccmd[3]_INST_0_i_21_n_0 ),
        .I3(ir0[3]),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(ir0[1]),
        .O(\badr[15]_INST_0_i_292_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \badr[15]_INST_0_i_293 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(ir0[8]),
        .I4(\badr[15]_INST_0_i_323_n_0 ),
        .I5(ir0[9]),
        .O(\badr[15]_INST_0_i_293_n_0 ));
  LUT6 #(
    .INIT(64'hFF0C3F1DFFCCFF3F)) 
    \badr[15]_INST_0_i_294 
       (.I0(fch_irq_req),
        .I1(ir0[2]),
        .I2(crdy),
        .I3(ir0[3]),
        .I4(ir0[1]),
        .I5(ir0[0]),
        .O(\badr[15]_INST_0_i_294_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_296 
       (.I0(ir0[13]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\badr[15]_INST_0_i_296_n_0 ));
  LUT5 #(
    .INIT(32'hC4FDFFFF)) 
    \badr[15]_INST_0_i_297 
       (.I0(ir0[2]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\badr[15]_INST_0_i_297_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAABAAAAAA)) 
    \badr[15]_INST_0_i_298 
       (.I0(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I1(ir0[10]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_12_n_0 ),
        .I5(\stat[2]_i_12_n_0 ),
        .O(\badr[15]_INST_0_i_298_n_0 ));
  LUT6 #(
    .INIT(64'hCFCFCFCCCF02CF02)) 
    \badr[15]_INST_0_i_299 
       (.I0(\sr_reg[15]_0 [6]),
        .I1(ir0[15]),
        .I2(ir0[14]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\sr_reg[15]_0 [7]),
        .I5(ir0[12]),
        .O(\badr[15]_INST_0_i_299_n_0 ));
  LUT5 #(
    .INIT(32'hCE4DCE5D)) 
    \badr[15]_INST_0_i_300 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(fch_irq_req),
        .O(\badr[15]_INST_0_i_300_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF04)) 
    \badr[15]_INST_0_i_301 
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .I2(\sr_reg[15]_0 [5]),
        .I3(ir1[13]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[15]),
        .O(\badr[15]_INST_0_i_301_n_0 ));
  LUT6 #(
    .INIT(64'h08000000FFFFFFFF)) 
    \badr[15]_INST_0_i_302 
       (.I0(ir1[6]),
        .I1(ir1[0]),
        .I2(\badr[15]_INST_0_i_251_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I4(ir1[9]),
        .I5(\badr[15]_INST_0_i_324_n_0 ),
        .O(\badr[15]_INST_0_i_302_n_0 ));
  LUT6 #(
    .INIT(64'h00000000002A0000)) 
    \badr[15]_INST_0_i_303 
       (.I0(\badr[15]_INST_0_i_250_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_17_n_0 ),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .I5(\badr[15]_INST_0_i_248_n_0 ),
        .O(\badr[15]_INST_0_i_303_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000005D)) 
    \badr[15]_INST_0_i_304 
       (.I0(ir1[9]),
        .I1(\badr[15]_INST_0_i_325_n_0 ),
        .I2(\badr[15]_INST_0_i_306_n_0 ),
        .I3(\badr[15]_INST_0_i_326_n_0 ),
        .I4(\badr[15]_INST_0_i_327_n_0 ),
        .I5(\badr[15]_INST_0_i_305_n_0 ),
        .O(\badr[15]_INST_0_i_304_n_0 ));
  LUT5 #(
    .INIT(32'h0000444F)) 
    \badr[15]_INST_0_i_305 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .I4(ir1[6]),
        .O(\badr[15]_INST_0_i_305_n_0 ));
  LUT5 #(
    .INIT(32'hAFBFBF30)) 
    \badr[15]_INST_0_i_306 
       (.I0(ir1[3]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[4]),
        .O(\badr[15]_INST_0_i_306_n_0 ));
  LUT5 #(
    .INIT(32'h0FD7FFFD)) 
    \badr[15]_INST_0_i_307 
       (.I0(ir0[1]),
        .I1(ir0[4]),
        .I2(ir0[3]),
        .I3(ir0[5]),
        .I4(ir0[6]),
        .O(\badr[15]_INST_0_i_307_n_0 ));
  LUT5 #(
    .INIT(32'hFEFF7EFF)) 
    \badr[15]_INST_0_i_308 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[1]),
        .I4(ir0[3]),
        .O(\badr[15]_INST_0_i_308_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[15]_INST_0_i_309 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .O(\badr[15]_INST_0_i_309_n_0 ));
  LUT6 #(
    .INIT(64'hEE00FA8022000A80)) 
    \badr[15]_INST_0_i_310 
       (.I0(ir0[1]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(ir0[4]),
        .O(\badr[15]_INST_0_i_310_n_0 ));
  LUT5 #(
    .INIT(32'hC0F8C7FF)) 
    \badr[15]_INST_0_i_311 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(ir0[1]),
        .I4(ir0[4]),
        .O(\badr[15]_INST_0_i_311_n_0 ));
  LUT6 #(
    .INIT(64'h1F1FF0FFBFBFFFFF)) 
    \badr[15]_INST_0_i_312 
       (.I0(ir0[6]),
        .I1(ir0[1]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[9]),
        .I5(ir0[4]),
        .O(\badr[15]_INST_0_i_312_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_313 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .O(\badr[15]_INST_0_i_313_n_0 ));
  LUT6 #(
    .INIT(64'hFFEBFFDFFBFEFFFA)) 
    \badr[15]_INST_0_i_314 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\badr[15]_INST_0_i_314_n_0 ));
  LUT6 #(
    .INIT(64'h8000808880008080)) 
    \badr[15]_INST_0_i_315 
       (.I0(ir0[8]),
        .I1(ir0[6]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[9]),
        .I4(ir0[7]),
        .I5(ir0[11]),
        .O(\badr[15]_INST_0_i_315_n_0 ));
  LUT6 #(
    .INIT(64'h4404000411045504)) 
    \badr[15]_INST_0_i_316 
       (.I0(ir0[15]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_0 [4]),
        .I3(ir0[14]),
        .I4(\sr_reg[15]_0 [7]),
        .I5(\sr_reg[15]_0 [5]),
        .O(\badr[15]_INST_0_i_316_n_0 ));
  LUT5 #(
    .INIT(32'h00003F02)) 
    \badr[15]_INST_0_i_317 
       (.I0(\sr_reg[15]_0 [6]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\badr[15]_INST_0_i_317_n_0 ));
  LUT6 #(
    .INIT(64'hFFBBFFFFFF0A0000)) 
    \badr[15]_INST_0_i_318 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(crdy),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\badr[15]_INST_0_i_318_n_0 ));
  LUT6 #(
    .INIT(64'hFFFCFDDCFFFFFFFC)) 
    \badr[15]_INST_0_i_319 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(ir0[7]),
        .O(\badr[15]_INST_0_i_319_n_0 ));
  LUT6 #(
    .INIT(64'h1000100010000000)) 
    \badr[15]_INST_0_i_320 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[3]),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .I4(ir0[7]),
        .I5(ir0[5]),
        .O(\badr[15]_INST_0_i_320_n_0 ));
  LUT5 #(
    .INIT(32'h0C50005D)) 
    \badr[15]_INST_0_i_321 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .O(\badr[15]_INST_0_i_321_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_322 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .O(\badr[15]_INST_0_i_322_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_323 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .O(\badr[15]_INST_0_i_323_n_0 ));
  LUT6 #(
    .INIT(64'h1DFFFFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_324 
       (.I0(ir1[0]),
        .I1(ir1[6]),
        .I2(ir1[3]),
        .I3(ir1[8]),
        .I4(ir1[10]),
        .I5(ir1[9]),
        .O(\badr[15]_INST_0_i_324_n_0 ));
  LUT5 #(
    .INIT(32'hFB00AA00)) 
    \badr[15]_INST_0_i_325 
       (.I0(ir1[0]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .O(\badr[15]_INST_0_i_325_n_0 ));
  LUT4 #(
    .INIT(16'h777F)) 
    \badr[15]_INST_0_i_326 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[3]),
        .I3(ir1[9]),
        .O(\badr[15]_INST_0_i_326_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \badr[15]_INST_0_i_327 
       (.I0(ir1[3]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(ir1[5]),
        .O(\badr[15]_INST_0_i_327_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \badr[15]_INST_0_i_35 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sel_cr[4]));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[15]_INST_0_i_37 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .O(a1bus_sel_cr[1]));
  LUT5 #(
    .INIT(32'h00040000)) 
    \badr[15]_INST_0_i_38 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\badr[15]_INST_0_i_26_n_0 ),
        .I4(\stat_reg[2]_15 ),
        .O(a1bus_sel_cr[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_39 
       (.I0(\stat_reg[2]_18 ),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF575555)) 
    \badr[15]_INST_0_i_40 
       (.I0(\badr[15]_INST_0_i_109_n_0 ),
        .I1(\badr[15]_INST_0_i_110_n_0 ),
        .I2(\badr[15]_INST_0_i_111_n_0 ),
        .I3(\badr[15]_INST_0_i_112_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(ctl_sela0_rn[1]));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_41 
       (.I0(ctl_sela0),
        .I1(\stat_reg[2]_20 ),
        .O(\badr[15]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_42 
       (.I0(\stat_reg[2]_18 ),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_51 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_18 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(a0bus_sel_cr[0]));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_56 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_18 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(a0bus_sel_cr[3]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_57 
       (.I0(ctl_sela0_rn[1]),
        .I1(ctl_sela0_rn[0]),
        .I2(\stat_reg[2]_18 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(a0bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_58 
       (.I0(\stat_reg[2]_18 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(a0bus_sel_cr[1]));
  LUT6 #(
    .INIT(64'h0100010100000000)) 
    \badr[15]_INST_0_i_59 
       (.I0(\badr[15]_INST_0_i_139_n_0 ),
        .I1(\stat_reg[2]_16 ),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(\badr[15]_INST_0_i_83_n_0 ),
        .I4(\badr[15]_INST_0_i_140_n_0 ),
        .I5(\badr[15]_INST_0_i_26_n_0 ),
        .O(a1bus_sel_0[1]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[15]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [15]),
        .O(a1bus_sr[15]));
  LUT6 #(
    .INIT(64'h4544000000000000)) 
    \badr[15]_INST_0_i_60 
       (.I0(\badr[15]_INST_0_i_139_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(\badr[15]_INST_0_i_83_n_0 ),
        .I3(\badr[15]_INST_0_i_140_n_0 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\badr[15]_INST_0_i_26_n_0 ),
        .O(a1bus_sel_0[2]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_61 
       (.I0(\badr[15]_INST_0_i_26_n_0 ),
        .I1(\badr[15]_INST_0_i_139_n_0 ),
        .O(\stat_reg[2]_14 ));
  LUT6 #(
    .INIT(64'h0200020200000000)) 
    \badr[15]_INST_0_i_62 
       (.I0(\badr[15]_INST_0_i_26_n_0 ),
        .I1(\badr[15]_INST_0_i_139_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(\badr[15]_INST_0_i_83_n_0 ),
        .I4(\badr[15]_INST_0_i_140_n_0 ),
        .I5(\stat_reg[2]_16 ),
        .O(a1bus_sel_0[3]));
  LUT4 #(
    .INIT(16'h088A)) 
    \badr[15]_INST_0_i_70 
       (.I0(ir1[2]),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .I3(ir1[3]),
        .O(\badr[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h030B090F00000000)) 
    \badr[15]_INST_0_i_71 
       (.I0(ir1[11]),
        .I1(ir1[12]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[14]),
        .I4(ir1[13]),
        .I5(ir1[15]),
        .O(\badr[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0F0F0D0D0F000)) 
    \badr[15]_INST_0_i_72 
       (.I0(ir1[8]),
        .I1(\badr[15]_INST_0_i_142_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[9]),
        .I5(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .O(\badr[15]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h01FF00FF01FFFFFF)) 
    \badr[15]_INST_0_i_73 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb[0]_i_18_n_0 ),
        .I2(\badr[15]_INST_0_i_143_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I4(ir1[10]),
        .I5(\badr[15]_INST_0_i_144_n_0 ),
        .O(\badr[15]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFCFFFCFCF)) 
    \badr[15]_INST_0_i_74 
       (.I0(\badr[15]_INST_0_i_25_0 ),
        .I1(ir1[15]),
        .I2(\badr[15]_INST_0_i_146_n_0 ),
        .I3(\sr_reg[15]_0 [5]),
        .I4(ir1[14]),
        .I5(ir1[12]),
        .O(\badr[15]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0A00AA0A0000A8A0)) 
    \badr[15]_INST_0_i_75 
       (.I0(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I1(fch_irq_req),
        .I2(ir1[1]),
        .I3(ir1[0]),
        .I4(ir1[3]),
        .I5(ir1[2]),
        .O(\badr[15]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8A808A8A)) 
    \badr[15]_INST_0_i_76 
       (.I0(ir1[13]),
        .I1(\badr[15]_INST_0_i_147_n_0 ),
        .I2(\bcmd[2]_INST_0_i_7_n_0 ),
        .I3(\badr[15]_INST_0_i_148_n_0 ),
        .I4(ir1[12]),
        .I5(\badr[15]_INST_0_i_149_n_0 ),
        .O(\badr[15]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBAAABA)) 
    \badr[15]_INST_0_i_77 
       (.I0(\rgf_selc1_wb_reg[0] ),
        .I1(\badr[15]_INST_0_i_150_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[14]),
        .I4(\badr[15]_INST_0_i_151_n_0 ),
        .I5(\badr[15]_INST_0_i_152_n_0 ),
        .O(\badr[15]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \badr[15]_INST_0_i_78 
       (.I0(\badr[15]_INST_0_i_153_n_0 ),
        .I1(\badr[15]_INST_0_i_154_n_0 ),
        .I2(ir1[9]),
        .I3(\fch_irq_lev[1]_i_5_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\badr[15]_INST_0_i_155_n_0 ),
        .O(\badr[15]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2F220000)) 
    \badr[15]_INST_0_i_79 
       (.I0(\badr[15]_INST_0_i_156_n_0 ),
        .I1(\bcmd[2]_INST_0_i_4_n_0 ),
        .I2(\badr[15]_INST_0_i_157_n_0 ),
        .I3(ir1[11]),
        .I4(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I5(\badr[15]_INST_0_i_158_n_0 ),
        .O(\badr[15]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hC400FFFFC400C400)) 
    \badr[15]_INST_0_i_80 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(ir1[15]),
        .I2(\badr[15]_INST_0_i_159_n_0 ),
        .I3(ir1[10]),
        .I4(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .I5(\badr[15]_INST_0_i_160_n_0 ),
        .O(\badr[15]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h0002220222222222)) 
    \badr[15]_INST_0_i_81 
       (.I0(\badr[15]_INST_0_i_161_n_0 ),
        .I1(\badr[15]_INST_0_i_162_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[2]),
        .I5(\badr[15]_INST_0_i_163_n_0 ),
        .O(\badr[15]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \badr[15]_INST_0_i_82 
       (.I0(\badr[15]_INST_0_i_164_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I5(\badr[15]_INST_0_i_165_n_0 ),
        .O(\badr[15]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h002000200020EEEE)) 
    \badr[15]_INST_0_i_83 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I3(\badr[15]_INST_0_i_166_n_0 ),
        .I4(ir1[15]),
        .I5(\badr[15]_INST_0_i_167_n_0 ),
        .O(\badr[15]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'hD555FFFFD555D555)) 
    \badr[15]_INST_0_i_84 
       (.I0(\sr_reg[4] ),
        .I1(\bdatw[9]_INST_0_i_69_n_0 ),
        .I2(fch_irq_req),
        .I3(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I4(\badr[15]_INST_0_i_168_n_0 ),
        .I5(ir1[8]),
        .O(\badr[15]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h0000AA08AAAAAAAA)) 
    \badr[15]_INST_0_i_85 
       (.I0(\stat[1]_i_6__0_n_0 ),
        .I1(\badr[15]_INST_0_i_169_n_0 ),
        .I2(\badr[15]_INST_0_i_170_n_0 ),
        .I3(ir1[11]),
        .I4(\badr[15]_INST_0_i_171_n_0 ),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h08A8000800000000)) 
    \badr[15]_INST_0_i_86 
       (.I0(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[1]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .I5(\badr[15]_INST_0_i_28_0 ),
        .O(\badr[15]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFABABFFAB)) 
    \badr[15]_INST_0_i_87 
       (.I0(\badr[15]_INST_0_i_173_n_0 ),
        .I1(\badr[15]_INST_0_i_174_n_0 ),
        .I2(\badr[15]_INST_0_i_175_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I4(\badr[15]_INST_0_i_176_n_0 ),
        .I5(\badr[15]_INST_0_i_177_n_0 ),
        .O(\badr[15]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h00FDFFFF00FD00FD)) 
    \badr[15]_INST_0_i_88 
       (.I0(\badr[15]_INST_0_i_178_n_0 ),
        .I1(\badr[15]_INST_0_i_179_n_0 ),
        .I2(\badr[15]_INST_0_i_180_n_0 ),
        .I3(ir1[11]),
        .I4(\badr[15]_INST_0_i_181_n_0 ),
        .I5(\badr[15]_INST_0_i_182_n_0 ),
        .O(\badr[15]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h4F0F4F0F4F0F4FFF)) 
    \badr[15]_INST_0_i_89 
       (.I0(\badr[15]_INST_0_i_183_n_0 ),
        .I1(\badr[15]_INST_0_i_184_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I3(ir1[9]),
        .I4(ir1[4]),
        .I5(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .O(\badr[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [15]),
        .I5(\iv_reg[15]_0 [15]),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \badr[15]_INST_0_i_90 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\rgf_selc1_wb_reg[1] [1]),
        .O(\badr[15]_INST_0_i_90_n_0 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[1]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[1]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[1]),
        .O(badr[0]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[1]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [1]),
        .O(a1bus_sr[1]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [1]),
        .I5(\iv_reg[15]_0 [1]),
        .O(\tr_reg[1] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[2]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[2]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[2]),
        .O(badr[1]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[2]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [2]),
        .O(a1bus_sr[2]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [2]),
        .I5(\iv_reg[15]_0 [2]),
        .O(\tr_reg[2] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[3]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[3]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[3]),
        .O(badr[2]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[3]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [3]),
        .O(a1bus_sr[3]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [3]),
        .I5(\iv_reg[15]_0 [3]),
        .O(\tr_reg[3] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[4]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[4]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[4]),
        .O(badr[3]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[4]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [4]),
        .O(a1bus_sr[4]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [4]),
        .I5(\iv_reg[15]_0 [4]),
        .O(\tr_reg[4]_1 ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[5]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[5]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[5]),
        .O(badr[4]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[5]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [5]),
        .O(a1bus_sr[5]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [5]),
        .I5(\iv_reg[15]_0 [5]),
        .O(\tr_reg[5] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[6]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[6]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[6]),
        .O(badr[5]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[6]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [6]),
        .O(a1bus_sr[6]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [6]),
        .I5(\iv_reg[15]_0 [6]),
        .O(\tr_reg[6] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[7]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[7]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[7]),
        .O(badr[6]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[7]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [7]),
        .O(a1bus_sr[7]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [7]),
        .I5(\iv_reg[15]_0 [7]),
        .O(\tr_reg[7] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[8]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[8]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[8]),
        .O(badr[7]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[8]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [8]),
        .O(a1bus_sr[8]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [8]),
        .I5(\iv_reg[15]_0 [8]),
        .O(\tr_reg[8] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[9]_INST_0 
       (.I0(\stat_reg[1]_5 [2]),
        .I1(\stat_reg[2]_5 ),
        .I2(a1bus_0[9]),
        .I3(\stat_reg[0]_48 ),
        .I4(a0bus_0[9]),
        .O(badr[8]));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[9]_INST_0_i_6 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_26_n_0 ),
        .I3(\stat_reg[2]_15 ),
        .I4(\stat_reg[2]_16 ),
        .I5(\sr_reg[15]_0 [9]),
        .O(a1bus_sr[9]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\tr_reg[15]_1 [9]),
        .I5(\iv_reg[15]_0 [9]),
        .O(\tr_reg[9] ));
  MUXF7 \badrx[15]_INST_0_i_1 
       (.I0(\badrx[15]_INST_0_i_2_n_0 ),
        .I1(\badrx[15]_INST_0_i_3_n_0 ),
        .O(\stat_reg[1]_4 ),
        .S(\stat_reg[0]_48 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \badrx[15]_INST_0_i_2 
       (.I0(tout__1_carry_i_22_0),
        .I1(ir1[11]),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(ir1[15]),
        .I4(\badrx[15]_INST_0_i_5_n_0 ),
        .I5(\badrx[15]_INST_0_i_6_n_0 ),
        .O(\badrx[15]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    \badrx[15]_INST_0_i_3 
       (.I0(ir0[12]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\badrx[15]_INST_0_i_7_n_0 ),
        .O(\badrx[15]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[15]_INST_0_i_5 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\badrx[15]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hBFFF)) 
    \badrx[15]_INST_0_i_6 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .O(\badrx[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \badrx[15]_INST_0_i_7 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(ir0[8]),
        .I2(ir0[15]),
        .I3(ir0[11]),
        .I4(\rgf_selc0_rn_wb_reg[0] [2]),
        .I5(rst_n_fl_reg_2),
        .O(\badrx[15]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[0]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\tr_reg[0]_0 ),
        .O(bbus_o[0]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[0]_INST_0_i_1 
       (.I0(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_3_n_0 ),
        .I2(bbus_o_0_sn_1),
        .I3(p_1_in3_in[0]),
        .I4(p_0_in2_in[0]),
        .I5(\bbus_o[0]_0 ),
        .O(\tr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFABAAAFAFFEFF)) 
    \bbus_o[0]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I4(\stat_reg[0]_7 ),
        .I5(ctl_selb0_0),
        .O(\bbus_o[0]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[0]_INST_0_i_22 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_0 [0]),
        .O(b0bus_sr[0]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[0]_INST_0_i_23 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20 [0]),
        .O(\grn_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[0]_INST_0_i_24 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20_0 [0]),
        .O(\grn_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[0]_INST_0_i_25 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21 [0]),
        .O(\grn_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[0]_INST_0_i_26 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21_0 [0]),
        .O(\grn_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[0]_INST_0_i_27 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22_0 [0]),
        .O(\grn_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[0]_INST_0_i_28 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[0]_INST_0_i_29 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23_0 [0]),
        .O(\grn_reg[0]_3 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[0]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[0]),
        .O(\bbus_o[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[0]_INST_0_i_30 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23 [0]),
        .O(\grn_reg[0]_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bbus_o[0]_INST_0_i_8 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .O(\bbus_o[0]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[10]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\bdatw[10]_0 ),
        .O(bbus_o[9]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[11]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(bdatw_11_sn_1),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[12]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(bdatw_12_sn_1),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[13]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(bbus_o_13_sn_1),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[14]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(bbus_o_14_sn_1),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[15]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\bdatw[15] ),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[1]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(bbus_o[1]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[1]_INST_0_i_1 
       (.I0(\bbus_o[1]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_3_n_0 ),
        .I2(bbus_o_1_sn_1),
        .I3(p_1_in3_in[1]),
        .I4(p_0_in2_in[1]),
        .I5(\bbus_o[1]_0 ),
        .O(\bbus_o[1]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEABFBFEFEABFB)) 
    \bbus_o[1]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I2(\stat_reg[0]_7 ),
        .I3(ir0[1]),
        .I4(ctl_selb0_0),
        .I5(ir0[0]),
        .O(\bbus_o[1]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[1]_INST_0_i_21 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_0 [1]),
        .O(b0bus_sr[1]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[1]_INST_0_i_22 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20 [1]),
        .O(\grn_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[1]_INST_0_i_23 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20_0 [1]),
        .O(\grn_reg[1]_7 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[1]_INST_0_i_24 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21 [1]),
        .O(\grn_reg[1]_5 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[1]_INST_0_i_25 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21_0 [1]),
        .O(\grn_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[1]_INST_0_i_26 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22_0 [1]),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[1]_INST_0_i_27 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[1]_INST_0_i_28 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23_0 [1]),
        .O(\grn_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[1]_INST_0_i_29 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23 [1]),
        .O(\grn_reg[1]_2 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[1]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[1]),
        .O(\bbus_o[1]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[2]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(bbus_o[2]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[2]_INST_0_i_1 
       (.I0(\bbus_o[2]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_3_n_0 ),
        .I2(bbus_o_2_sn_1),
        .I3(p_1_in3_in[2]),
        .I4(p_0_in2_in[2]),
        .I5(\bbus_o[2]_0 ),
        .O(\bbus_o[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFAEAAAFAFFBFF)) 
    \bbus_o[2]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(\bbus_o[2]_INST_0_i_8_n_0 ),
        .I2(ir0[2]),
        .I3(ir0[1]),
        .I4(\stat_reg[0]_7 ),
        .I5(ctl_selb0_0),
        .O(\bbus_o[2]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[2]_INST_0_i_22 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_0 [2]),
        .O(b0bus_sr[2]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[2]_INST_0_i_23 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20 [2]),
        .O(\grn_reg[2]_4 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[2]_INST_0_i_24 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20_0 [2]),
        .O(\grn_reg[2]_7 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[2]_INST_0_i_25 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21 [2]),
        .O(\grn_reg[2]_5 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[2]_INST_0_i_26 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21_0 [2]),
        .O(\grn_reg[2]_6 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[2]_INST_0_i_27 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22_0 [2]),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[2]_INST_0_i_28 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[2]_INST_0_i_29 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23_0 [2]),
        .O(\grn_reg[2]_3 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[2]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[2]),
        .O(\bbus_o[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[2]_INST_0_i_30 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23 [2]),
        .O(\grn_reg[2]_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bbus_o[2]_INST_0_i_8 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .O(\bbus_o[2]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[3]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(bbus_o[3]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[3]_INST_0_i_1 
       (.I0(\bbus_o[3]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_3_n_0 ),
        .I2(bbus_o_3_sn_1),
        .I3(p_1_in3_in[3]),
        .I4(p_0_in2_in[3]),
        .I5(\bbus_o[3]_0 ),
        .O(\bbus_o[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAFFBBAFFFAFEE)) 
    \bbus_o[3]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(\bbus_o[3]_INST_0_i_8_n_0 ),
        .I2(ir0[3]),
        .I3(\stat_reg[0]_7 ),
        .I4(ir0[2]),
        .I5(ctl_selb0_0),
        .O(\bbus_o[3]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[3]_INST_0_i_22 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_0 [3]),
        .O(b0bus_sr[3]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[3]_INST_0_i_23 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20 [3]),
        .O(\grn_reg[3]_4 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[3]_INST_0_i_24 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20_0 [3]),
        .O(\grn_reg[3]_7 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[3]_INST_0_i_25 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21 [3]),
        .O(\grn_reg[3]_5 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[3]_INST_0_i_26 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21_0 [3]),
        .O(\grn_reg[3]_6 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[3]_INST_0_i_27 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22_0 [3]),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[3]_INST_0_i_28 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[3]_INST_0_i_29 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23_0 [3]),
        .O(\grn_reg[3]_3 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[3]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[3]),
        .O(\bbus_o[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[3]_INST_0_i_30 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23 [3]),
        .O(\grn_reg[3]_2 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \bbus_o[3]_INST_0_i_8 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .O(\bbus_o[3]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[4]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\tr_reg[4] ),
        .O(bbus_o[4]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[4]_INST_0_i_1 
       (.I0(\bbus_o[4]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[13]_0 ),
        .I3(p_1_in3_in[4]),
        .I4(p_0_in2_in[4]),
        .I5(\rgf_c0bus_wb_reg[13]_1 ),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hAAFFBFAAEEFFBFAA)) 
    \bbus_o[4]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ir0[4]),
        .I3(\bbus_o[4]_INST_0_i_8_n_0 ),
        .I4(ctl_selb0_0),
        .I5(ir0[3]),
        .O(\bbus_o[4]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[4]_INST_0_i_24 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\sr_reg[15]_0 [4]),
        .O(b0bus_sr[4]));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bbus_o[4]_INST_0_i_25 
       (.I0(ctl_selb0_0),
        .I1(\stat_reg[0]_7 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[2]_17 ),
        .I4(ctl_selb0_rn[1]),
        .I5(ctl_selb0_rn[0]),
        .O(b0bus_sel_0[1]));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bbus_o[4]_INST_0_i_26 
       (.I0(ctl_selb0_0),
        .I1(\stat_reg[0]_7 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[2]_17 ),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(b0bus_sel_0[0]));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[4]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[4]),
        .O(\bbus_o[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[4]_INST_0_i_31 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20 [4]),
        .O(\grn_reg[4]_4 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[4]_INST_0_i_32 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_20_0 [4]),
        .O(\grn_reg[4]_7 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[4]_INST_0_i_35 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21 [4]),
        .O(\grn_reg[4]_5 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[4]_INST_0_i_36 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(\i_/bbus_o[0]_INST_0_i_18 ),
        .I5(\i_/bbus_o[4]_INST_0_i_21_0 [4]),
        .O(\grn_reg[4]_6 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[4]_INST_0_i_38 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(\stat_reg[2]_17 ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22_0 [4]),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[4]_INST_0_i_39 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[0]),
        .I3(\stat_reg[0]_21 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_22 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bbus_o[4]_INST_0_i_42 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I2(\sr_reg[5] ),
        .I3(\stat_reg[0]_22 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23_0 [4]),
        .O(\grn_reg[4]_3 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bbus_o[4]_INST_0_i_43 
       (.I0(\bbus_o[4]_INST_0_i_45_n_0 ),
        .I1(\sr_reg[5] ),
        .I2(ctl_selb0_rn[1]),
        .I3(\stat_reg[0]_23 ),
        .I4(bank_sel),
        .I5(\i_/bbus_o[4]_INST_0_i_23 [4]),
        .O(\grn_reg[4]_2 ));
  LUT6 #(
    .INIT(64'hFEFFFEFEFEFFFEFF)) 
    \bbus_o[4]_INST_0_i_45 
       (.I0(\bbus_o[4]_INST_0_i_48_n_0 ),
        .I1(\bdatw[15]_INST_0_i_60_n_0 ),
        .I2(\bdatw[15]_INST_0_i_67_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\bbus_o[4]_INST_0_i_49_n_0 ),
        .I5(\bdatw[15]_INST_0_i_64_n_0 ),
        .O(\bbus_o[4]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5F5F5F4F4F4FF)) 
    \bbus_o[4]_INST_0_i_46 
       (.I0(\bdatw[15]_INST_0_i_160_n_0 ),
        .I1(\bdatw[15]_INST_0_i_171_n_0 ),
        .I2(\bdatw[15]_INST_0_i_163_n_0 ),
        .I3(\bdatw[15]_INST_0_i_172_n_0 ),
        .I4(\bdatw[15]_INST_0_i_173_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\stat_reg[0]_32 ));
  LUT6 #(
    .INIT(64'hFF55FF54FF55FFFF)) 
    \bbus_o[4]_INST_0_i_47 
       (.I0(\bdatw[15]_INST_0_i_163_n_0 ),
        .I1(\bdatw[15]_INST_0_i_172_n_0 ),
        .I2(\bdatw[15]_INST_0_i_173_n_0 ),
        .I3(\bdatw[15]_INST_0_i_160_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\bdatw[15]_INST_0_i_171_n_0 ),
        .O(\stat_reg[0]_31 ));
  LUT6 #(
    .INIT(64'hFFFF7F7700000000)) 
    \bbus_o[4]_INST_0_i_48 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(\bdatw[15]_INST_0_i_142_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_50_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_51_n_0 ),
        .I5(ir0[12]),
        .O(\bbus_o[4]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF02)) 
    \bbus_o[4]_INST_0_i_49 
       (.I0(\bdatw[15]_INST_0_i_150_n_0 ),
        .I1(\bdatw[15]_INST_0_i_151_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_52_n_0 ),
        .I3(rst_n_fl_reg_2),
        .I4(\bbus_o[4]_INST_0_i_53_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_54_n_0 ),
        .O(\bbus_o[4]_INST_0_i_49_n_0 ));
  MUXF7 \bbus_o[4]_INST_0_i_50 
       (.I0(\bdatw[15]_INST_0_i_145_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_55_n_0 ),
        .O(\bbus_o[4]_INST_0_i_50_n_0 ),
        .S(ir0[11]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAA2AAAAA)) 
    \bbus_o[4]_INST_0_i_51 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[11]),
        .I5(\ccmd[4]_INST_0_i_20_n_0 ),
        .O(\bbus_o[4]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBFB0000)) 
    \bbus_o[4]_INST_0_i_52 
       (.I0(\bbus_o[4]_INST_0_i_56_n_0 ),
        .I1(ir0[9]),
        .I2(\bbus_o[4]_INST_0_i_57_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_58_n_0 ),
        .I4(ir0[11]),
        .I5(\bdatw[15]_INST_0_i_154_n_0 ),
        .O(\bbus_o[4]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFA959FFFF)) 
    \bbus_o[4]_INST_0_i_53 
       (.I0(ir0[11]),
        .I1(\sr_reg[15]_0 [4]),
        .I2(ir0[14]),
        .I3(\bbus_o[4]_INST_0_i_49_0 ),
        .I4(ir0[12]),
        .I5(ir0[13]),
        .O(\bbus_o[4]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h1110FFFF11101110)) 
    \bbus_o[4]_INST_0_i_54 
       (.I0(ir0[6]),
        .I1(\bdatw[15]_INST_0_i_223_n_0 ),
        .I2(\ccmd[4]_INST_0_i_12_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_59_n_0 ),
        .I4(\bdatw[15]_INST_0_i_148_n_0 ),
        .I5(ir0[13]),
        .O(\bbus_o[4]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055555501)) 
    \bbus_o[4]_INST_0_i_55 
       (.I0(\bdatw[15]_INST_0_i_224_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_60_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_61_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_62_n_0 ),
        .I4(\badr[15]_INST_0_i_274_n_0 ),
        .I5(\bdatw[15]_INST_0_i_225_n_0 ),
        .O(\bbus_o[4]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \bbus_o[4]_INST_0_i_56 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[5]),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(ir0[4]),
        .O(\bbus_o[4]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hD050)) 
    \bbus_o[4]_INST_0_i_57 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .O(\bbus_o[4]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h80888800)) 
    \bbus_o[4]_INST_0_i_58 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .I4(ir0[4]),
        .O(\bbus_o[4]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \bbus_o[4]_INST_0_i_59 
       (.I0(ir0[14]),
        .I1(ir0[13]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .O(\bbus_o[4]_INST_0_i_59_n_0 ));
  LUT3 #(
    .INIT(8'h62)) 
    \bbus_o[4]_INST_0_i_60 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .O(\bbus_o[4]_INST_0_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h56)) 
    \bbus_o[4]_INST_0_i_61 
       (.I0(ir0[6]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .O(\bbus_o[4]_INST_0_i_61_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \bbus_o[4]_INST_0_i_62 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\bbus_o[4]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \bbus_o[4]_INST_0_i_8 
       (.I0(\stat_reg[0]_7 ),
        .I1(ir0[2]),
        .I2(ir0[0]),
        .I3(ir0[3]),
        .I4(ir0[1]),
        .O(\bbus_o[4]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[5]_INST_0_i_18 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [5]),
        .O(b0bus_sr[5]));
  LUT6 #(
    .INIT(64'h5500405511004055)) 
    \bbus_o[5]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ir0[5]),
        .I3(\bbus_o[5]_INST_0_i_8_n_0 ),
        .I4(ctl_selb0_0),
        .I5(ir0[4]),
        .O(\stat_reg[0]_30 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[5]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[5]),
        .O(\stat_reg[0]_34 ));
  LUT5 #(
    .INIT(32'hFFFBFFFF)) 
    \bbus_o[5]_INST_0_i_8 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .I2(ir0[3]),
        .I3(\stat_reg[0]_7 ),
        .I4(ir0[2]),
        .O(\bbus_o[5]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[6]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(bbus_o_6_sn_1),
        .O(bbus_o[5]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[6]_INST_0_i_18 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [6]),
        .O(b0bus_sr[6]));
  LUT6 #(
    .INIT(64'h4455514000115140)) 
    \bbus_o[6]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ir0[6]),
        .I3(\bbus_o[6]_INST_0_i_8_n_0 ),
        .I4(ctl_selb0_0),
        .I5(ir0[5]),
        .O(\stat_reg[0]_29 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[6]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[6]),
        .O(\stat_reg[0]_35 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bbus_o[6]_INST_0_i_8 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[2]),
        .O(\bbus_o[6]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[7]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(bbus_o_7_sn_1),
        .O(bbus_o[6]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[7]_INST_0_i_18 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [7]),
        .O(b0bus_sr[7]));
  LUT6 #(
    .INIT(64'hAAFFBFAAEEFFBFAA)) 
    \bbus_o[7]_INST_0_i_2 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ir0[7]),
        .I3(\bbus_o[7]_INST_0_i_8_n_0 ),
        .I4(ctl_selb0_0),
        .I5(ir0[6]),
        .O(\stat_reg[0]_10 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bbus_o[7]_INST_0_i_3 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[7]),
        .O(\stat_reg[0]_36 ));
  LUT5 #(
    .INIT(32'hFFDFFFFF)) 
    \bbus_o[7]_INST_0_i_8 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(ir0[0]),
        .I3(\stat_reg[0]_7 ),
        .I4(ir0[2]),
        .O(\bbus_o[7]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[8]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\bdatw[8]_0 ),
        .O(bbus_o[7]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[9]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(bdatw_9_sn_1),
        .O(bbus_o[8]));
  MUXF7 \bcmd[0]_INST_0 
       (.I0(\bcmd[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_2_n_0 ),
        .O(\stat_reg[1]_5 [2]),
        .S(\stat_reg[0]_48 ));
  LUT6 #(
    .INIT(64'h0100010F01000100)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\bcmd[0]_INST_0_i_4_n_0 ),
        .I2(\bcmd[0]_INST_0_i_5_n_0 ),
        .I3(ir1[12]),
        .I4(\bcmd[0]_INST_0_i_6_n_0 ),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBDFBFBFFFDFBFBFF)) 
    \bcmd[0]_INST_0_i_10 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(ir0[5]),
        .O(\bcmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2A7FFF00)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(ir0[6]),
        .I1(ir0[3]),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .I5(\bcmd[1] ),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAA40AA44AA44AA44)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(ir0[10]),
        .I1(\bcmd[0]_INST_0_i_21_n_0 ),
        .I2(\bcmd[0]_INST_0_i_22_n_0 ),
        .I3(ir0[7]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\bcmd[0]_INST_0_i_23_n_0 ),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC0FF0000C000A0A0)) 
    \bcmd[0]_INST_0_i_13 
       (.I0(ir1[10]),
        .I1(ir1[3]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[8]),
        .I5(ir1[9]),
        .O(\bcmd[0]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[0]_INST_0_i_14 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\bcmd[0]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[0]_INST_0_i_15 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .O(\bcmd[0]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00100000)) 
    \bcmd[0]_INST_0_i_16 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(ir1[1]),
        .I3(ir1[3]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\bcmd[0]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[0]_INST_0_i_17 
       (.I0(ir1[7]),
        .I1(ir1[5]),
        .I2(ir1[8]),
        .I3(ir1[4]),
        .O(\bcmd[0]_INST_0_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_18 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[13]),
        .O(\bcmd[0]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_19 
       (.I0(ir0[6]),
        .I1(ir0[5]),
        .O(\bcmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00AE00AE00AE0000)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(\bcmd[0]_INST_0_i_8_n_0 ),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .I2(\bcmd[0]_INST_0_i_10_n_0 ),
        .I3(\bcmd[0]_INST_0_i_11_n_0 ),
        .I4(ir0[8]),
        .I5(\bcmd[0]_INST_0_i_12_n_0 ),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_20 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .O(\bcmd[0]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[0]_INST_0_i_21 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .O(\bcmd[0]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_22 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .O(\bcmd[0]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \bcmd[0]_INST_0_i_23 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[2]),
        .I3(ir0[1]),
        .O(\bcmd[0]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .O(\bcmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFBF6BFFFFBFEBFF)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(ir1[6]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[5]),
        .O(\bcmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h45FF45FFFFFF45FF)) 
    \bcmd[0]_INST_0_i_5 
       (.I0(\bcmd[0]_INST_0_i_13_n_0 ),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(\bcmd[0]_INST_0_i_15_n_0 ),
        .I3(\bcmd[1]_0 ),
        .I4(\bcmd[0]_INST_0_i_16_n_0 ),
        .I5(\bcmd[0]_INST_0_i_17_n_0 ),
        .O(\bcmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(ir1[14]),
        .I1(ir1[11]),
        .I2(ir1[13]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(ir1[2]),
        .O(\bcmd[0]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .O(\bcmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(\bcmd[0]_INST_0_i_18_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[4]),
        .I3(\bcmd[0]_INST_0_i_19_n_0 ),
        .I4(ir0[14]),
        .I5(\bcmd[0]_INST_0_i_20_n_0 ),
        .O(\bcmd[0]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[0]_INST_0_i_9 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(ir0[13]),
        .O(\bcmd[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4500450045FF4500)) 
    \bcmd[1]_INST_0 
       (.I0(\bcmd[1] ),
        .I1(\bcmd[1]_INST_0_i_2_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\stat_reg[0]_48 ),
        .I4(\bcmd[1]_0 ),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\stat_reg[2]_5 ));
  LUT6 #(
    .INIT(64'hFFFFFBFFFBFFFFFF)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(\bcmd[1]_INST_0_i_14_n_0 ),
        .I1(ir0[6]),
        .I2(rst_n_fl_reg_2),
        .I3(ir0[12]),
        .I4(ir0[9]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFBFFFBFFFFFF)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(\bcmd[1]_INST_0_i_16_n_0 ),
        .I1(ir1[12]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\bcmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hEEFFFFFFEEFFFFEF)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(\bcmd[1]_INST_0_i_17_n_0 ),
        .I1(\bcmd[1]_INST_0_i_18_n_0 ),
        .I2(ir1[0]),
        .I3(ir1[7]),
        .I4(ir1[3]),
        .I5(ir1[1]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD0000000D000D000)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(ir0[9]),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(ir0[3]),
        .I5(ir0[5]),
        .O(\bcmd[1]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .O(rst_n_fl_reg_2));
  LUT6 #(
    .INIT(64'h7A5FFF5F5FFF5FFF)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(ir1[8]),
        .I1(\bcmd[1]_INST_0_i_19_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .I4(ir1[7]),
        .I5(ir1[11]),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFFFFFFFF7E)) 
    \bcmd[1]_INST_0_i_17 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .I4(ir1[9]),
        .I5(ir1[10]),
        .O(\bcmd[1]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFF3FFFFFFFFFFFE)) 
    \bcmd[1]_INST_0_i_18 
       (.I0(ir1[2]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(\stat[2]_i_10__0_n_0 ),
        .I4(ir1[8]),
        .I5(ir1[7]),
        .O(\bcmd[1]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_19 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .O(\bcmd[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000FE)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(fch_irq_req),
        .I2(\bcmd[1]_INST_0_i_6_n_0 ),
        .I3(\bcmd[1]_INST_0_i_7_n_0 ),
        .I4(\bcmd[1]_INST_0_i_8_n_0 ),
        .I5(\bcmd[1]_INST_0_i_9_n_0 ),
        .O(\bcmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1FF79FFF)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[7]),
        .I5(\bcmd[1]_INST_0_i_10_n_0 ),
        .O(\bcmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8AAAAAAAA888A)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(fch_irq_req),
        .I4(ir1[11]),
        .I5(ir1[12]),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .O(\bcmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF3FFE3FFF)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(ir0[1]),
        .I1(ir0[8]),
        .I2(ir0[3]),
        .I3(ir0[7]),
        .I4(ir0[0]),
        .I5(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFE7FFE)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\bcmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h3EFFFFFFFFFFFF3E)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(ir0[2]),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .I5(ir0[13]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  MUXF7 \bcmd[2]_INST_0 
       (.I0(\bcmd[2]_INST_0_i_2_n_0 ),
        .I1(\bcmd[2]_INST_0_i_3_n_0 ),
        .O(\stat_reg[1]_5 [1]),
        .S(\stat_reg[0]_48 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[2]_INST_0_i_11 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\bcmd[2]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(\bcmd[2]_INST_0_i_4_n_0 ),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[7]),
        .I4(\read_cyc_reg[1] ),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\bcmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(\bcmd[2]_INST_0_i_8_n_0 ),
        .I3(\bcmd[2]_INST_0_i_9_n_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(\bcmd[2]_INST_0_i_11_n_0 ),
        .O(\bcmd[2]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF77F)) 
    \bcmd[2]_INST_0_i_4 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(ir1[11]),
        .O(\bcmd[2]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[2]_INST_0_i_5 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .O(\bcmd[2]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[2]_INST_0_i_7 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .O(\bcmd[2]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[2]_INST_0_i_8 
       (.I0(ir0[9]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\bcmd[2]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[2]_INST_0_i_9 
       (.I0(ir0[13]),
        .I1(ir0[12]),
        .O(\bcmd[2]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[0]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .O(bdatw[0]));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[10]_INST_0 
       (.I0(\bdatw[10]_0 ),
        .I1(\stat_reg[0]_48 ),
        .I2(bdatw_10_sn_1),
        .I3(\bcmd[2]_INST_0_0 ),
        .I4(\bdatw[10]_INST_0_i_3_n_0 ),
        .I5(\bcmd[1]_INST_0_0 ),
        .O(bdatw[10]));
  LUT6 #(
    .INIT(64'h808000002A2AAA00)) 
    \bdatw[10]_INST_0_i_10 
       (.I0(\stat_reg[0]_11 ),
        .I1(\bdatw[14]_INST_0_i_29_n_0 ),
        .I2(\bdatw[10]_INST_0_i_29_n_0 ),
        .I3(ir1[9]),
        .I4(ctl_selb1_0),
        .I5(\stat_reg[0]_12 ),
        .O(rst_n_fl_reg_3));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_11 
       (.I0(eir[10]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_2));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \bdatw[10]_INST_0_i_16 
       (.I0(\bdatw[10]_INST_0_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_9_0 ),
        .I2(b1bus_b02[2]),
        .I3(\rgf_c1bus_wb[5]_i_9_1 ),
        .I4(\rgf_c1bus_wb[5]_i_9_2 ),
        .I5(\bdatw[10]_INST_0_i_45_n_0 ),
        .O(\bdatw[10]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[10]_INST_0_i_17 
       (.I0(ir0[2]),
        .I1(ir0[0]),
        .O(\bdatw[10]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[10]_INST_0_i_18 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .O(\bdatw[10]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[10]_INST_0_i_28 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [10]),
        .O(b0bus_sr[10]));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[10]_INST_0_i_29 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .O(\bdatw[10]_INST_0_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_48 ),
        .I2(\bdatw[10]_INST_0_i_16_n_0 ),
        .O(\bdatw[10]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[10]_INST_0_i_39 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [10]),
        .O(b1bus_sr[10]));
  LUT6 #(
    .INIT(64'h4044401140444044)) 
    \bdatw[10]_INST_0_i_4 
       (.I0(\sr_reg[5] ),
        .I1(ctl_selb0_0),
        .I2(ir0[9]),
        .I3(\stat_reg[0]_7 ),
        .I4(\bdatw[10]_INST_0_i_17_n_0 ),
        .I5(\bdatw[10]_INST_0_i_18_n_0 ),
        .O(\stat_reg[0]_6 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_40 
       (.I0(eir[2]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(\bdatw[10]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \bdatw[10]_INST_0_i_45 
       (.I0(ir1[1]),
        .I1(ctl_selb1_0),
        .I2(\bdatw[10]_INST_0_i_70_n_0 ),
        .I3(\stat_reg[0]_12 ),
        .I4(ir1[2]),
        .I5(\stat_reg[0]_11 ),
        .O(\bdatw[10]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[10]_INST_0_i_5 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[10]),
        .O(\stat_reg[0]_39 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[10]_INST_0_i_64 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_117_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_0 [2]),
        .O(b1bus_sr[2]));
  LUT4 #(
    .INIT(16'h0004)) 
    \bdatw[10]_INST_0_i_70 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(ir1[2]),
        .I3(ir1[0]),
        .O(\bdatw[10]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bdatw[10]_INST_0_i_73 
       (.I0(\stat_reg[0]_19 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [2]),
        .O(\sr_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bdatw[10]_INST_0_i_74 
       (.I0(\stat_reg[0]_20 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_64 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[11]_INST_0 
       (.I0(bdatw_11_sn_1),
        .I1(\stat_reg[0]_48 ),
        .I2(\bdatw[11]_0 ),
        .I3(\bcmd[2]_INST_0_0 ),
        .I4(\bdatw[11]_INST_0_i_3_n_0 ),
        .I5(\bcmd[1]_INST_0_0 ),
        .O(bdatw[11]));
  LUT6 #(
    .INIT(64'h08080000A2A2AA00)) 
    \bdatw[11]_INST_0_i_10 
       (.I0(\stat_reg[0]_11 ),
        .I1(\bdatw[11]_INST_0_i_28_n_0 ),
        .I2(\bdatw[11]_INST_0_i_29_n_0 ),
        .I3(ir1[10]),
        .I4(ctl_selb1_0),
        .I5(\stat_reg[0]_12 ),
        .O(rst_n_fl_reg_4));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_11 
       (.I0(eir[11]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_1));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[11]_INST_0_i_16 
       (.I0(\bdatw[11]_INST_0_i_40_n_0 ),
        .I1(\bdatw[11]_INST_0_i_41_n_0 ),
        .I2(\sr[4]_i_102_1 ),
        .I3(b1bus_b02[3]),
        .I4(\sr[4]_i_102_2 ),
        .I5(\sr[4]_i_102_3 ),
        .O(\bdatw[11]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_17 
       (.I0(ir0[1]),
        .I1(ir0[2]),
        .O(\bdatw[11]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[11]_INST_0_i_27 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [11]),
        .O(b0bus_sr[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_28 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .O(\bdatw[11]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[11]_INST_0_i_29 
       (.I0(ir1[2]),
        .I1(ir1[1]),
        .O(\bdatw[11]_INST_0_i_29_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[11]_INST_0_i_3 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_48 ),
        .I2(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\bdatw[11]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_39 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [11]),
        .O(b1bus_sr[11]));
  LUT6 #(
    .INIT(64'hBAAAEFFFFEEEEFFF)) 
    \bdatw[11]_INST_0_i_4 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(\bdatw[11]_INST_0_i_17_n_0 ),
        .I3(\bdatw[15]_INST_0_i_19_n_0 ),
        .I4(ctl_selb0_0),
        .I5(ir0[10]),
        .O(\stat_reg[0]_28 ));
  LUT6 #(
    .INIT(64'h0CF13FF1FFFFFFFF)) 
    \bdatw[11]_INST_0_i_40 
       (.I0(ir1[2]),
        .I1(ctl_selb1_0),
        .I2(\bdatw[11]_INST_0_i_58_n_0 ),
        .I3(\stat_reg[0]_12 ),
        .I4(ir1[3]),
        .I5(\stat_reg[0]_11 ),
        .O(\bdatw[11]_INST_0_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_41 
       (.I0(eir[3]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(\bdatw[11]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[11]_INST_0_i_5 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[11]),
        .O(\stat_reg[0]_40 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[11]_INST_0_i_58 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .I3(ir1[2]),
        .O(\bdatw[11]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[11]_INST_0_i_65 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_117_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_0 [3]),
        .O(b1bus_sr[3]));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bdatw[11]_INST_0_i_73 
       (.I0(\stat_reg[0]_19 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [3]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bdatw[11]_INST_0_i_74 
       (.I0(\stat_reg[0]_20 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_64 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[12]_INST_0 
       (.I0(bdatw_12_sn_1),
        .I1(\stat_reg[0]_48 ),
        .I2(\bdatw[12]_0 ),
        .I3(\bcmd[2]_INST_0_0 ),
        .I4(\bdatw[12]_INST_0_i_3_n_0 ),
        .I5(\bcmd[1]_INST_0_0 ),
        .O(bdatw[12]));
  LUT6 #(
    .INIT(64'h2220828022202220)) 
    \bdatw[12]_INST_0_i_10 
       (.I0(\stat_reg[0]_11 ),
        .I1(\stat_reg[0]_12 ),
        .I2(ctl_selb1_0),
        .I3(ir1[10]),
        .I4(\bdatw[13]_INST_0_i_28_n_0 ),
        .I5(\bdatw[14]_INST_0_i_30_n_0 ),
        .O(\stat_reg[0]_13 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[12]_INST_0_i_11 
       (.I0(eir[12]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(rst_n_fl_reg_8));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[12]_INST_0_i_16 
       (.I0(\bdatw[12]_INST_0_i_38_n_0 ),
        .I1(\bdatw[12]_INST_0_i_39_n_0 ),
        .I2(\rgf_c1bus_wb_reg[13]_3 ),
        .I3(b1bus_b02[4]),
        .I4(\rgf_c1bus_wb_reg[13]_4 ),
        .I5(\rgf_c1bus_wb_reg[13]_5 ),
        .O(\tr_reg[4]_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[12]_INST_0_i_17 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(ir0[2]),
        .I3(ir0[0]),
        .O(\bdatw[12]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[12]_INST_0_i_27 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [12]),
        .O(b0bus_sr[12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(\tr_reg[4] ),
        .I1(\stat_reg[0]_48 ),
        .I2(\tr_reg[4]_0 ),
        .O(\bdatw[12]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_37 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [12]),
        .O(b1bus_sr[12]));
  LUT6 #(
    .INIT(64'h0CF13FF1FFFFFFFF)) 
    \bdatw[12]_INST_0_i_38 
       (.I0(ir1[3]),
        .I1(ctl_selb1_0),
        .I2(\bdatw[12]_INST_0_i_56_n_0 ),
        .I3(\stat_reg[0]_12 ),
        .I4(ir1[4]),
        .I5(\stat_reg[0]_11 ),
        .O(\bdatw[12]_INST_0_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[12]_INST_0_i_39 
       (.I0(eir[4]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(\bdatw[12]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hBAEFFEEF)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(\bdatw[12]_INST_0_i_17_n_0 ),
        .I3(ctl_selb0_0),
        .I4(ir0[10]),
        .O(\stat_reg[0]_27 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[12]_INST_0_i_5 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[12]),
        .O(\stat_reg[0]_41 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[12]_INST_0_i_56 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .O(\bdatw[12]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[12]_INST_0_i_63 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_117_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_0 [4]),
        .O(b1bus_sr[4]));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bdatw[12]_INST_0_i_71 
       (.I0(\stat_reg[0]_19 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [4]),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bdatw[12]_INST_0_i_72 
       (.I0(\stat_reg[0]_20 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_64 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h202000008A8AAA00)) 
    \bdatw[13]_INST_0_i_10 
       (.I0(\stat_reg[0]_11 ),
        .I1(\bdatw[13]_INST_0_i_28_n_0 ),
        .I2(\bdatw[13]_INST_0_i_29_n_0 ),
        .I3(ir1[10]),
        .I4(ctl_selb1_0),
        .I5(\stat_reg[0]_12 ),
        .O(rst_n_fl_reg_5));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_11 
       (.I0(eir[13]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(rst_n_fl_reg_7));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_17 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .O(\bdatw[13]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[13]_INST_0_i_27 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [13]),
        .O(b0bus_sr[13]));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[13]_INST_0_i_28 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .O(\bdatw[13]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[13]_INST_0_i_29 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .O(\bdatw[13]_INST_0_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[13]_INST_0_i_39 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [13]),
        .O(b1bus_sr[13]));
  LUT6 #(
    .INIT(64'hBAAAEFFFFEEEEFFF)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(\bdatw[13]_INST_0_i_17_n_0 ),
        .I3(\bdatw[14]_INST_0_i_17_n_0 ),
        .I4(ctl_selb0_0),
        .I5(ir0[10]),
        .O(\stat_reg[0]_26 ));
  LUT6 #(
    .INIT(64'hAA0A08A8A00008A8)) 
    \bdatw[13]_INST_0_i_40 
       (.I0(\stat_reg[0]_11 ),
        .I1(ir1[4]),
        .I2(ctl_selb1_0),
        .I3(\bdatw[13]_INST_0_i_58_n_0 ),
        .I4(\stat_reg[0]_12 ),
        .I5(ir1[5]),
        .O(rst_n_fl_reg_10));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_41 
       (.I0(eir[5]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_7));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[13]_INST_0_i_5 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[13]),
        .O(\stat_reg[0]_42 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[13]_INST_0_i_58 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .I2(ir1[2]),
        .I3(ir1[0]),
        .O(\bdatw[13]_INST_0_i_58_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[13]_INST_0_i_68 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [5]),
        .O(b1bus_sr[5]));
  LUT6 #(
    .INIT(64'h808000002A2AAA00)) 
    \bdatw[14]_INST_0_i_10 
       (.I0(\stat_reg[0]_11 ),
        .I1(\bdatw[14]_INST_0_i_29_n_0 ),
        .I2(\bdatw[14]_INST_0_i_30_n_0 ),
        .I3(ir1[10]),
        .I4(ctl_selb1_0),
        .I5(\stat_reg[0]_12 ),
        .O(rst_n_fl_reg_6));
  LUT5 #(
    .INIT(32'h2A020000)) 
    \bdatw[14]_INST_0_i_105 
       (.I0(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[1]),
        .I3(ir1[0]),
        .I4(ir1[2]),
        .O(\bdatw[14]_INST_0_i_105_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4444FFF4)) 
    \bdatw[14]_INST_0_i_106 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_5_0 ),
        .I2(rst_n_fl_reg_9),
        .I3(\bdatw[15]_INST_0_i_252_n_0 ),
        .I4(\bdatw[14]_INST_0_i_109_n_0 ),
        .I5(\bdatw[14]_INST_0_i_110_n_0 ),
        .O(\bdatw[14]_INST_0_i_106_n_0 ));
  LUT6 #(
    .INIT(64'h55555555FFDFFFFF)) 
    \bdatw[14]_INST_0_i_107 
       (.I0(\read_cyc_reg[1] ),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(\bcmd[0]_INST_0_i_7_n_0 ),
        .I3(\bdatw[15]_INST_0_i_199_n_0 ),
        .I4(\badr[15]_INST_0_i_70_n_0 ),
        .I5(\bdatw[15]_INST_0_i_185_n_0 ),
        .O(\bdatw[14]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1FFFFFFFFFFF1)) 
    \bdatw[14]_INST_0_i_108 
       (.I0(\stat[1]_i_11__0_n_0 ),
        .I1(\stat[2]_i_9__0_n_0 ),
        .I2(\bdatw[15]_INST_0_i_248_n_0 ),
        .I3(\bdatw[14]_INST_0_i_111_n_0 ),
        .I4(ir1[7]),
        .I5(ir1[10]),
        .O(\bdatw[14]_INST_0_i_108_n_0 ));
  LUT4 #(
    .INIT(16'hFFF7)) 
    \bdatw[14]_INST_0_i_109 
       (.I0(ir1[13]),
        .I1(ir1[14]),
        .I2(ir1[6]),
        .I3(ir1[8]),
        .O(\bdatw[14]_INST_0_i_109_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_11 
       (.I0(eir[14]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_0));
  LUT4 #(
    .INIT(16'h0802)) 
    \bdatw[14]_INST_0_i_110 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(ir1[14]),
        .I3(\sr_reg[15]_0 [7]),
        .O(\bdatw[14]_INST_0_i_110_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[14]_INST_0_i_111 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .O(\bdatw[14]_INST_0_i_111_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_17 
       (.I0(ir0[3]),
        .I1(ir0[2]),
        .O(\bdatw[14]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_18 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .O(\bdatw[14]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[14]_INST_0_i_28 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [14]),
        .O(b0bus_sr[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_29 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .O(\bdatw[14]_INST_0_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_30 
       (.I0(ir1[2]),
        .I1(ir1[0]),
        .O(\bdatw[14]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBAAAEFFFFEEEEFFF)) 
    \bdatw[14]_INST_0_i_4 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(\bdatw[14]_INST_0_i_17_n_0 ),
        .I3(\bdatw[14]_INST_0_i_18_n_0 ),
        .I4(ctl_selb0_0),
        .I5(ir0[10]),
        .O(\stat_reg[0]_25 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_44 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [14]),
        .O(b1bus_sr[14]));
  LUT6 #(
    .INIT(64'h2A2A8A8020208A80)) 
    \bdatw[14]_INST_0_i_45 
       (.I0(\stat_reg[0]_11 ),
        .I1(\bdatw[14]_INST_0_i_77_n_0 ),
        .I2(ctl_selb1_0),
        .I3(ir1[5]),
        .I4(\stat_reg[0]_12 ),
        .I5(ir1[6]),
        .O(rst_n_fl_reg_11));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_46 
       (.I0(eir[6]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_6));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[14]_INST_0_i_5 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[14]),
        .O(\stat_reg[0]_43 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFABFFFF)) 
    \bdatw[14]_INST_0_i_59 
       (.I0(ctl_selb1_rn[2]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\bdatw[14]_INST_0_i_89_n_0 ),
        .I3(\bdatw[14]_INST_0_i_90_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\stat_reg[0]_11 ),
        .O(\stat_reg[0]_19 ));
  LUT6 #(
    .INIT(64'hFFBFFFBFFFBBFFFF)) 
    \bdatw[14]_INST_0_i_60 
       (.I0(\stat_reg[0]_11 ),
        .I1(ctl_selb1_0),
        .I2(\bdatw[15]_INST_0_i_99_n_0 ),
        .I3(ir1[15]),
        .I4(\bdatw[14]_INST_0_i_89_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\stat_reg[0]_20 ));
  LUT4 #(
    .INIT(16'hFBFF)) 
    \bdatw[14]_INST_0_i_77 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .O(\bdatw[14]_INST_0_i_77_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_87 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [6]),
        .O(b1bus_sr[6]));
  LUT6 #(
    .INIT(64'h555555FDFFFFFFFF)) 
    \bdatw[14]_INST_0_i_88 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_205_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\bdatw[15]_INST_0_i_204_n_0 ),
        .I4(\bdatw[14]_INST_0_i_105_n_0 ),
        .I5(\bcmd[1]_0 ),
        .O(\stat_reg[0]_47 ));
  LUT6 #(
    .INIT(64'h00000000BABABABB)) 
    \bdatw[14]_INST_0_i_89 
       (.I0(\bdatw[14]_INST_0_i_106_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[15]_INST_0_i_182_n_0 ),
        .I3(\bdatw[15]_INST_0_i_181_n_0 ),
        .I4(\bdatw[15]_INST_0_i_180_n_0 ),
        .I5(\bdatw[14]_INST_0_i_107_n_0 ),
        .O(\bdatw[14]_INST_0_i_89_n_0 ));
  LUT5 #(
    .INIT(32'hFFFBAAAA)) 
    \bdatw[14]_INST_0_i_90 
       (.I0(ir1[15]),
        .I1(\bdatw[15]_INST_0_i_177_n_0 ),
        .I2(\bdatw[14]_INST_0_i_108_n_0 ),
        .I3(\bdatw[15]_INST_0_i_179_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\bdatw[14]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[15]_INST_0 
       (.I0(\bdatw[15] ),
        .I1(\stat_reg[0]_48 ),
        .I2(fch_leir_nir_reg),
        .I3(\bcmd[2]_INST_0_0 ),
        .I4(\bdatw[15]_0 ),
        .I5(\bcmd[1]_INST_0_0 ),
        .O(bdatw[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00F1)) 
    \bdatw[15]_INST_0_i_100 
       (.I0(\bdatw[15]_INST_0_i_180_n_0 ),
        .I1(\bdatw[15]_INST_0_i_181_n_0 ),
        .I2(\bdatw[15]_INST_0_i_182_n_0 ),
        .I3(\bcmd[0]_INST_0_i_3_n_0 ),
        .I4(\bdatw[15]_INST_0_i_183_n_0 ),
        .I5(\bdatw[15]_INST_0_i_184_n_0 ),
        .O(\bdatw[15]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAEAAAA)) 
    \bdatw[15]_INST_0_i_101 
       (.I0(\bdatw[15]_INST_0_i_185_n_0 ),
        .I1(\badr[15]_INST_0_i_70_n_0 ),
        .I2(\bdatw[15]_INST_0_i_186_n_0 ),
        .I3(ir1[13]),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(\bcmd[0]_INST_0_i_14_n_0 ),
        .O(\bdatw[15]_INST_0_i_101_n_0 ));
  LUT6 #(
    .INIT(64'h55757757FFFFFFFF)) 
    \bdatw[15]_INST_0_i_103 
       (.I0(\bdatw[15]_INST_0_i_187_n_0 ),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(\sr_reg[15]_0 [5]),
        .I4(ir1[11]),
        .I5(\rgf_selc1_wb[1]_i_5_0 ),
        .O(\bdatw[15]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA88AAAAA)) 
    \bdatw[15]_INST_0_i_104 
       (.I0(ir1[14]),
        .I1(\bdatw[15]_INST_0_i_188_n_0 ),
        .I2(ir1[5]),
        .I3(ir1[4]),
        .I4(ir1[7]),
        .I5(\bdatw[15]_INST_0_i_189_n_0 ),
        .O(\bdatw[15]_INST_0_i_104_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAFBEFEFE)) 
    \bdatw[15]_INST_0_i_105 
       (.I0(\bdatw[15]_INST_0_i_187_n_0 ),
        .I1(ir1[14]),
        .I2(ir1[11]),
        .I3(\sr_reg[15]_0 [7]),
        .I4(ir1[12]),
        .I5(ir1[15]),
        .O(\bdatw[15]_INST_0_i_105_n_0 ));
  LUT6 #(
    .INIT(64'hBBBB0A00AAAA0B00)) 
    \bdatw[15]_INST_0_i_106 
       (.I0(\bdatw[15]_INST_0_i_190_n_0 ),
        .I1(\bdatw[15]_INST_0_i_191_n_0 ),
        .I2(ir1[11]),
        .I3(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\bdatw[15]_INST_0_i_106_n_0 ));
  LUT6 #(
    .INIT(64'h888888888888888A)) 
    \bdatw[15]_INST_0_i_107 
       (.I0(ir1[11]),
        .I1(\bdatw[15]_INST_0_i_192_n_0 ),
        .I2(\bdatw[15]_INST_0_i_193_n_0 ),
        .I3(\bdatw[15]_INST_0_i_194_n_0 ),
        .I4(\bdatw[15]_INST_0_i_195_n_0 ),
        .I5(\bdatw[15]_INST_0_i_196_n_0 ),
        .O(\bdatw[15]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFAAAAAAAA)) 
    \bdatw[15]_INST_0_i_108 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I2(\bdatw[15]_INST_0_i_197_n_0 ),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\bdatw[15]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000EA0000)) 
    \bdatw[15]_INST_0_i_109 
       (.I0(\bdatw[15]_INST_0_i_198_n_0 ),
        .I1(fch_irq_req),
        .I2(\bdatw[9]_INST_0_i_69_n_0 ),
        .I3(\bcmd[0]_INST_0_i_14_n_0 ),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(\bdatw[15]_INST_0_i_199_n_0 ),
        .O(\bdatw[15]_INST_0_i_109_n_0 ));
  LUT6 #(
    .INIT(64'h00000008AA00AA08)) 
    \bdatw[15]_INST_0_i_114 
       (.I0(\bcmd[1]_0 ),
        .I1(ir1[12]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\bdatw[15]_INST_0_i_202_n_0 ),
        .I5(\bdatw[15]_INST_0_i_203_n_0 ),
        .O(ctl_selb1_rn[1]));
  LUT6 #(
    .INIT(64'hAA80AA80AA80AAAA)) 
    \bdatw[15]_INST_0_i_115 
       (.I0(\bcmd[1]_0 ),
        .I1(\badr[15]_INST_0_i_70_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I3(\bdatw[15]_INST_0_i_204_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\bdatw[15]_INST_0_i_205_n_0 ),
        .O(ctl_selb1_rn[0]));
  LUT6 #(
    .INIT(64'hFFAEAEAEAAAAAAAA)) 
    \bdatw[15]_INST_0_i_116 
       (.I0(\bdatw[15]_INST_0_i_206_n_0 ),
        .I1(\badr[15]_INST_0_i_90_n_0 ),
        .I2(\bdatw[15]_INST_0_i_207_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I4(\bdatw[15]_INST_0_i_208_n_0 ),
        .I5(\bdatw[15]_INST_0_i_209_n_0 ),
        .O(ctl_selb1_rn[2]));
  LUT3 #(
    .INIT(8'hBF)) 
    \bdatw[15]_INST_0_i_117 
       (.I0(\stat_reg[0]_11 ),
        .I1(\stat_reg[0]_12 ),
        .I2(ctl_selb1_0),
        .O(\bdatw[15]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \bdatw[15]_INST_0_i_118 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_0),
        .I4(\stat_reg[0]_12 ),
        .I5(\stat_reg[0]_11 ),
        .O(b1bus_sel_cr[5]));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \bdatw[15]_INST_0_i_119 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_0),
        .I4(\stat_reg[0]_12 ),
        .I5(\stat_reg[0]_11 ),
        .O(b1bus_sel_cr[2]));
  LUT6 #(
    .INIT(64'h37333333F7FFFFFF)) 
    \bdatw[15]_INST_0_i_12 
       (.I0(\stat_reg[0]_12 ),
        .I1(\stat_reg[0]_11 ),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(ir1[1]),
        .I4(ir1[2]),
        .I5(\bdatw[15]_INST_0_i_41_n_0 ),
        .O(\bdatw[15]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \bdatw[15]_INST_0_i_120 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[2]),
        .I2(ctl_selb1_rn[0]),
        .I3(ctl_selb1_0),
        .I4(\stat_reg[0]_12 ),
        .I5(\stat_reg[0]_11 ),
        .O(b1bus_sel_cr[1]));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[15]_INST_0_i_129 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(ir1[2]),
        .I3(ir1[0]),
        .O(\bdatw[15]_INST_0_i_129_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bdatw[15]_INST_0_i_13 
       (.I0(\stat_reg[0]_12 ),
        .I1(ctl_selb1_0),
        .I2(\stat_reg[0]_11 ),
        .O(\bdatw[15]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_139 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [7]),
        .O(b1bus_sr[7]));
  LUT6 #(
    .INIT(64'h0000000008800000)) 
    \bdatw[15]_INST_0_i_140 
       (.I0(ir0[9]),
        .I1(\ccmd[3]_INST_0_i_20_n_0 ),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[10]),
        .I5(ir0[6]),
        .O(\bdatw[15]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAEAEAEAEAEAEA)) 
    \bdatw[15]_INST_0_i_141 
       (.I0(\bdatw[15]_INST_0_i_222_n_0 ),
        .I1(fch_irq_req),
        .I2(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I3(\ccmd[4]_INST_0_i_13_n_0 ),
        .I4(ir0[0]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\bdatw[15]_INST_0_i_141_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200003032)) 
    \bdatw[15]_INST_0_i_142 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[10]),
        .I3(ir0[6]),
        .I4(\bdatw[15]_INST_0_i_223_n_0 ),
        .I5(ir0[9]),
        .O(\bdatw[15]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF9DFFBD)) 
    \bdatw[15]_INST_0_i_143 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(\badr[15]_INST_0_i_274_n_0 ),
        .I4(ir0[6]),
        .I5(\bdatw[15]_INST_0_i_224_n_0 ),
        .O(\bdatw[15]_INST_0_i_143_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABBBAABBABAA)) 
    \bdatw[15]_INST_0_i_144 
       (.I0(\bdatw[15]_INST_0_i_225_n_0 ),
        .I1(\badr[15]_INST_0_i_274_n_0 ),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[6]),
        .I5(ir0[3]),
        .O(\bdatw[15]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF07F7FFFFFFFF)) 
    \bdatw[15]_INST_0_i_145 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(crdy),
        .I2(ir0[8]),
        .I3(ir0[10]),
        .I4(\bdatw[15]_INST_0_i_226_n_0 ),
        .I5(ir0[6]),
        .O(\bdatw[15]_INST_0_i_145_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0A00CF30)) 
    \bdatw[15]_INST_0_i_146 
       (.I0(\sr_reg[15]_0 [6]),
        .I1(\sr_reg[15]_0 [5]),
        .I2(ir0[14]),
        .I3(ir0[11]),
        .I4(ir0[13]),
        .I5(ir0[12]),
        .O(\bdatw[15]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FFF7FFF7)) 
    \bdatw[15]_INST_0_i_147 
       (.I0(\bdatw[15]_INST_0_i_227_n_0 ),
        .I1(\badr[15]_INST_0_i_195_n_0 ),
        .I2(\bcmd[0]_INST_0_i_22_n_0 ),
        .I3(\badr[15]_INST_0_i_264_n_0 ),
        .I4(\sr_reg[15]_0 [6]),
        .I5(ir0[13]),
        .O(\bdatw[15]_INST_0_i_147_n_0 ));
  LUT3 #(
    .INIT(8'hDE)) 
    \bdatw[15]_INST_0_i_148 
       (.I0(\sr_reg[15]_0 [7]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .O(\bdatw[15]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000F10000)) 
    \bdatw[15]_INST_0_i_149 
       (.I0(rst_n_fl_reg_2),
        .I1(\ccmd[4]_INST_0_i_20_n_0 ),
        .I2(\ccmd[4]_INST_0_i_12_n_0 ),
        .I3(ir0[8]),
        .I4(crdy),
        .I5(ir0[6]),
        .O(\bdatw[15]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h5D5DFDFFFDFDFDFF)) 
    \bdatw[15]_INST_0_i_150 
       (.I0(\bdatw[15]_INST_0_i_228_n_0 ),
        .I1(\ccmd[4]_INST_0_i_17_n_0 ),
        .I2(ir0[8]),
        .I3(\ccmd[4]_INST_0_i_12_n_0 ),
        .I4(ir0[10]),
        .I5(\stat[0]_i_18_n_0 ),
        .O(\bdatw[15]_INST_0_i_150_n_0 ));
  LUT5 #(
    .INIT(32'h40040004)) 
    \bdatw[15]_INST_0_i_151 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .O(\bdatw[15]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'h10000000FFFFFFFF)) 
    \bdatw[15]_INST_0_i_152 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[5]),
        .I4(\ccmd[1]_INST_0_i_18_n_0 ),
        .I5(ir0[9]),
        .O(\bdatw[15]_INST_0_i_152_n_0 ));
  LUT6 #(
    .INIT(64'hAA222222A0222222)) 
    \bdatw[15]_INST_0_i_153 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .I2(\bdatw[15]_INST_0_i_229_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(\fadr[15]_INST_0_i_13_n_0 ),
        .O(\bdatw[15]_INST_0_i_153_n_0 ));
  LUT6 #(
    .INIT(64'h000000001D1DAA00)) 
    \bdatw[15]_INST_0_i_154 
       (.I0(ir0[7]),
        .I1(ir0[10]),
        .I2(crdy),
        .I3(ir0[6]),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\bdatw[15]_INST_0_i_154_n_0 ));
  LUT6 #(
    .INIT(64'h7000000000000070)) 
    \bdatw[15]_INST_0_i_155 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [2]),
        .I2(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I3(ir0[12]),
        .I4(ir0[11]),
        .I5(ir0[13]),
        .O(\bdatw[15]_INST_0_i_155_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF3E)) 
    \bdatw[15]_INST_0_i_156 
       (.I0(ir0[5]),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .I3(\bdatw[15]_INST_0_i_67_0 ),
        .I4(\bdatw[15]_INST_0_i_231_n_0 ),
        .O(\bdatw[15]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'h0000000008008908)) 
    \bdatw[15]_INST_0_i_157 
       (.I0(\stat_reg[0]_50 ),
        .I1(ir0[2]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ir0[3]),
        .I5(ir0[6]),
        .O(\bdatw[15]_INST_0_i_157_n_0 ));
  LUT4 #(
    .INIT(16'h00FD)) 
    \bdatw[15]_INST_0_i_158 
       (.I0(crdy),
        .I1(ir0[11]),
        .I2(\bdatw[15]_INST_0_i_232_n_0 ),
        .I3(\bdatw[15]_INST_0_i_167_n_0 ),
        .O(\bdatw[15]_INST_0_i_158_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \bdatw[15]_INST_0_i_159 
       (.I0(\bdatw[15]_INST_0_i_233_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[11]),
        .O(\bdatw[15]_INST_0_i_159_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAFBAAFBAAFBAA)) 
    \bdatw[15]_INST_0_i_160 
       (.I0(\bcmd[1] ),
        .I1(\bdatw[15]_INST_0_i_234_n_0 ),
        .I2(\bdatw[15]_INST_0_i_235_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I5(\badr[15]_INST_0_i_282_n_0 ),
        .O(\bdatw[15]_INST_0_i_160_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEFEEEAAAAAAAA)) 
    \bdatw[15]_INST_0_i_161 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\badr[15]_INST_0_i_201_n_0 ),
        .I2(ir0[2]),
        .I3(crdy),
        .I4(\bdatw[15]_INST_0_i_236_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .O(\bdatw[15]_INST_0_i_161_n_0 ));
  LUT6 #(
    .INIT(64'h8F88888800000000)) 
    \bdatw[15]_INST_0_i_162 
       (.I0(ir0[0]),
        .I1(\bdatw[15]_INST_0_i_237_n_0 ),
        .I2(\bdatw[15]_INST_0_i_238_n_0 ),
        .I3(ir0[9]),
        .I4(\ccmd[3]_INST_0_i_20_n_0 ),
        .I5(\stat[0]_i_7_n_0 ),
        .O(\bdatw[15]_INST_0_i_162_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFFAAAAAAAA)) 
    \bdatw[15]_INST_0_i_163 
       (.I0(\bcmd[1] ),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[0]),
        .I4(\bdatw[15]_INST_0_i_235_n_0 ),
        .I5(\bdatw[15]_INST_0_i_239_n_0 ),
        .O(\bdatw[15]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    \bdatw[15]_INST_0_i_164 
       (.I0(\bdatw[15]_INST_0_i_240_n_0 ),
        .I1(ir0[13]),
        .I2(\ccmd[3]_INST_0_i_18_n_0 ),
        .I3(\ccmd[2]_INST_0_i_3_0 ),
        .I4(ir0[15]),
        .I5(\ccmd[4]_INST_0_i_18_n_0 ),
        .O(\bdatw[15]_INST_0_i_164_n_0 ));
  LUT6 #(
    .INIT(64'h8A88888888888888)) 
    \bdatw[15]_INST_0_i_165 
       (.I0(\stat[0]_i_7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_237_n_0 ),
        .I2(\bdatw[15]_INST_0_i_241_n_0 ),
        .I3(ir0[9]),
        .I4(ir0[6]),
        .I5(\ccmd[3]_INST_0_i_20_n_0 ),
        .O(\bdatw[15]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'h15541555FFFFFFFF)) 
    \bdatw[15]_INST_0_i_166 
       (.I0(\bdatw[15]_INST_0_i_242_n_0 ),
        .I1(\bdatw[15]_INST_0_i_243_n_0 ),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(\ccmd[4]_INST_0_i_12_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .O(\bdatw[15]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFCC3FA0008000)) 
    \bdatw[15]_INST_0_i_167 
       (.I0(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(\bdatw[15]_INST_0_i_244_n_0 ),
        .O(\bdatw[15]_INST_0_i_167_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    \bdatw[15]_INST_0_i_168 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[12]),
        .I2(rst_n_fl_reg_2),
        .I3(ir0[2]),
        .I4(ir0[15]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\bdatw[15]_INST_0_i_168_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFDFDFFFDFF)) 
    \bdatw[15]_INST_0_i_169 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bcmd[1] ),
        .I2(\bdatw[15]_INST_0_i_245_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\bdatw[15]_INST_0_i_246_n_0 ),
        .I5(\bcmd[0]_INST_0_i_9_n_0 ),
        .O(\stat_reg[0]_46 ));
  LUT6 #(
    .INIT(64'hA2A2A280FFFFFFFF)) 
    \bdatw[15]_INST_0_i_17 
       (.I0(\bdatw[15]_INST_0_i_57_n_0 ),
        .I1(ir0[15]),
        .I2(\bcmd[0]_INST_0_i_9_n_0 ),
        .I3(\bdatw[15]_INST_0_i_58_n_0 ),
        .I4(\bdatw[15]_INST_0_i_59_n_0 ),
        .I5(ctl_fetch0_fl_reg_0),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDFDDDF)) 
    \bdatw[15]_INST_0_i_170 
       (.I0(\stat_reg[2]_17 ),
        .I1(\bdatw[15]_INST_0_i_163_n_0 ),
        .I2(\bdatw[15]_INST_0_i_172_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I4(\bdatw[15]_INST_0_i_247_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\stat_reg[0]_23 ));
  LUT6 #(
    .INIT(64'h8088AAAA80888088)) 
    \bdatw[15]_INST_0_i_171 
       (.I0(\bcmd[0]_INST_0_i_9_n_0 ),
        .I1(ir0[1]),
        .I2(\bdatw[15]_INST_0_i_167_n_0 ),
        .I3(\bdatw[15]_INST_0_i_166_n_0 ),
        .I4(\bdatw[15]_INST_0_i_233_n_0 ),
        .I5(\stat[0]_i_7_n_0 ),
        .O(\bdatw[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA8A888888888)) 
    \bdatw[15]_INST_0_i_172 
       (.I0(\bcmd[0]_INST_0_i_9_n_0 ),
        .I1(\bdatw[15]_INST_0_i_162_n_0 ),
        .I2(\bdatw[15]_INST_0_i_167_n_0 ),
        .I3(\bdatw[15]_INST_0_i_232_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I5(ir0[0]),
        .O(\bdatw[15]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA200020002000)) 
    \bdatw[15]_INST_0_i_173 
       (.I0(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I1(\bdatw[15]_INST_0_i_236_n_0 ),
        .I2(crdy),
        .I3(ir0[2]),
        .I4(fch_irq_req),
        .I5(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .O(\bdatw[15]_INST_0_i_173_n_0 ));
  LUT6 #(
    .INIT(64'h10111010FFFFFFFF)) 
    \bdatw[15]_INST_0_i_174 
       (.I0(\bcmd[1] ),
        .I1(\bdatw[15]_INST_0_i_245_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\bdatw[15]_INST_0_i_246_n_0 ),
        .I4(\bcmd[0]_INST_0_i_9_n_0 ),
        .I5(\stat_reg[2]_17 ),
        .O(\stat_reg[0]_21 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40C40010)) 
    \bdatw[15]_INST_0_i_177 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(\read_cyc_reg[1] ),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_177_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF7776)) 
    \bdatw[15]_INST_0_i_178 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .I4(\bdatw[15]_INST_0_i_248_n_0 ),
        .O(\bdatw[15]_INST_0_i_178_n_0 ));
  LUT6 #(
    .INIT(64'h7F77FFFF7F77BFBB)) 
    \bdatw[15]_INST_0_i_179 
       (.I0(ir1[11]),
        .I1(\bdatw[15]_INST_0_i_197_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(ir1[10]),
        .I5(ir1[5]),
        .O(\bdatw[15]_INST_0_i_179_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEAEEEAAAA)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_60_n_0 ),
        .I1(ir0[12]),
        .I2(\bdatw[15]_INST_0_i_61_n_0 ),
        .I3(\bdatw[15]_INST_0_i_62_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\bdatw[15]_INST_0_i_63_n_0 ),
        .O(\stat_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h1F001F0055000000)) 
    \bdatw[15]_INST_0_i_180 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .I2(\bdatw[15]_INST_0_i_249_n_0 ),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(ir1[10]),
        .O(\bdatw[15]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'h00001C10FFFFFFFF)) 
    \bdatw[15]_INST_0_i_181 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(ir1[11]),
        .O(\bdatw[15]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'hA2A2020082820200)) 
    \bdatw[15]_INST_0_i_182 
       (.I0(\bdatw[15]_INST_0_i_250_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(rst_n_fl_reg_9),
        .I4(ir1[10]),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_182_n_0 ));
  LUT6 #(
    .INIT(64'h44C444C444C44444)) 
    \bdatw[15]_INST_0_i_183 
       (.I0(\bdatw[15]_INST_0_i_251_n_0 ),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .I3(\stat[1]_i_18_n_0 ),
        .I4(\bdatw[15]_INST_0_i_252_n_0 ),
        .I5(rst_n_fl_reg_9),
        .O(\bdatw[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'h0000A959FFFFFFFF)) 
    \bdatw[15]_INST_0_i_184 
       (.I0(ir1[11]),
        .I1(\sr_reg[15]_0 [4]),
        .I2(ir1[14]),
        .I3(\bbus_o[4]_INST_0_i_49_0 ),
        .I4(ir1[13]),
        .I5(ir1[12]),
        .O(\bdatw[15]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF3B04FFFF0B34)) 
    \bdatw[15]_INST_0_i_185 
       (.I0(\sr_reg[15]_0 [5]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[12]),
        .I5(\sr_reg[15]_0 [6]),
        .O(\bdatw[15]_INST_0_i_185_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[15]_INST_0_i_186 
       (.I0(ir1[14]),
        .I1(ir1[11]),
        .O(\bdatw[15]_INST_0_i_186_n_0 ));
  LUT4 #(
    .INIT(16'h0F2F)) 
    \bdatw[15]_INST_0_i_187 
       (.I0(\sr_reg[15]_0 [6]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .O(\bdatw[15]_INST_0_i_187_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[15]_INST_0_i_188 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .O(\bdatw[15]_INST_0_i_188_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_189 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .O(\bdatw[15]_INST_0_i_189_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_19 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .O(\bdatw[15]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h00011011)) 
    \bdatw[15]_INST_0_i_190 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .O(\bdatw[15]_INST_0_i_190_n_0 ));
  LUT5 #(
    .INIT(32'hFF46FFFF)) 
    \bdatw[15]_INST_0_i_191 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .I3(ir1[11]),
        .I4(ir1[6]),
        .O(\bdatw[15]_INST_0_i_191_n_0 ));
  LUT5 #(
    .INIT(32'h2F2C3D3F)) 
    \bdatw[15]_INST_0_i_192 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(ir1[8]),
        .O(\bdatw[15]_INST_0_i_192_n_0 ));
  LUT4 #(
    .INIT(16'h0041)) 
    \bdatw[15]_INST_0_i_193 
       (.I0(ir1[3]),
        .I1(ir1[6]),
        .I2(ir1[4]),
        .I3(ir1[5]),
        .O(\bdatw[15]_INST_0_i_193_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \bdatw[15]_INST_0_i_194 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\bdatw[15]_INST_0_i_194_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \bdatw[15]_INST_0_i_195 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .O(\bdatw[15]_INST_0_i_195_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \bdatw[15]_INST_0_i_196 
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .I2(ir1[3]),
        .I3(ir1[6]),
        .O(\bdatw[15]_INST_0_i_196_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[15]_INST_0_i_197 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\bdatw[15]_INST_0_i_197_n_0 ));
  LUT5 #(
    .INIT(32'h3F030200)) 
    \bdatw[15]_INST_0_i_198 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[3]),
        .I2(ir1[1]),
        .I3(ir1[0]),
        .I4(ir1[2]),
        .O(\bdatw[15]_INST_0_i_198_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bdatw[15]_INST_0_i_199 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(ir1[14]),
        .O(\bdatw[15]_INST_0_i_199_n_0 ));
  LUT5 #(
    .INIT(32'h000000A2)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(\bdatw[15]_INST_0_i_12_n_0 ),
        .I1(eir[15]),
        .I2(\bdatw[15]_INST_0_i_13_n_0 ),
        .I3(\bdatw[15]_1 ),
        .I4(\bdatw[15]_2 ),
        .O(fch_leir_nir_reg));
  LUT6 #(
    .INIT(64'h0000000000005DDD)) 
    \bdatw[15]_INST_0_i_202 
       (.I0(ir1[1]),
        .I1(\bdatw[15]_INST_0_i_253_n_0 ),
        .I2(ir1[10]),
        .I3(\bdatw[15]_INST_0_i_254_n_0 ),
        .I4(\bdatw[15]_INST_0_i_255_n_0 ),
        .I5(\bdatw[15]_INST_0_i_208_n_0 ),
        .O(\bdatw[15]_INST_0_i_202_n_0 ));
  LUT6 #(
    .INIT(64'h0000F7FFF7FFF7FF)) 
    \bdatw[15]_INST_0_i_203 
       (.I0(\bdatw[15]_INST_0_i_256_n_0 ),
        .I1(ir1[1]),
        .I2(\bdatw[15]_INST_0_i_257_n_0 ),
        .I3(ir1[14]),
        .I4(\badr[15]_INST_0_i_70_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .O(\bdatw[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \bdatw[15]_INST_0_i_204 
       (.I0(\bdatw[15]_INST_0_i_256_n_0 ),
        .I1(ir1[14]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[0]),
        .O(\bdatw[15]_INST_0_i_204_n_0 ));
  LUT6 #(
    .INIT(64'h0000D5DDD5DDD5DD)) 
    \bdatw[15]_INST_0_i_205 
       (.I0(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I1(\bdatw[15]_INST_0_i_258_n_0 ),
        .I2(\bdatw[15]_INST_0_i_207_n_0 ),
        .I3(ir1[0]),
        .I4(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I5(\badr[15]_INST_0_i_160_n_0 ),
        .O(\bdatw[15]_INST_0_i_205_n_0 ));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \bdatw[15]_INST_0_i_206 
       (.I0(\bdatw[15]_INST_0_i_259_n_0 ),
        .I1(\badr[15]_INST_0_i_90_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(\bdatw[15]_INST_0_i_260_n_0 ),
        .O(\bdatw[15]_INST_0_i_206_n_0 ));
  LUT6 #(
    .INIT(64'h0000000044454545)) 
    \bdatw[15]_INST_0_i_207 
       (.I0(\bdatw[15]_INST_0_i_261_n_0 ),
        .I1(ir1[11]),
        .I2(\bdatw[15]_INST_0_i_262_n_0 ),
        .I3(rst_n_fl_reg_9),
        .I4(\bdatw[15]_INST_0_i_263_n_0 ),
        .I5(\bdatw[15]_INST_0_i_264_n_0 ),
        .O(\bdatw[15]_INST_0_i_207_n_0 ));
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \bdatw[15]_INST_0_i_208 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(ir1[6]),
        .O(\bdatw[15]_INST_0_i_208_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_209 
       (.I0(ir1[2]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .O(\bdatw[15]_INST_0_i_209_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF888A)) 
    \bdatw[15]_INST_0_i_21 
       (.I0(\bdatw[15]_INST_0_i_64_n_0 ),
        .I1(\bdatw[15]_INST_0_i_65_n_0 ),
        .I2(rst_n_fl_reg_2),
        .I3(\bdatw[15]_INST_0_i_66_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\bdatw[15]_INST_0_i_67_n_0 ),
        .O(ctl_selb0_0));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_22 
       (.I0(ctl_selb0_rn[1]),
        .I1(ctl_selb0_rn[0]),
        .I2(\stat_reg[2]_17 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .O(b0bus_sel_cr[3]));
  LUT6 #(
    .INIT(64'h2B002B002B000000)) 
    \bdatw[15]_INST_0_i_222 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .I4(crdy),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\bdatw[15]_INST_0_i_222_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_223 
       (.I0(ir0[8]),
        .I1(crdy),
        .O(\bdatw[15]_INST_0_i_223_n_0 ));
  LUT4 #(
    .INIT(16'h2023)) 
    \bdatw[15]_INST_0_i_224 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .O(\bdatw[15]_INST_0_i_224_n_0 ));
  LUT5 #(
    .INIT(32'h00BB00C3)) 
    \bdatw[15]_INST_0_i_225 
       (.I0(crdy),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[9]),
        .I4(ir0[10]),
        .O(\bdatw[15]_INST_0_i_225_n_0 ));
  LUT3 #(
    .INIT(8'h1A)) 
    \bdatw[15]_INST_0_i_226 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .O(\bdatw[15]_INST_0_i_226_n_0 ));
  LUT4 #(
    .INIT(16'h2A02)) 
    \bdatw[15]_INST_0_i_227 
       (.I0(crdy),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .O(\bdatw[15]_INST_0_i_227_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_228 
       (.I0(ir0[6]),
        .I1(ir0[11]),
        .O(\bdatw[15]_INST_0_i_228_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[15]_INST_0_i_229 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(ir0[5]),
        .O(\bdatw[15]_INST_0_i_229_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_23 
       (.I0(ctl_selb0_rn[1]),
        .I1(ctl_selb0_rn[0]),
        .I2(\stat_reg[2]_17 ),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .O(b0bus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h3FFA)) 
    \bdatw[15]_INST_0_i_231 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .O(\bdatw[15]_INST_0_i_231_n_0 ));
  LUT6 #(
    .INIT(64'h3FFD0DCD3FFDCDCD)) 
    \bdatw[15]_INST_0_i_232 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[6]),
        .I4(ir0[9]),
        .I5(ir0[7]),
        .O(\bdatw[15]_INST_0_i_232_n_0 ));
  LUT6 #(
    .INIT(64'hAF30FFF0FF30FFFF)) 
    \bdatw[15]_INST_0_i_233 
       (.I0(\bdatw[15]_INST_0_i_241_n_0 ),
        .I1(crdy),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(ir0[1]),
        .I5(\rgf_selc0_rn_wb[1]_i_27_n_0 ),
        .O(\bdatw[15]_INST_0_i_233_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bdatw[15]_INST_0_i_234 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[1]),
        .O(\bdatw[15]_INST_0_i_234_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_235 
       (.I0(ir0[11]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(ir0[10]),
        .I5(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .O(\bdatw[15]_INST_0_i_235_n_0 ));
  LUT3 #(
    .INIT(8'hD4)) 
    \bdatw[15]_INST_0_i_236 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[3]),
        .O(\bdatw[15]_INST_0_i_236_n_0 ));
  LUT5 #(
    .INIT(32'h40454545)) 
    \bdatw[15]_INST_0_i_237 
       (.I0(ir0[9]),
        .I1(crdy),
        .I2(ir0[8]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .O(\bdatw[15]_INST_0_i_237_n_0 ));
  LUT5 #(
    .INIT(32'hC6FBFFFB)) 
    \bdatw[15]_INST_0_i_238 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .I4(ir0[0]),
        .O(\bdatw[15]_INST_0_i_238_n_0 ));
  LUT6 #(
    .INIT(64'h2AAAAAAAAAAAAAAA)) 
    \bdatw[15]_INST_0_i_239 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .I4(\ccmd[4]_INST_0_i_15_n_0 ),
        .I5(\badr[15]_INST_0_i_282_n_0 ),
        .O(\bdatw[15]_INST_0_i_239_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \bdatw[15]_INST_0_i_240 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(ir0[2]),
        .I3(ir0[6]),
        .O(\bdatw[15]_INST_0_i_240_n_0 ));
  LUT3 #(
    .INIT(8'hC6)) 
    \bdatw[15]_INST_0_i_241 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(ir0[5]),
        .O(\bdatw[15]_INST_0_i_241_n_0 ));
  LUT5 #(
    .INIT(32'h0000D500)) 
    \bdatw[15]_INST_0_i_242 
       (.I0(ir0[8]),
        .I1(ir0[6]),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(ir0[9]),
        .O(\bdatw[15]_INST_0_i_242_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_243 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .O(\bdatw[15]_INST_0_i_243_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_244 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\bdatw[15]_INST_0_i_244_n_0 ));
  LUT6 #(
    .INIT(64'h7000707070707070)) 
    \bdatw[15]_INST_0_i_245 
       (.I0(\badr[15]_INST_0_i_282_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\bdatw[15]_INST_0_i_235_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_27_n_0 ),
        .I5(ir0[1]),
        .O(\bdatw[15]_INST_0_i_245_n_0 ));
  LUT6 #(
    .INIT(64'h0000DD0DDDDDDDDD)) 
    \bdatw[15]_INST_0_i_246 
       (.I0(\stat[0]_i_7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_233_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I3(\bdatw[15]_INST_0_i_232_n_0 ),
        .I4(\bdatw[15]_INST_0_i_167_n_0 ),
        .I5(ir0[1]),
        .O(\bdatw[15]_INST_0_i_246_n_0 ));
  LUT6 #(
    .INIT(64'hFF3F3F1DFFFFFF3F)) 
    \bdatw[15]_INST_0_i_247 
       (.I0(fch_irq_req),
        .I1(ir0[2]),
        .I2(crdy),
        .I3(ir0[3]),
        .I4(ir0[1]),
        .I5(ir0[0]),
        .O(\bdatw[15]_INST_0_i_247_n_0 ));
  LUT4 #(
    .INIT(16'hFEE6)) 
    \bdatw[15]_INST_0_i_248 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\rgf_selc1_wb_reg[1] [2]),
        .O(\bdatw[15]_INST_0_i_248_n_0 ));
  LUT6 #(
    .INIT(64'h1D33000000000000)) 
    \bdatw[15]_INST_0_i_249 
       (.I0(ir1[6]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[8]),
        .I5(ir1[7]),
        .O(\bdatw[15]_INST_0_i_249_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_250 
       (.I0(ir1[6]),
        .I1(ir1[11]),
        .O(\bdatw[15]_INST_0_i_250_n_0 ));
  LUT3 #(
    .INIT(8'hDE)) 
    \bdatw[15]_INST_0_i_251 
       (.I0(\sr_reg[15]_0 [7]),
        .I1(ir1[14]),
        .I2(ir1[11]),
        .O(\bdatw[15]_INST_0_i_251_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_252 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\bdatw[15]_INST_0_i_252_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00DF)) 
    \bdatw[15]_INST_0_i_253 
       (.I0(\badr[15]_INST_0_i_244_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_14_n_0 ),
        .I2(rst_n_fl_reg_9),
        .I3(\bdatw[15]_INST_0_i_262_n_0 ),
        .I4(ir1[11]),
        .I5(\bdatw[15]_INST_0_i_261_n_0 ),
        .O(\bdatw[15]_INST_0_i_253_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_254 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .O(\bdatw[15]_INST_0_i_254_n_0 ));
  LUT6 #(
    .INIT(64'h3900000000000000)) 
    \bdatw[15]_INST_0_i_255 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .I2(ir1[5]),
        .I3(\badr[15]_INST_0_i_243_n_0 ),
        .I4(ir1[6]),
        .I5(ir1[1]),
        .O(\bdatw[15]_INST_0_i_255_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \bdatw[15]_INST_0_i_256 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .I2(ir1[13]),
        .I3(ir1[10]),
        .I4(ir1[8]),
        .I5(ir1[9]),
        .O(\bdatw[15]_INST_0_i_256_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[15]_INST_0_i_257 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .O(\bdatw[15]_INST_0_i_257_n_0 ));
  LUT6 #(
    .INIT(64'hDDFF7DF7FFFFFFF7)) 
    \bdatw[15]_INST_0_i_258 
       (.I0(\badr[15]_INST_0_i_243_n_0 ),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .I4(ir1[5]),
        .I5(ir1[0]),
        .O(\bdatw[15]_INST_0_i_258_n_0 ));
  LUT3 #(
    .INIT(8'h63)) 
    \bdatw[15]_INST_0_i_259 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .I2(ir1[4]),
        .O(\bdatw[15]_INST_0_i_259_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \bdatw[15]_INST_0_i_260 
       (.I0(ir1[9]),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[2]),
        .O(\bdatw[15]_INST_0_i_260_n_0 ));
  LUT6 #(
    .INIT(64'h00DD000000B50000)) 
    \bdatw[15]_INST_0_i_261 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .I5(ir1[9]),
        .O(\bdatw[15]_INST_0_i_261_n_0 ));
  LUT5 #(
    .INIT(32'hC80F0000)) 
    \bdatw[15]_INST_0_i_262 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[10]),
        .O(\bdatw[15]_INST_0_i_262_n_0 ));
  LUT4 #(
    .INIT(16'h0111)) 
    \bdatw[15]_INST_0_i_263 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .O(\bdatw[15]_INST_0_i_263_n_0 ));
  LUT6 #(
    .INIT(64'h0808080800080808)) 
    \bdatw[15]_INST_0_i_264 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(ir1[8]),
        .O(\bdatw[15]_INST_0_i_264_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(\stat_reg[2]_5 ),
        .I1(\stat_reg[1]_5 [1]),
        .O(\bcmd[2]_INST_0_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[15]_INST_0_i_37 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [15]),
        .O(b0bus_sr[15]));
  LUT6 #(
    .INIT(64'hDDDDDDDDCFFFFFFF)) 
    \bdatw[15]_INST_0_i_38 
       (.I0(\bdatw[15]_INST_0_i_99_n_0 ),
        .I1(ir1[15]),
        .I2(\bdatw[15]_INST_0_i_100_n_0 ),
        .I3(\bdatw[15]_INST_0_i_101_n_0 ),
        .I4(\read_cyc_reg[1] ),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\stat_reg[0]_12 ));
  LUT6 #(
    .INIT(64'h22A222A222A2AAAA)) 
    \bdatw[15]_INST_0_i_39 
       (.I0(\stat[0]_i_2__1_0 ),
        .I1(\bdatw[15]_INST_0_i_103_n_0 ),
        .I2(ir1[15]),
        .I3(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I4(\bdatw[15]_INST_0_i_104_n_0 ),
        .I5(\bdatw[15]_INST_0_i_105_n_0 ),
        .O(\stat_reg[0]_11 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \bdatw[15]_INST_0_i_40 
       (.I0(ctl_selb1_0),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .O(\bdatw[15]_INST_0_i_40_n_0 ));
  LUT3 #(
    .INIT(8'h54)) 
    \bdatw[15]_INST_0_i_41 
       (.I0(\stat_reg[0]_12 ),
        .I1(ctl_selb1_0),
        .I2(ir1[10]),
        .O(\bdatw[15]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0E00FF000E000000)) 
    \bdatw[15]_INST_0_i_42 
       (.I0(\bdatw[15]_INST_0_i_106_n_0 ),
        .I1(\bdatw[15]_INST_0_i_107_n_0 ),
        .I2(\bdatw[15]_INST_0_i_108_n_0 ),
        .I3(\bcmd[1]_0 ),
        .I4(ir1[12]),
        .I5(\bdatw[15]_INST_0_i_109_n_0 ),
        .O(ctl_selb1_0));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_45 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .O(b1bus_sel_cr[3]));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_46 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .O(b1bus_sel_cr[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_5 
       (.I0(\stat_reg[1]_5 [1]),
        .I1(\stat_reg[2]_5 ),
        .O(\bcmd[1]_INST_0_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bdatw[15]_INST_0_i_50 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .O(b1bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'hAA0A08A8A00008A8)) 
    \bdatw[15]_INST_0_i_51 
       (.I0(\stat_reg[0]_11 ),
        .I1(ir1[6]),
        .I2(ctl_selb1_0),
        .I3(\bdatw[15]_INST_0_i_129_n_0 ),
        .I4(\stat_reg[0]_12 ),
        .I5(ir1[7]),
        .O(rst_n_fl_reg_12));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_52 
       (.I0(eir[7]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_5));
  LUT6 #(
    .INIT(64'h55757757FFFFFFFF)) 
    \bdatw[15]_INST_0_i_57 
       (.I0(\bdatw[15]_INST_0_i_59_n_0 ),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(\sr_reg[15]_0 [5]),
        .I4(ir0[11]),
        .I5(\rgf_selc0_wb[1]_i_4_1 ),
        .O(\bdatw[15]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h1EFCDEFC)) 
    \bdatw[15]_INST_0_i_58 
       (.I0(\sr_reg[15]_0 [7]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(\bdatw[15]_INST_0_i_140_n_0 ),
        .O(\bdatw[15]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'h02FF)) 
    \bdatw[15]_INST_0_i_59 
       (.I0(\sr_reg[15]_0 [6]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[13]),
        .O(\bdatw[15]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hBAAAEFFFFEEEEFFF)) 
    \bdatw[15]_INST_0_i_6 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(fctl_n_133),
        .I4(ctl_selb0_0),
        .I5(ir0[10]),
        .O(\stat_reg[0]_24 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFBFFFF)) 
    \bdatw[15]_INST_0_i_60 
       (.I0(\bcmd[1] ),
        .I1(\bdatw[15]_INST_0_i_141_n_0 ),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .I4(\ccmd[0]_INST_0_i_23_n_0 ),
        .I5(ir0[12]),
        .O(\bdatw[15]_INST_0_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[15]_INST_0_i_61 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\bdatw[15]_INST_0_i_61_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[15]_INST_0_i_62 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[8]),
        .O(\bdatw[15]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hAABABBBBAABAAAAA)) 
    \bdatw[15]_INST_0_i_63 
       (.I0(rst_n_fl_reg_2),
        .I1(\bdatw[15]_INST_0_i_142_n_0 ),
        .I2(\bdatw[15]_INST_0_i_143_n_0 ),
        .I3(\bdatw[15]_INST_0_i_144_n_0 ),
        .I4(ir0[11]),
        .I5(\bdatw[15]_INST_0_i_145_n_0 ),
        .O(\bdatw[15]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h1010101010101011)) 
    \bdatw[15]_INST_0_i_64 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(\bdatw[15]_INST_0_i_146_n_0 ),
        .I3(\bdatw[15]_INST_0_i_147_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[14]),
        .O(\bdatw[15]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'hDFFFDCDC)) 
    \bdatw[15]_INST_0_i_65 
       (.I0(\bdatw[15]_INST_0_i_148_n_0 ),
        .I1(\bdatw[15]_INST_0_i_149_n_0 ),
        .I2(ir0[13]),
        .I3(ir0[12]),
        .I4(\rgf_selc0_wb[1]_i_4_1 ),
        .O(\bdatw[15]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h2222222200022222)) 
    \bdatw[15]_INST_0_i_66 
       (.I0(\bdatw[15]_INST_0_i_150_n_0 ),
        .I1(\bdatw[15]_INST_0_i_151_n_0 ),
        .I2(\bdatw[15]_INST_0_i_152_n_0 ),
        .I3(\bdatw[15]_INST_0_i_153_n_0 ),
        .I4(ir0[11]),
        .I5(\bdatw[15]_INST_0_i_154_n_0 ),
        .O(\bdatw[15]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFDD00DF00)) 
    \bdatw[15]_INST_0_i_67 
       (.I0(\bdatw[15]_INST_0_i_155_n_0 ),
        .I1(\bdatw[15]_INST_0_i_156_n_0 ),
        .I2(ir0[7]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\bdatw[15]_INST_0_i_157_n_0 ),
        .I5(ir0[15]),
        .O(\bdatw[15]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF08AA)) 
    \bdatw[15]_INST_0_i_68 
       (.I0(\bcmd[0]_INST_0_i_9_n_0 ),
        .I1(ir0[1]),
        .I2(\bdatw[15]_INST_0_i_158_n_0 ),
        .I3(\bdatw[15]_INST_0_i_159_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\bdatw[15]_INST_0_i_160_n_0 ),
        .O(ctl_selb0_rn[1]));
  LUT6 #(
    .INIT(64'h00000000EAEEEAEA)) 
    \bdatw[15]_INST_0_i_69 
       (.I0(\bdatw[15]_INST_0_i_161_n_0 ),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .I2(\bdatw[15]_INST_0_i_162_n_0 ),
        .I3(\bdatw[15]_INST_0_i_158_n_0 ),
        .I4(ir0[0]),
        .I5(\bdatw[15]_INST_0_i_163_n_0 ),
        .O(ctl_selb0_rn[0]));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[15]),
        .O(\stat_reg[0]_44 ));
  LUT6 #(
    .INIT(64'h4444444455555455)) 
    \bdatw[15]_INST_0_i_70 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\bdatw[15]_INST_0_i_164_n_0 ),
        .I2(\bdatw[15]_INST_0_i_165_n_0 ),
        .I3(\bdatw[15]_INST_0_i_166_n_0 ),
        .I4(\bdatw[15]_INST_0_i_167_n_0 ),
        .I5(\bdatw[15]_INST_0_i_168_n_0 ),
        .O(\stat_reg[2]_17 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \bdatw[15]_INST_0_i_71 
       (.I0(ctl_selb0_0),
        .I1(\stat_reg[0]_7 ),
        .I2(\sr_reg[5] ),
        .O(\bdatw[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F5F5F4F4F4F44)) 
    \bdatw[15]_INST_0_i_75 
       (.I0(\bdatw[15]_INST_0_i_160_n_0 ),
        .I1(\bdatw[15]_INST_0_i_171_n_0 ),
        .I2(\bdatw[15]_INST_0_i_163_n_0 ),
        .I3(\bdatw[15]_INST_0_i_172_n_0 ),
        .I4(\bdatw[15]_INST_0_i_173_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\stat_reg[0]_45 ));
  LUT6 #(
    .INIT(64'hFAFAFAFAFBFBFBFF)) 
    \bdatw[15]_INST_0_i_76 
       (.I0(\bdatw[15]_INST_0_i_160_n_0 ),
        .I1(\bdatw[15]_INST_0_i_171_n_0 ),
        .I2(\bdatw[15]_INST_0_i_163_n_0 ),
        .I3(\bdatw[15]_INST_0_i_172_n_0 ),
        .I4(\bdatw[15]_INST_0_i_173_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\stat_reg[0]_22 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \bdatw[15]_INST_0_i_84 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[5] ),
        .I4(\stat_reg[0]_7 ),
        .I5(ctl_selb0_0),
        .O(b0bus_sel_cr[4]));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \bdatw[15]_INST_0_i_85 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\sr_reg[5] ),
        .I4(\stat_reg[0]_7 ),
        .I5(ctl_selb0_0),
        .O(b0bus_sel_cr[1]));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \bdatw[15]_INST_0_i_86 
       (.I0(ctl_selb0_rn[1]),
        .I1(\stat_reg[2]_17 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\sr_reg[5] ),
        .I4(\stat_reg[0]_7 ),
        .I5(ctl_selb0_0),
        .O(b0bus_sel_cr[0]));
  LUT6 #(
    .INIT(64'h0000000000008002)) 
    \bdatw[15]_INST_0_i_99 
       (.I0(\bdatw[15]_INST_0_i_177_n_0 ),
        .I1(ir1[13]),
        .I2(ir1[11]),
        .I3(ir1[12]),
        .I4(\bdatw[15]_INST_0_i_178_n_0 ),
        .I5(\bdatw[15]_INST_0_i_179_n_0 ),
        .O(\bdatw[15]_INST_0_i_99_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[1]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[9]_INST_0_i_3_n_0 ),
        .O(bdatw[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[2]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[10]_INST_0_i_3_n_0 ),
        .O(bdatw[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[3]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[11]_INST_0_i_3_n_0 ),
        .O(bdatw[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[4]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[12]_INST_0_i_3_n_0 ),
        .O(bdatw[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[5]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bdatw_5_sn_1),
        .O(bdatw[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[6]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(bdatw_6_sn_1),
        .O(bdatw[6]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[7]_INST_0 
       (.I0(\stat_reg[2]_5 ),
        .I1(\bdatw[15]_0 ),
        .O(bdatw[7]));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[8]_INST_0 
       (.I0(\bdatw[8]_0 ),
        .I1(\stat_reg[0]_48 ),
        .I2(bdatw_8_sn_1),
        .I3(\bcmd[2]_INST_0_0 ),
        .I4(\bdatw[8]_INST_0_i_3_n_0 ),
        .I5(\bcmd[1]_INST_0_0 ),
        .O(bdatw[8]));
  LUT5 #(
    .INIT(32'h82828280)) 
    \bdatw[8]_INST_0_i_10 
       (.I0(\stat_reg[0]_11 ),
        .I1(\stat_reg[0]_12 ),
        .I2(\bdatw[8]_INST_0_i_28_n_0 ),
        .I3(ir1[7]),
        .I4(ctl_selb1_0),
        .O(\stat_reg[0]_33 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_11 
       (.I0(eir[8]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_4));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[8]_INST_0_i_16 
       (.I0(\bdatw[8]_INST_0_i_39_n_0 ),
        .I1(\bdatw[8]_INST_0_i_40_n_0 ),
        .I2(\sr[6]_i_16 ),
        .I3(b1bus_b02[0]),
        .I4(\sr[6]_i_16_0 ),
        .I5(\sr[6]_i_16_1 ),
        .O(\tr_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    \bdatw[8]_INST_0_i_17 
       (.I0(ir0[0]),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .I3(ir0[3]),
        .I4(\stat_reg[0]_7 ),
        .O(\bdatw[8]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[8]_INST_0_i_27 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [8]),
        .O(b0bus_sr[8]));
  LUT5 #(
    .INIT(32'h00000200)) 
    \bdatw[8]_INST_0_i_28 
       (.I0(ctl_selb1_0),
        .I1(ir1[1]),
        .I2(ir1[2]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .O(\bdatw[8]_INST_0_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(\tr_reg[0]_0 ),
        .I1(\stat_reg[0]_48 ),
        .I2(\tr_reg[0] ),
        .O(\bdatw[8]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[8]_INST_0_i_38 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [8]),
        .O(b1bus_sr[8]));
  LUT6 #(
    .INIT(64'hAAA655FFFFFFFFFF)) 
    \bdatw[8]_INST_0_i_39 
       (.I0(\stat_reg[0]_12 ),
        .I1(\bdatw[8]_INST_0_i_57_n_0 ),
        .I2(ir1[2]),
        .I3(ir1[0]),
        .I4(ctl_selb1_0),
        .I5(\stat_reg[0]_11 ),
        .O(\bdatw[8]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hBEFEBEBE)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[8]_INST_0_i_17_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ir0[7]),
        .I4(\stat_reg[0]_7 ),
        .O(\stat_reg[0]_9 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_40 
       (.I0(eir[0]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(\bdatw[8]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[8]_INST_0_i_5 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[8]),
        .O(\stat_reg[0]_37 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[8]_INST_0_i_57 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .O(\bdatw[8]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[8]_INST_0_i_64 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_117_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_0 [0]),
        .O(b1bus_sr[0]));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bdatw[8]_INST_0_i_72 
       (.I0(\stat_reg[0]_19 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [0]),
        .O(\sr_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bdatw[8]_INST_0_i_73 
       (.I0(\stat_reg[0]_20 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_64 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[9]_INST_0 
       (.I0(bdatw_9_sn_1),
        .I1(\stat_reg[0]_48 ),
        .I2(\bdatw[9]_0 ),
        .I3(\bcmd[2]_INST_0_0 ),
        .I4(\bdatw[9]_INST_0_i_3_n_0 ),
        .I5(\bcmd[1]_INST_0_0 ),
        .O(bdatw[9]));
  LUT6 #(
    .INIT(64'h8280222022202220)) 
    \bdatw[9]_INST_0_i_10 
       (.I0(\stat_reg[0]_11 ),
        .I1(\stat_reg[0]_12 ),
        .I2(ctl_selb1_0),
        .I3(ir1[8]),
        .I4(\bdatw[11]_INST_0_i_28_n_0 ),
        .I5(fctl_n_95),
        .O(\stat_reg[0]_14 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[9]_INST_0_i_11 
       (.I0(eir[9]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(fch_leir_nir_reg_3));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \bdatw[9]_INST_0_i_16 
       (.I0(\bdatw[9]_INST_0_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_28_0 ),
        .I2(b1bus_b02[1]),
        .I3(\rgf_c1bus_wb[14]_i_28_1 ),
        .I4(\rgf_c1bus_wb[14]_i_28_2 ),
        .I5(\bdatw[9]_INST_0_i_44_n_0 ),
        .O(\bdatw[9]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[9]_INST_0_i_17 
       (.I0(ir0[1]),
        .I1(ir0[0]),
        .I2(ir0[3]),
        .I3(ir0[2]),
        .O(\bdatw[9]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[9]_INST_0_i_27 
       (.I0(\stat_reg[2]_17 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_71_n_0 ),
        .I4(\sr_reg[15]_0 [9]),
        .O(b0bus_sr[9]));
  LUT3 #(
    .INIT(8'h8B)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_48 ),
        .I2(\bdatw[9]_INST_0_i_16_n_0 ),
        .O(\bdatw[9]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[9]_INST_0_i_38 
       (.I0(b1bus_sel_cr[0]),
        .I1(\sr_reg[15]_0 [9]),
        .O(b1bus_sr[9]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[9]_INST_0_i_39 
       (.I0(eir[1]),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .O(\bdatw[9]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hAEFBFEFB)) 
    \bdatw[9]_INST_0_i_4 
       (.I0(\sr_reg[5] ),
        .I1(\bdatw[9]_INST_0_i_17_n_0 ),
        .I2(\stat_reg[0]_7 ),
        .I3(ctl_selb0_0),
        .I4(ir0[8]),
        .O(\stat_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \bdatw[9]_INST_0_i_44 
       (.I0(ir1[0]),
        .I1(ctl_selb1_0),
        .I2(\bdatw[9]_INST_0_i_69_n_0 ),
        .I3(\stat_reg[0]_12 ),
        .I4(ir1[1]),
        .I5(\stat_reg[0]_11 ),
        .O(\bdatw[9]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \bdatw[9]_INST_0_i_5 
       (.I0(\sr_reg[5] ),
        .I1(\stat_reg[0]_7 ),
        .I2(ctl_selb0_0),
        .I3(eir[9]),
        .O(\stat_reg[0]_38 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[9]_INST_0_i_63 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_117_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\sr_reg[15]_0 [1]),
        .O(b1bus_sr[1]));
  LUT4 #(
    .INIT(16'h0004)) 
    \bdatw[9]_INST_0_i_69 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(ir1[2]),
        .I3(ir1[3]),
        .O(\bdatw[9]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bdatw[9]_INST_0_i_72 
       (.I0(\stat_reg[0]_19 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [1]),
        .O(\sr_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bdatw[9]_INST_0_i_73 
       (.I0(\stat_reg[0]_20 ),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(bank_sel),
        .I5(\i_/bdatw[12]_INST_0_i_64 [1]),
        .O(\grn_reg[1] ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(ccmd[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF5050505C)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(\ccmd[0]_INST_0_i_2_n_0 ),
        .I1(\ccmd[0]_INST_0_i_3_n_0 ),
        .I2(\ccmd[0]_INST_0_i_4_n_0 ),
        .I3(\ccmd[0]_INST_0_i_5_n_0 ),
        .I4(\ccmd[0]_INST_0_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(\ccmd[0]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(ir0[14]),
        .I1(ir0[15]),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(ir0[14]),
        .I1(ir0[12]),
        .I2(ir0[15]),
        .I3(\ccmd[0]_INST_0_i_23_n_0 ),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000008EA58E)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(ir0[11]),
        .I1(crdy),
        .I2(ir0[8]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\ccmd[4]_INST_0_i_12_n_0 ),
        .I5(\ccmd[0]_INST_0_i_24_n_0 ),
        .O(\ccmd[0]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h41)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[11]),
        .O(\ccmd[0]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(ir0[7]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F5F5F755D5555)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(ir0[3]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[6]),
        .I3(ir0[4]),
        .I4(ir0[7]),
        .I5(ir0[5]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hA0A0AAAAA3E0ABAA)) 
    \ccmd[0]_INST_0_i_19 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(ir0[5]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\ccmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h5444444454445444)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(ir0[15]),
        .I1(\ccmd[0]_INST_0_i_7_n_0 ),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(\ccmd[0]_INST_0_i_8_n_0 ),
        .I5(\ccmd[0]_INST_0_i_9_n_0 ),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFEFFFFFFFC)) 
    \ccmd[0]_INST_0_i_21 
       (.I0(ir0[9]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(ir0[10]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[6]),
        .I5(ir0[11]),
        .O(\ccmd[0]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_22 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[0]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \ccmd[0]_INST_0_i_23 
       (.I0(ir0[6]),
        .I1(ir0[4]),
        .I2(ir0[5]),
        .I3(ir0[7]),
        .I4(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .O(\ccmd[0]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF14101414)) 
    \ccmd[0]_INST_0_i_24 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[11]),
        .I5(\ccmd[0]_INST_0_i_25_n_0 ),
        .O(\ccmd[0]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFBFBFFFBFBFB)) 
    \ccmd[0]_INST_0_i_25 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[7]),
        .I5(crdy),
        .O(\ccmd[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFFFFFEF)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(\ccmd[0]_INST_0_i_1_1 ),
        .I5(ir0[15]),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAA2A)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(ir0[13]),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\ccmd[0]_INST_0_i_11_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[12]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0001010104111011)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(\ccmd[0]_INST_0_i_12_n_0 ),
        .I1(\ccmd[0]_INST_0_i_1_2 ),
        .I2(ir0[1]),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(ir0[0]),
        .I5(ir0[3]),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h28882288)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(\ccmd[0]_INST_0_i_1_0 ),
        .I1(ir0[11]),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .I4(\sr_reg[15]_0 [5]),
        .O(\ccmd[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000210003)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(\sr_reg[15]_0 [7]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[12]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\ccmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAEAEAEAEAEAEA)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(\ccmd[0]_INST_0_i_15_n_0 ),
        .I1(\ccmd[0]_INST_0_i_16_n_0 ),
        .I2(\ccmd[0]_INST_0_i_17_n_0 ),
        .I3(\ccmd[0]_INST_0_i_18_n_0 ),
        .I4(\ccmd[0]_INST_0_i_19_n_0 ),
        .I5(fctl_n_94),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0FDFDFFF0F5F5)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(ir0[9]),
        .I2(\ccmd[0]_INST_0_i_21_n_0 ),
        .I3(\ccmd[0]_INST_0_i_22_n_0 ),
        .I4(ir0[11]),
        .I5(ir0[8]),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[1]_INST_0 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'h00000000AAAAFF03)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_3_n_0 ),
        .I2(\ccmd[1]_INST_0_i_4_n_0 ),
        .I3(\ccmd[1]_INST_0_i_5_n_0 ),
        .I4(\ccmd[1]_INST_0_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\ccmd[1]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .O(\ccmd[1]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[4]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(\ccmd[0]_INST_0_i_11_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(\ccmd[1]_INST_0_i_9_n_0 ),
        .O(\ccmd[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF4FFF1F1F4FFF3FF)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(ir0[10]),
        .I1(ir0[6]),
        .I2(\ccmd[1]_INST_0_i_19_n_0 ),
        .I3(crdy),
        .I4(ir0[7]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(ir0[13]),
        .I1(ir0[11]),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4044404440404000)) 
    \ccmd[1]_INST_0_i_15 
       (.I0(\ccmd[4]_INST_0_i_20_n_0 ),
        .I1(ir0[8]),
        .I2(crdy),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\ccmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000001100004213)) 
    \ccmd[1]_INST_0_i_16 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(ir0[9]),
        .O(\ccmd[1]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFBF23FF)) 
    \ccmd[1]_INST_0_i_17 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .I3(ir0[7]),
        .I4(ir0[5]),
        .O(\ccmd[1]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[1]_INST_0_i_18 
       (.I0(ir0[10]),
        .I1(ir0[8]),
        .O(\ccmd[1]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFF8F)) 
    \ccmd[1]_INST_0_i_19 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .O(\ccmd[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000EEE00000000)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(\ccmd[1]_INST_0_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_8_n_0 ),
        .I2(ir0[13]),
        .I3(ir0[15]),
        .I4(\rgf_selc0_rn_wb_reg[0] [2]),
        .I5(ir0[14]),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0009)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[15]),
        .I3(\ccmd[1]_INST_0_i_9_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFFFFF00AAFFBF)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(ir0[11]),
        .I1(crdy),
        .I2(\ccmd[4]_INST_0_i_16_n_0 ),
        .I3(ir0[13]),
        .I4(ir0[15]),
        .I5(ir0[14]),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0E000)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(\ccmd[1]_INST_0_i_10_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I2(\ccmd[1]_INST_0_i_11_n_0 ),
        .I3(ir0[2]),
        .I4(\rgf_selc0_rn_wb_reg[0] [2]),
        .I5(\ccmd[1]_INST_0_i_12_n_0 ),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[11]),
        .I3(ir0[15]),
        .O(\ccmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0F004F4F0F004F44)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(ir0[13]),
        .I1(ir0[15]),
        .I2(\ccmd[1]_INST_0_i_13_n_0 ),
        .I3(\ccmd[4]_INST_0_i_18_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\ccmd[4]_INST_0_i_12_n_0 ),
        .O(\ccmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA8A8A8A8A8A8)) 
    \ccmd[1]_INST_0_i_8 
       (.I0(\ccmd[1]_INST_0_i_14_n_0 ),
        .I1(\ccmd[1]_INST_0_i_15_n_0 ),
        .I2(\ccmd[1]_INST_0_i_16_n_0 ),
        .I3(\ccmd[1]_INST_0_i_17_n_0 ),
        .I4(\bcmd[2]_INST_0_i_8_n_0 ),
        .I5(\ccmd[1]_INST_0_i_18_n_0 ),
        .O(\ccmd[1]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(ir0[13]),
        .I1(ir0[11]),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(ccmd[2]));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF7)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\rgf_selc0_rn_wb_reg[0] [2]),
        .I4(\ccmd[2]_INST_0_i_2_n_0 ),
        .I5(\ccmd[2]_INST_0_i_3_n_0 ),
        .O(\ccmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h1FFFFFF11FF1FFF1)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(crdy),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(ir0[7]),
        .I5(ir0[6]),
        .O(\ccmd[2]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(ir0[6]),
        .I1(ir0[10]),
        .O(\ccmd[2]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00008000C0C08000)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(ir0[7]),
        .I2(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I3(ir0[6]),
        .I4(ir0[10]),
        .I5(ir0[9]),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000090)) 
    \ccmd[2]_INST_0_i_13 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[11]),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(ir0[10]),
        .I5(\ccmd[2]_INST_0_i_16_n_0 ),
        .O(\ccmd[2]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000077061706)) 
    \ccmd[2]_INST_0_i_14 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(\ccmd[2]_INST_0_i_17_n_0 ),
        .I3(\ccmd[2]_INST_0_i_18_n_0 ),
        .I4(ir0[0]),
        .I5(\ccmd[2]_INST_0_i_19_n_0 ),
        .O(\ccmd[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAEAAAAAA)) 
    \ccmd[2]_INST_0_i_16 
       (.I0(ir0[8]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(ir0[11]),
        .I3(ir0[10]),
        .I4(ir0[7]),
        .I5(ir0[9]),
        .O(\ccmd[2]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    \ccmd[2]_INST_0_i_17 
       (.I0(\ccmd[0]_INST_0_i_11_n_0 ),
        .I1(ir0[13]),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(ir0[0]),
        .I4(ir0[11]),
        .I5(ir0[5]),
        .O(\ccmd[2]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000054)) 
    \ccmd[2]_INST_0_i_18 
       (.I0(ir0[14]),
        .I1(crdy),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(ir0[15]),
        .I5(\ccmd[2]_INST_0_i_20_n_0 ),
        .O(\ccmd[2]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    \ccmd[2]_INST_0_i_19 
       (.I0(ir0[4]),
        .I1(ir0[10]),
        .I2(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I3(ir0[2]),
        .I4(ir0[6]),
        .I5(ir0[7]),
        .O(\ccmd[2]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFCAAFFFFFFAAFF)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(\ccmd[2]_INST_0_i_5_n_0 ),
        .I3(ir0[15]),
        .I4(ir0[14]),
        .I5(\ccmd[2]_INST_0_i_6_n_0 ),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \ccmd[2]_INST_0_i_20 
       (.I0(ir0[5]),
        .I1(ir0[11]),
        .I2(ir0[13]),
        .O(\ccmd[2]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(ir0[12]),
        .I1(\rgf_selc0_rn_wb_reg[0] [2]),
        .I2(\ccmd[2]_INST_0_i_7_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I4(\ccmd[2]_INST_0_i_8_n_0 ),
        .I5(\ccmd[2]_INST_0_i_9_n_0 ),
        .O(\ccmd[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h4044404040444044)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(ir0[11]),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(\ccmd[4]_INST_0_i_12_n_0 ),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA82AAAAAAA8)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(\stat[2]_i_12_n_0 ),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .I3(\ccmd[2]_INST_0_i_11_n_0 ),
        .I4(\ccmd[2]_INST_0_i_2_0 ),
        .I5(ir0[7]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FF02)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(ir0[11]),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(\ccmd[2]_INST_0_i_12_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(\ccmd[2]_INST_0_i_13_n_0 ),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF70500000)) 
    \ccmd[2]_INST_0_i_7 
       (.I0(ir0[13]),
        .I1(ir0[11]),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .I4(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I5(\ccmd[2]_INST_0_i_14_n_0 ),
        .O(\ccmd[2]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFFFFFFF)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(\bcmd[0]_INST_0_i_20_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [2]),
        .I2(\ccmd[2]_INST_0_i_3_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I4(ir0[13]),
        .I5(\ccmd[0]_INST_0_i_11_n_0 ),
        .O(\ccmd[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0400040000000400)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I2(ir0[13]),
        .I3(ir0[15]),
        .I4(ir0[11]),
        .I5(ir0[14]),
        .O(\ccmd[2]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(ccmd[3]));
  LUT6 #(
    .INIT(64'h00000000FFFFFF07)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(\ccmd[3]_INST_0_i_2_n_0 ),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(ir0[15]),
        .I4(\rgf_selc0_rn_wb_reg[0] [2]),
        .I5(\ccmd[3]_INST_0_i_4_n_0 ),
        .O(\ccmd[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBAABAAAAAAABA)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[8]),
        .I5(crdy),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[9]),
        .O(\ccmd[3]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF003030A8)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(\ccmd[3]_INST_0_i_3_0 ),
        .I1(ir0[0]),
        .I2(ir0[2]),
        .I3(ir0[1]),
        .I4(ir0[3]),
        .I5(ir0[6]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(crdy),
        .O(\ccmd[3]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCC4CCC7FFF7FFF7)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(\ccmd[3]_INST_0_i_20_n_0 ),
        .I1(ir0[12]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(crdy),
        .I5(\ccmd[3]_INST_0_i_21_n_0 ),
        .O(\ccmd[3]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_17 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .O(\ccmd[3]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[3]_INST_0_i_18 
       (.I0(ir0[11]),
        .I1(ir0[7]),
        .O(\ccmd[3]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFEFEFF)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(\ccmd[3]_INST_0_i_5_n_0 ),
        .I1(\ccmd[3]_INST_0_i_6_n_0 ),
        .I2(\ccmd[3]_INST_0_i_7_n_0 ),
        .I3(\ccmd[3]_INST_0_i_8_n_0 ),
        .I4(\ccmd[3]_INST_0_i_9_n_0 ),
        .I5(\ccmd[3]_INST_0_i_10_n_0 ),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[3]_INST_0_i_20 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .O(\ccmd[3]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \ccmd[3]_INST_0_i_21 
       (.I0(ir0[7]),
        .I1(ir0[8]),
        .I2(ir0[4]),
        .I3(ir0[5]),
        .O(\ccmd[3]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040404000)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(\ccmd[3]_INST_0_i_11_n_0 ),
        .I1(\ccmd[3]_INST_0_i_12_n_0 ),
        .I2(\ccmd[3]_INST_0_i_13_n_0 ),
        .I3(\ccmd[4]_INST_0_i_15_n_0 ),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\ccmd[3]_INST_0_i_15_n_0 ),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0CC04C0000000000)) 
    \ccmd[3]_INST_0_i_4 
       (.I0(ir0[11]),
        .I1(ctl_fetch0_fl_reg_0),
        .I2(ir0[13]),
        .I3(ir0[14]),
        .I4(ir0[12]),
        .I5(ir0[15]),
        .O(\ccmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\ccmd[4]_INST_0_i_12_n_0 ),
        .I2(crdy),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(ir0[11]),
        .I5(\ccmd[3]_INST_0_i_17_n_0 ),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000006000000000)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I3(ir0[7]),
        .I4(ir0[9]),
        .I5(ir0[11]),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h02220200)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .I1(ir0[11]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(crdy),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFDFFDDEEDDEE)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(ir0[10]),
        .I1(\ccmd[3]_INST_0_i_18_n_0 ),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\ccmd[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBBBFFFBFFFFB)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(ir0[5]),
        .I1(\stat[2]_i_12_n_0 ),
        .I2(ir0[3]),
        .I3(ir0[4]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(ir0[6]),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(ccmd[4]));
  LUT6 #(
    .INIT(64'h00000000AFAE00AE)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(\ccmd[4]_INST_0_i_3_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\ccmd[4]_INST_0_i_5_n_0 ),
        .I3(ir0[11]),
        .I4(\ccmd[4]_INST_0_i_6_n_0 ),
        .I5(\ccmd[4]_INST_0_i_7_n_0 ),
        .O(\stat_reg[0]_3 ));
  LUT4 #(
    .INIT(16'h9DDD)) 
    \ccmd[4]_INST_0_i_11 
       (.I0(ir0[15]),
        .I1(ir0[12]),
        .I2(ir0[8]),
        .I3(ir0[7]),
        .O(\ccmd[4]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \ccmd[4]_INST_0_i_12 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .I4(ir0[13]),
        .I5(ir0[12]),
        .O(\ccmd[4]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[4]_INST_0_i_13 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .O(\ccmd[4]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hAA02)) 
    \ccmd[4]_INST_0_i_14 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(ir0[3]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .O(\ccmd[4]_INST_0_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[4]_INST_0_i_15 
       (.I0(ir0[14]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .O(\ccmd[4]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \ccmd[4]_INST_0_i_16 
       (.I0(ir0[4]),
        .I1(ir0[10]),
        .I2(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I3(ir0[2]),
        .I4(ir0[6]),
        .I5(\fadr[15]_INST_0_i_18_n_0 ),
        .O(\ccmd[4]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \ccmd[4]_INST_0_i_17 
       (.I0(ir0[9]),
        .I1(crdy),
        .O(\ccmd[4]_INST_0_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \ccmd[4]_INST_0_i_18 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\ccmd[4]_INST_0_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \ccmd[4]_INST_0_i_19 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(ir0[9]),
        .O(\ccmd[4]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFF45FF45FFFFFF55)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(\ccmd[4]_INST_0_i_8_n_0 ),
        .I1(\ccmd[4]_INST_0_i_9_n_0 ),
        .I2(crdy),
        .I3(ccmd_4_sn_1),
        .I4(\ccmd[4]_INST_0_i_11_n_0 ),
        .I5(\ccmd[4]_INST_0_i_12_n_0 ),
        .O(\ccmd[4]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \ccmd[4]_INST_0_i_20 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .O(\ccmd[4]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h000000004F000000)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(\ccmd[4]_INST_0_i_14_n_0 ),
        .I3(\ccmd[4]_INST_0_i_15_n_0 ),
        .I4(\ccmd[4]_INST_0_i_16_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_3_n_0 ),
        .O(\ccmd[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00FF001700)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(ir0[8]),
        .I1(ir0[10]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(\bcmd[0]_INST_0_i_9_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\ccmd[4]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0010033011113333)) 
    \ccmd[4]_INST_0_i_5 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(ir0[11]),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(ir0[7]),
        .I4(crdy),
        .I5(\ccmd[4]_INST_0_i_18_n_0 ),
        .O(\ccmd[4]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0080008888800080)) 
    \ccmd[4]_INST_0_i_6 
       (.I0(\ccmd[4]_INST_0_i_19_n_0 ),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .I2(crdy),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(ir0[7]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\ccmd[4]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[4]_INST_0_i_7 
       (.I0(ir0[15]),
        .I1(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(\ccmd[4]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000003300001033)) 
    \ccmd[4]_INST_0_i_8 
       (.I0(\ccmd[4]_INST_0_i_20_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(ir0[6]),
        .I3(ir0[12]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\ccmd[4]_INST_0_i_12_n_0 ),
        .O(\ccmd[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h9999989888989898)) 
    \ccmd[4]_INST_0_i_9 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(ir0[9]),
        .O(\ccmd[4]_INST_0_i_9_n_0 ));
  FDRE ctl_bcc_take0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take0_fl_reg_0),
        .Q(ctl_bcc_take0_fl),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE ctl_bcc_take1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take1_fl_reg_0),
        .Q(ctl_bcc_take1_fl),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE ctl_fetch0_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch0),
        .Q(ctl_fetch0_fl),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'h01)) 
    ctl_fetch1_fl_i_20
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .O(ctl_fetch1_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch1_fl_i_36
       (.I0(ir1[4]),
        .I1(ir1[5]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(ir1[7]),
        .O(ctl_fetch1_fl_i_36_n_0));
  FDRE ctl_fetch1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch1),
        .Q(ctl_fetch1_fl),
        .R(\<const0> ));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_ext_fl_i_1
       (.I0(fctl_n_67),
        .O(ctl_fetch_ext_fl_i_1_n_0));
  FDRE ctl_fetch_ext_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_ext_fl_i_1_n_0),
        .Q(ctl_fetch_ext_fl),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hFB)) 
    \eir_fl[15]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .I2(fch_irq_lev0),
        .O(\eir_fl[15]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(irq_vec[0]),
        .I1(fch_irq_lev0),
        .I2(eir[1]),
        .O(\eir_fl[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(irq_vec[1]),
        .I1(fch_irq_lev0),
        .I2(eir[2]),
        .O(\eir_fl[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(irq_vec[2]),
        .I1(fch_irq_lev0),
        .I2(eir[3]),
        .O(\eir_fl[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(irq_vec[3]),
        .I1(fch_irq_lev0),
        .I2(eir[4]),
        .O(\eir_fl[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(irq_vec[4]),
        .I1(fch_irq_lev0),
        .I2(eir[5]),
        .O(\eir_fl[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \eir_fl[6]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .O(\eir_fl[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_2 
       (.I0(irq_vec[5]),
        .I1(fch_irq_lev0),
        .I2(eir[6]),
        .O(\eir_fl[6]_i_2_n_0 ));
  FDRE \eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[0]),
        .Q(\eir_fl_reg_n_0_[0] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[10]),
        .Q(\eir_fl_reg_n_0_[10] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[11]),
        .Q(\eir_fl_reg_n_0_[11] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[12]),
        .Q(\eir_fl_reg_n_0_[12] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[13]),
        .Q(\eir_fl_reg_n_0_[13] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[14]),
        .Q(\eir_fl_reg_n_0_[14] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[15]),
        .Q(\eir_fl_reg_n_0_[15] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[1]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[1] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[2]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[2] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[3]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[3] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[4]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[4] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[5]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[5] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[6]_i_2_n_0 ),
        .Q(\eir_fl_reg_n_0_[6] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[7]),
        .Q(\eir_fl_reg_n_0_[7] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[8]),
        .Q(\eir_fl_reg_n_0_[8] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[9]),
        .Q(\eir_fl_reg_n_0_[9] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBFFF)) 
    \fadr[15]_INST_0_i_11 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I3(\fadr[15]_INST_0_i_18_n_0 ),
        .I4(ir0[4]),
        .I5(ir0[6]),
        .O(\fadr[15]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_13 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .O(\fadr[15]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_16 
       (.I0(ir1[5]),
        .I1(ir1[7]),
        .O(\fadr[15]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_18 
       (.I0(ir0[5]),
        .I1(ir0[7]),
        .O(\fadr[15]_INST_0_i_18_n_0 ));
  FDRE fadr_1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fadr[1]),
        .Q(fadr_1_fl),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(fch_irq_lev0),
        .I2(fch_irq_lev[0]),
        .O(\fch_irq_lev[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(fch_irq_lev0),
        .I2(fch_irq_lev[1]),
        .O(\fch_irq_lev[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00002000AAAAAAAA)) 
    \fch_irq_lev[1]_i_2 
       (.I0(fch_irq_req),
        .I1(\stat_reg[0]_48 ),
        .I2(brdy),
        .I3(fctl_n_89),
        .I4(\fch_irq_lev[1]_i_3_n_0 ),
        .I5(\fch_irq_lev[1]_i_4_n_0 ),
        .O(fch_irq_lev0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \fch_irq_lev[1]_i_3 
       (.I0(\rgf_selc1_rn_wb[0]_i_22_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[4]),
        .I3(\rgf_selc1_wb_reg[1] [2]),
        .I4(ir1[11]),
        .I5(\fch_irq_lev[1]_i_5_n_0 ),
        .O(\fch_irq_lev[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    \fch_irq_lev[1]_i_4 
       (.I0(\rgf_selc0_wb[0]_i_5_n_0 ),
        .I1(\fch_irq_lev[1]_i_2_0 ),
        .I2(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I3(ir0[4]),
        .I4(ir0[1]),
        .I5(\sr[13]_i_8_n_0 ),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \fch_irq_lev[1]_i_5 
       (.I0(ir1[3]),
        .I1(ir1[0]),
        .I2(ir1[1]),
        .O(\fch_irq_lev[1]_i_5_n_0 ));
  FDRE \fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[0]_i_1_n_0 ),
        .Q(fch_irq_lev[0]),
        .R(SR));
  FDRE \fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[1]_i_1_n_0 ),
        .Q(fch_irq_lev[1]),
        .R(SR));
  FDRE fch_irq_req_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(fch_irq_req_fl),
        .R(\<const0> ));
  FDRE fch_issu1_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_issu1_ir),
        .Q(fch_issu1_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'hF7570000FFFFFFFF)) 
    fch_issu1_inferred_i_100
       (.I0(fdatx[10]),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fch_issu1_inferred_i_97_n_0),
        .I4(fch_issu1_inferred_i_168_n_0),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_100_n_0));
  LUT6 #(
    .INIT(64'h44C0FFFFFFFFFFFF)) 
    fch_issu1_inferred_i_101
       (.I0(fch_issu1_inferred_i_169_n_0),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(fdatx[12]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_101_n_0));
  LUT6 #(
    .INIT(64'hAAFEAAAAAABAAAAA)) 
    fch_issu1_inferred_i_102
       (.I0(fch_issu1_inferred_i_101_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .I5(fdatx[2]),
        .O(fch_issu1_inferred_i_102_n_0));
  LUT6 #(
    .INIT(64'h5DDDDDDD55D5D5D5)) 
    fch_issu1_inferred_i_103
       (.I0(fch_issu1_inferred_i_168_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[8]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[2]),
        .O(fch_issu1_inferred_i_103_n_0));
  LUT6 #(
    .INIT(64'hAA3F0FFF00000000)) 
    fch_issu1_inferred_i_104
       (.I0(fch_issu1_inferred_i_170_n_0),
        .I1(fdatx[1]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .I5(fch_issu1_inferred_i_171_n_0),
        .O(fch_issu1_inferred_i_104_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBBFFFFFFF)) 
    fch_issu1_inferred_i_105
       (.I0(fdatx[11]),
        .I1(fdatx[12]),
        .I2(fch_issu1_inferred_i_161_n_0),
        .I3(fdatx[9]),
        .I4(fdatx[7]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_105_n_0));
  LUT6 #(
    .INIT(64'hCCCCCCCC08C8C8C8)) 
    fch_issu1_inferred_i_106
       (.I0(fdatx[1]),
        .I1(fdatx[10]),
        .I2(fdatx[8]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_106_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_107
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_107_n_0));
  LUT6 #(
    .INIT(64'h0A002A8002020202)) 
    fch_issu1_inferred_i_108
       (.I0(fdatx[8]),
        .I1(fdatx[4]),
        .I2(fdatx[5]),
        .I3(fdatx[7]),
        .I4(fdatx[3]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_108_n_0));
  LUT6 #(
    .INIT(64'h00000000DDDFDDDD)) 
    fch_issu1_inferred_i_109
       (.I0(fdat[3]),
        .I1(fdat[9]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fch_issu1_inferred_i_172_n_0),
        .O(fch_issu1_inferred_i_109_n_0));
  LUT6 #(
    .INIT(64'hFFFF3F703058FFFF)) 
    fch_issu1_inferred_i_110
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[11]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_110_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    fch_issu1_inferred_i_111
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .O(fch_issu1_inferred_i_111_n_0));
  LUT6 #(
    .INIT(64'h0FDDFFDDFFDDFFDD)) 
    fch_issu1_inferred_i_113
       (.I0(fdatx[3]),
        .I1(fch_issu1_inferred_i_173_n_0),
        .I2(fdatx[0]),
        .I3(fdatx[9]),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_174_n_0),
        .O(fch_issu1_inferred_i_113_n_0));
  LUT4 #(
    .INIT(16'hCAF7)) 
    fch_issu1_inferred_i_114
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .O(fch_issu1_inferred_i_114_n_0));
  LUT6 #(
    .INIT(64'h0515444455555555)) 
    fch_issu1_inferred_i_115
       (.I0(fdatx[11]),
        .I1(fdatx[9]),
        .I2(fdatx[6]),
        .I3(fdatx[7]),
        .I4(fdatx[8]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_115_n_0));
  LUT6 #(
    .INIT(64'hEEE0E0E0E0E0E0E0)) 
    fch_issu1_inferred_i_116
       (.I0(fch_issu1_inferred_i_107_n_0),
        .I1(fdatx[5]),
        .I2(fch_issu1_inferred_i_175_n_0),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .I5(fch_issu1_inferred_i_176_n_0),
        .O(fch_issu1_inferred_i_116_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    fch_issu1_inferred_i_117
       (.I0(fch_issu1_inferred_i_54_n_0),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .O(fch_issu1_inferred_i_117_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFFFBF)) 
    fch_issu1_inferred_i_118
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_177_n_0),
        .I2(fdatx_5_sn_1),
        .I3(fdatx[6]),
        .I4(fch_issu1_inferred_i_135_n_0),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_118_n_0));
  LUT4 #(
    .INIT(16'hEAAA)) 
    fch_issu1_inferred_i_119
       (.I0(fdatx[10]),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .I3(fdatx[14]),
        .O(fch_issu1_inferred_i_119_n_0));
  LUT6 #(
    .INIT(64'h5555555155555555)) 
    fch_issu1_inferred_i_120
       (.I0(fdat[15]),
        .I1(fdat[0]),
        .I2(fdat[12]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fch_issu1_inferred_i_126_n_0),
        .O(fch_issu1_inferred_i_120_n_0));
  LUT6 #(
    .INIT(64'hA2A2A2A0A2A2A2A2)) 
    fch_issu1_inferred_i_121
       (.I0(fch_issu1_inferred_i_178_n_0),
        .I1(fdat[5]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_121_n_0));
  LUT6 #(
    .INIT(64'h80FFFFFF80000000)) 
    fch_issu1_inferred_i_122
       (.I0(fdat[6]),
        .I1(fdat[9]),
        .I2(fch_issu1_inferred_i_179_n_0),
        .I3(fdat[10]),
        .I4(fdat[11]),
        .I5(fdat[5]),
        .O(fch_issu1_inferred_i_122_n_0));
  LUT6 #(
    .INIT(64'h0000000003233333)) 
    fch_issu1_inferred_i_123
       (.I0(fdat[11]),
        .I1(fadr_1_fl),
        .I2(fdat[12]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_123_n_0));
  LUT6 #(
    .INIT(64'h4474F0F0F0F0F0F0)) 
    fch_issu1_inferred_i_124
       (.I0(fch_issu1_inferred_i_180_n_0),
        .I1(fdat[9]),
        .I2(fdat[4]),
        .I3(\nir_id[14]_i_12_n_0 ),
        .I4(fdat[11]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_124_n_0));
  LUT6 #(
    .INIT(64'h0000FF00D5D5D5D5)) 
    fch_issu1_inferred_i_125
       (.I0(fdatx[4]),
        .I1(fch_issu1_inferred_i_161_n_0),
        .I2(fdatx[7]),
        .I3(fch_issu1_inferred_i_181_n_0),
        .I4(fch_issu1_inferred_i_182_n_0),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_125_n_0));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    fch_issu1_inferred_i_126
       (.I0(fdat[9]),
        .I1(\nir_id[19]_i_7_n_0 ),
        .I2(fch_issu1_inferred_i_183_n_0),
        .I3(fdat_5_sn_1),
        .I4(fdat[2]),
        .I5(fdat[3]),
        .O(fch_issu1_inferred_i_126_n_0));
  LUT6 #(
    .INIT(64'hFFEFFFFF1F9F0000)) 
    fch_issu1_inferred_i_127
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[8]),
        .I3(fdat[3]),
        .I4(fdat[9]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_127_n_0));
  LUT6 #(
    .INIT(64'h6900EFEE69006F66)) 
    fch_issu1_inferred_i_128
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .I4(fdat[6]),
        .I5(\nir_id[17]_i_6_n_0 ),
        .O(fch_issu1_inferred_i_128_n_0));
  LUT6 #(
    .INIT(64'h8F88888888888888)) 
    fch_issu1_inferred_i_129
       (.I0(fdat[11]),
        .I1(fdat[15]),
        .I2(fdat[5]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_129_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000F700)) 
    fch_issu1_inferred_i_130
       (.I0(fch_issu1_inferred_i_184_n_0),
        .I1(fdat[8]),
        .I2(fdat[15]),
        .I3(fdat[14]),
        .I4(fdat[11]),
        .I5(fch_issu1_inferred_i_142_n_0),
        .O(fch_issu1_inferred_i_130_n_0));
  LUT6 #(
    .INIT(64'h91996060F1F9F1F9)) 
    fch_issu1_inferred_i_131
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .I2(fdatx[6]),
        .I3(fch_issu1_inferred_i_154_n_0),
        .I4(fdatx[10]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_131_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000E600)) 
    fch_issu1_inferred_i_132
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[8]),
        .I4(fdatx[7]),
        .I5(fch_issu1_inferred_i_185_n_0),
        .O(fch_issu1_inferred_i_132_n_0));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    fch_issu1_inferred_i_133
       (.I0(fdatx[4]),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[3]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_133_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000BF00)) 
    fch_issu1_inferred_i_134
       (.I0(fdatx[15]),
        .I1(fdatx[8]),
        .I2(fch_issu1_inferred_i_186_n_0),
        .I3(fdatx[14]),
        .I4(fdatx[11]),
        .I5(fch_issu1_inferred_i_140_n_0),
        .O(fch_issu1_inferred_i_134_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    fch_issu1_inferred_i_135
       (.I0(fdatx[11]),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .O(fch_issu1_inferred_i_135_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    fch_issu1_inferred_i_136
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[2]),
        .I3(fdatx[3]),
        .O(fch_issu1_inferred_i_136_n_0));
  LUT5 #(
    .INIT(32'h00080000)) 
    fch_issu1_inferred_i_137
       (.I0(fdatx[6]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[7]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_137_n_0));
  LUT6 #(
    .INIT(64'hFFEFEFFEAAAAAAAA)) 
    fch_issu1_inferred_i_138
       (.I0(fch_issu1_inferred_i_187_n_0),
        .I1(fdatx[6]),
        .I2(fdatx[7]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .I5(fch_issu1_inferred_i_107_n_0),
        .O(fch_issu1_inferred_i_138_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_139
       (.I0(fdatx[8]),
        .I1(fdatx[10]),
        .O(fch_issu1_inferred_i_139_n_0));
  LUT6 #(
    .INIT(64'h5D55555555555555)) 
    fch_issu1_inferred_i_14
       (.I0(fch_issu1_inferred_i_43_n_0),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[11]),
        .I4(fdat[8]),
        .I5(fch_issu1_inferred_i_44_n_0),
        .O(fch_issu1_inferred_i_14_n_0));
  LUT5 #(
    .INIT(32'h44CC7FDD)) 
    fch_issu1_inferred_i_140
       (.I0(fdatx[13]),
        .I1(fdatx[15]),
        .I2(fdatx[11]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .O(fch_issu1_inferred_i_140_n_0));
  LUT6 #(
    .INIT(64'h000000000441FFFF)) 
    fch_issu1_inferred_i_141
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(\nir_id[16]_i_3_n_0 ),
        .I5(fch_issu1_inferred_i_188_n_0),
        .O(fch_issu1_inferred_i_141_n_0));
  LUT5 #(
    .INIT(32'h44CC7FDD)) 
    fch_issu1_inferred_i_142
       (.I0(fdat[13]),
        .I1(fdat[15]),
        .I2(fdat[11]),
        .I3(fdat[14]),
        .I4(fdat[12]),
        .O(fch_issu1_inferred_i_142_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_143
       (.I0(fdat[8]),
        .I1(fdat[10]),
        .O(fch_issu1_inferred_i_143_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_145
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .O(fch_issu1_inferred_i_145_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_146
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_146_n_0));
  LUT4 #(
    .INIT(16'h0040)) 
    fch_issu1_inferred_i_147
       (.I0(fdat[7]),
        .I1(fdat[5]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .O(fch_issu1_inferred_i_147_n_0));
  LUT6 #(
    .INIT(64'hFCECFC4CFCECFCEC)) 
    fch_issu1_inferred_i_148
       (.I0(fdatx[9]),
        .I1(fdatx[5]),
        .I2(fch_issu1_inferred_i_107_n_0),
        .I3(fch_issu1_inferred_i_152_n_0),
        .I4(fch_issu1_inferred_i_189_n_0),
        .I5(fch_issu1_inferred_i_190_n_0),
        .O(fch_issu1_inferred_i_148_n_0));
  LUT5 #(
    .INIT(32'hAAAA8AAA)) 
    fch_issu1_inferred_i_149
       (.I0(fdatx[15]),
        .I1(fdatx[12]),
        .I2(fdatx[11]),
        .I3(fdatx[13]),
        .I4(fdatx[14]),
        .O(fch_issu1_inferred_i_149_n_0));
  LUT6 #(
    .INIT(64'h555555555555D555)) 
    fch_issu1_inferred_i_15
       (.I0(fch_issu1_inferred_i_45_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[6]),
        .I3(fch_issu1_inferred_i_46_n_0),
        .I4(fdatx[9]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_15_n_0));
  LUT6 #(
    .INIT(64'h110F0000110F000F)) 
    fch_issu1_inferred_i_150
       (.I0(fdatx[0]),
        .I1(fch_issu1_inferred_i_189_n_0),
        .I2(fdatx[3]),
        .I3(fdatx[9]),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_97_n_0),
        .O(fch_issu1_inferred_i_150_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0B00FFFF)) 
    fch_issu1_inferred_i_151
       (.I0(fdatx[6]),
        .I1(fdatx[3]),
        .I2(fch_issu1_inferred_i_182_n_0),
        .I3(fch_issu1_inferred_i_191_n_0),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_192_n_0),
        .O(fch_issu1_inferred_i_151_n_0));
  LUT4 #(
    .INIT(16'h1000)) 
    fch_issu1_inferred_i_152
       (.I0(fdatx[9]),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .O(fch_issu1_inferred_i_152_n_0));
  LUT6 #(
    .INIT(64'hFFFFF7FFFFFFFEFF)) 
    fch_issu1_inferred_i_153
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[7]),
        .I3(fdatx[8]),
        .I4(fdatx[3]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_153_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_154
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(fch_issu1_inferred_i_154_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_155
       (.I0(fdatx[5]),
        .I1(fdatx[3]),
        .O(fch_issu1_inferred_i_155_n_0));
  LUT6 #(
    .INIT(64'h4400044044400440)) 
    fch_issu1_inferred_i_156
       (.I0(fdatx[11]),
        .I1(fdatx[10]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_156_n_0));
  LUT6 #(
    .INIT(64'h0E0C0000020E0000)) 
    fch_issu1_inferred_i_157
       (.I0(fdatx[7]),
        .I1(fdatx[8]),
        .I2(fdatx[10]),
        .I3(fdatx[11]),
        .I4(fdatx[9]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_157_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    fch_issu1_inferred_i_158
       (.I0(fdat[14]),
        .I1(fdat[13]),
        .I2(fdat[12]),
        .O(fch_issu1_inferred_i_158_n_0));
  LUT6 #(
    .INIT(64'h0000000301020202)) 
    fch_issu1_inferred_i_159
       (.I0(fdatx[1]),
        .I1(fch_issu1_inferred_i_193_n_0),
        .I2(fdatx[13]),
        .I3(fdatx[3]),
        .I4(fdatx[2]),
        .I5(fdatx[0]),
        .O(fch_issu1_inferred_i_159_n_0));
  LUT5 #(
    .INIT(32'h08000008)) 
    fch_issu1_inferred_i_16
       (.I0(fch_issu1_inferred_i_47_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[11]),
        .O(fch_issu1_inferred_i_16_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_160
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_160_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_161
       (.I0(fdatx[8]),
        .I1(fdatx[6]),
        .O(fch_issu1_inferred_i_161_n_0));
  LUT6 #(
    .INIT(64'h5EFFFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_162
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[10]),
        .I3(fdatx[12]),
        .I4(fdatx[11]),
        .I5(fdatx[8]),
        .O(fch_issu1_inferred_i_162_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_163
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .O(fch_issu1_inferred_i_163_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    fch_issu1_inferred_i_164
       (.I0(fdatx[14]),
        .I1(fdatx[13]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[8]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_164_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    fch_issu1_inferred_i_165
       (.I0(fdatx[11]),
        .I1(fdatx[10]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .O(fch_issu1_inferred_i_165_n_0));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFFBFFFF)) 
    fch_issu1_inferred_i_167
       (.I0(fch_issu1_inferred_i_165_n_0),
        .I1(fdatx_5_sn_1),
        .I2(fdatx[2]),
        .I3(fdatx[3]),
        .I4(fdatx[0]),
        .I5(fdatx[1]),
        .O(fch_issu1_inferred_i_167_n_0));
  LUT6 #(
    .INIT(64'h000000004A0A0000)) 
    fch_issu1_inferred_i_168
       (.I0(fdatx[10]),
        .I1(fdatx[7]),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_161_n_0),
        .I4(fdatx[12]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_168_n_0));
  LUT6 #(
    .INIT(64'hAA0A2000AAA8000A)) 
    fch_issu1_inferred_i_169
       (.I0(fdatx[8]),
        .I1(fdatx[3]),
        .I2(fdatx[4]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_169_n_0));
  LUT6 #(
    .INIT(64'h0020000000000020)) 
    fch_issu1_inferred_i_17
       (.I0(fdat_12_sn_1),
        .I1(fdat[15]),
        .I2(fdat[10]),
        .I3(fdat[9]),
        .I4(fdat[8]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'h0400C0C000C0C00C)) 
    fch_issu1_inferred_i_170
       (.I0(fdatx[3]),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .I4(fdatx[5]),
        .I5(fdatx[4]),
        .O(fch_issu1_inferred_i_170_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_171
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_171_n_0));
  LUT6 #(
    .INIT(64'h000000005FDD5DDD)) 
    fch_issu1_inferred_i_172
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[3]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fch_issu1_inferred_i_194_n_0),
        .O(fch_issu1_inferred_i_172_n_0));
  LUT3 #(
    .INIT(8'h10)) 
    fch_issu1_inferred_i_173
       (.I0(fdatx[6]),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .O(fch_issu1_inferred_i_173_n_0));
  LUT5 #(
    .INIT(32'h08C80B8B)) 
    fch_issu1_inferred_i_174
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[5]),
        .I3(fdatx[3]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_174_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0F00DF00)) 
    fch_issu1_inferred_i_175
       (.I0(fdatx_5_sn_1),
        .I1(fdatx[2]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .I5(fch_issu1_inferred_i_195_n_0),
        .O(fch_issu1_inferred_i_175_n_0));
  LUT6 #(
    .INIT(64'hFABBFBBBFABAFABA)) 
    fch_issu1_inferred_i_176
       (.I0(fdatx[2]),
        .I1(fdatx[7]),
        .I2(fdatx[3]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_176_n_0));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    fch_issu1_inferred_i_177
       (.I0(fdatx[12]),
        .I1(fdatx[7]),
        .I2(fch_issu1_inferred_i_196_n_0),
        .I3(fdatx[1]),
        .I4(fdatx[13]),
        .I5(fdatx[0]),
        .O(fch_issu1_inferred_i_177_n_0));
  LUT6 #(
    .INIT(64'hB3B3B3B3B3B3B3F3)) 
    fch_issu1_inferred_i_178
       (.I0(fdat[6]),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(fdat[2]),
        .I4(fdat[5]),
        .I5(fdat[4]),
        .O(fch_issu1_inferred_i_178_n_0));
  LUT6 #(
    .INIT(64'hFABBFBBBFABAFABA)) 
    fch_issu1_inferred_i_179
       (.I0(fdat[2]),
        .I1(fdat[7]),
        .I2(fdat[3]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_179_n_0));
  LUT6 #(
    .INIT(64'h0000DD000000F000)) 
    fch_issu1_inferred_i_180
       (.I0(fch_issu1_inferred_i_197_n_0),
        .I1(fch_issu1_inferred_i_147_n_0),
        .I2(fdat_5_sn_1),
        .I3(fdat[8]),
        .I4(fdat[1]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_180_n_0));
  LUT6 #(
    .INIT(64'h0000FFFF0ECCFFFF)) 
    fch_issu1_inferred_i_181
       (.I0(fdatx[4]),
        .I1(fdatx[7]),
        .I2(fdatx[3]),
        .I3(fdatx[5]),
        .I4(fdatx[6]),
        .I5(fdatx[1]),
        .O(fch_issu1_inferred_i_181_n_0));
  LUT5 #(
    .INIT(32'h5F5F5F4F)) 
    fch_issu1_inferred_i_182
       (.I0(fdatx[6]),
        .I1(fdatx[1]),
        .I2(fdatx[8]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_182_n_0));
  LUT4 #(
    .INIT(16'h0004)) 
    fch_issu1_inferred_i_183
       (.I0(fdat[8]),
        .I1(fdat[1]),
        .I2(fdat[11]),
        .I3(fdat[10]),
        .O(fch_issu1_inferred_i_183_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_184
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_184_n_0));
  LUT6 #(
    .INIT(64'hFF40FF40FF00FFFF)) 
    fch_issu1_inferred_i_185
       (.I0(fdatx[5]),
        .I1(fdatx[6]),
        .I2(fdatx[8]),
        .I3(fch_issu1_inferred_i_198_n_0),
        .I4(fdatx[7]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_185_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_186
       (.I0(fdatx[10]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_186_n_0));
  LUT6 #(
    .INIT(64'hCCCFDFFFFFCFDFFF)) 
    fch_issu1_inferred_i_187
       (.I0(fdatx[7]),
        .I1(fdatx[15]),
        .I2(fdatx[6]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_187_n_0));
  LUT6 #(
    .INIT(64'hABBBBBFFEFFFBBFF)) 
    fch_issu1_inferred_i_188
       (.I0(fdat[15]),
        .I1(fdat[9]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_188_n_0));
  LUT5 #(
    .INIT(32'h55FFF57E)) 
    fch_issu1_inferred_i_189
       (.I0(fdatx[6]),
        .I1(fdatx[4]),
        .I2(fdatx[5]),
        .I3(fdatx[7]),
        .I4(fdatx[3]),
        .O(fch_issu1_inferred_i_189_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_190
       (.I0(fdatx[8]),
        .I1(fdatx[2]),
        .O(fch_issu1_inferred_i_190_n_0));
  LUT6 #(
    .INIT(64'h000000000008FFFF)) 
    fch_issu1_inferred_i_191
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[1]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_191_n_0));
  LUT6 #(
    .INIT(64'h00000000D0000000)) 
    fch_issu1_inferred_i_192
       (.I0(fdatx[5]),
        .I1(fdatx[3]),
        .I2(fdatx[6]),
        .I3(fdatx[7]),
        .I4(fdatx[8]),
        .I5(fdatx[1]),
        .O(fch_issu1_inferred_i_192_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    fch_issu1_inferred_i_193
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[9]),
        .I3(fdatx[7]),
        .O(fch_issu1_inferred_i_193_n_0));
  LUT6 #(
    .INIT(64'h0EFFFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_194
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .I2(fdat[6]),
        .I3(fdat[0]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_194_n_0));
  LUT6 #(
    .INIT(64'h33333333BBBBBBFB)) 
    fch_issu1_inferred_i_195
       (.I0(fdatx[5]),
        .I1(fch_issu1_inferred_i_107_n_0),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .I4(fdatx[8]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_195_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_196
       (.I0(fdatx[3]),
        .I1(fdatx[2]),
        .O(fch_issu1_inferred_i_196_n_0));
  LUT3 #(
    .INIT(8'h8F)) 
    fch_issu1_inferred_i_197
       (.I0(fdat[5]),
        .I1(fdat[3]),
        .I2(fdat[7]),
        .O(fch_issu1_inferred_i_197_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_198
       (.I0(fdatx[15]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_198_n_0));
  LUT4 #(
    .INIT(16'h0080)) 
    fch_issu1_inferred_i_25
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fch_issu1_inferred_i_56_n_0),
        .O(fch_issu1_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'h400040C040004000)) 
    fch_issu1_inferred_i_26
       (.I0(fch_issu1_inferred_i_57_n_0),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[9]),
        .I4(fdat[8]),
        .I5(fch_issu1_inferred_i_58_n_0),
        .O(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF88082800)) 
    fch_issu1_inferred_i_27
       (.I0(fdat[15]),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(fadr_1_fl),
        .O(fch_issu1_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF5500C000)) 
    fch_issu1_inferred_i_36
       (.I0(fch_issu1_inferred_i_85_n_0),
        .I1(fch_issu1_inferred_i_86_n_0),
        .I2(fch_issu1_inferred_i_87_n_0),
        .I3(fdatx[11]),
        .I4(fdatx[10]),
        .I5(fch_issu1_inferred_i_88_n_0),
        .O(fch_issu1_inferred_i_36_n_0));
  LUT5 #(
    .INIT(32'h2A820AAA)) 
    fch_issu1_inferred_i_37
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[11]),
        .O(fch_issu1_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'h2000200020002002)) 
    fch_issu1_inferred_i_39
       (.I0(fch_issu1_inferred_i_92_n_0),
        .I1(fch_issu1_inferred_i_93_n_0),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'h000F0F0F0A0D0000)) 
    fch_issu1_inferred_i_43
       (.I0(fdat[8]),
        .I1(\nir_id[18]_i_8_n_0 ),
        .I2(fch_issu1_inferred_i_96_n_0),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_43_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_44
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_44_n_0));
  LUT6 #(
    .INIT(64'h0CFBF0F000000000)) 
    fch_issu1_inferred_i_45
       (.I0(fch_issu1_inferred_i_97_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[11]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .I5(fch_issu1_inferred_i_47_n_0),
        .O(fch_issu1_inferred_i_45_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_46
       (.I0(fdatx[11]),
        .I1(fdatx[10]),
        .O(fch_issu1_inferred_i_46_n_0));
  LUT4 #(
    .INIT(16'h4000)) 
    fch_issu1_inferred_i_47
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .O(fch_issu1_inferred_i_47_n_0));
  LUT6 #(
    .INIT(64'h888A8A8A8A8A8A8A)) 
    fch_issu1_inferred_i_49
       (.I0(fch_issu1_inferred_i_99_n_0),
        .I1(fch_issu1_inferred_i_100_n_0),
        .I2(fch_issu1_inferred_i_101_n_0),
        .I3(fdatx[10]),
        .I4(fdatx[0]),
        .I5(fch_issu1_inferred_i_87_n_0),
        .O(fch_issu1_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h4000400040004040)) 
    fch_issu1_inferred_i_51
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_104_n_0),
        .I4(fch_issu1_inferred_i_105_n_0),
        .I5(fch_issu1_inferred_i_106_n_0),
        .O(fch_issu1_inferred_i_51_n_0));
  LUT5 #(
    .INIT(32'hAAAAA2AA)) 
    fch_issu1_inferred_i_52
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[11]),
        .O(fch_issu1_inferred_i_52_n_0));
  LUT4 #(
    .INIT(16'hC060)) 
    fch_issu1_inferred_i_53
       (.I0(fdatx[11]),
        .I1(fdatx[12]),
        .I2(fdatx[14]),
        .I3(fdatx[13]),
        .O(fch_issu1_inferred_i_53_n_0));
  LUT6 #(
    .INIT(64'h000037F03508FFFF)) 
    fch_issu1_inferred_i_54
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[11]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'h00020000888A8888)) 
    fch_issu1_inferred_i_55
       (.I0(fch_issu1_inferred_i_107_n_0),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fch_issu1_inferred_i_108_n_0),
        .O(fch_issu1_inferred_i_55_n_0));
  LUT6 #(
    .INIT(64'h1135733117317731)) 
    fch_issu1_inferred_i_56
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_56_n_0));
  LUT6 #(
    .INIT(64'h0A002A8002020202)) 
    fch_issu1_inferred_i_57
       (.I0(fdat[8]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_57_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_58
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .O(fch_issu1_inferred_i_58_n_0));
  LUT6 #(
    .INIT(64'h4400440074F044F0)) 
    fch_issu1_inferred_i_62
       (.I0(fch_issu1_inferred_i_113_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[3]),
        .I3(fdatx[11]),
        .I4(fch_issu1_inferred_i_114_n_0),
        .I5(fch_issu1_inferred_i_115_n_0),
        .O(fch_issu1_inferred_i_62_n_0));
  LUT6 #(
    .INIT(64'hFFA80000FFA8FFA8)) 
    fch_issu1_inferred_i_63
       (.I0(fdatx[14]),
        .I1(fch_issu1_inferred_i_116_n_0),
        .I2(fch_issu1_inferred_i_117_n_0),
        .I3(fch_issu1_inferred_i_118_n_0),
        .I4(fch_issu1_inferred_i_119_n_0),
        .I5(fch_issu1_inferred_i_52_n_0),
        .O(fch_issu1_inferred_i_63_n_0));
  LUT6 #(
    .INIT(64'hAAAA2000AAAAAAAA)) 
    fch_issu1_inferred_i_64
       (.I0(fch_issu1_inferred_i_120_n_0),
        .I1(fch_issu1_inferred_i_121_n_0),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .I4(fch_issu1_inferred_i_122_n_0),
        .I5(fch_issu1_inferred_i_25_n_0),
        .O(fch_issu1_inferred_i_64_n_0));
  LUT5 #(
    .INIT(32'h03233333)) 
    fch_issu1_inferred_i_65
       (.I0(fdat[11]),
        .I1(fadr_1_fl),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .I4(fdat[12]),
        .O(fch_issu1_inferred_i_65_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_66
       (.I0(fadr_1_fl),
        .I1(fdat[15]),
        .O(fch_issu1_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'h0000AB00ABABABAB)) 
    fch_issu1_inferred_i_67
       (.I0(fch_issu1_inferred_i_123_n_0),
        .I1(fadr_1_fl),
        .I2(fdat[15]),
        .I3(fch_issu1_inferred_i_25_n_0),
        .I4(fch_issu1_inferred_i_124_n_0),
        .I5(fch_issu1_inferred_i_120_n_0),
        .O(fch_issu1_inferred_i_67_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    fch_issu1_inferred_i_68
       (.I0(fdatx[14]),
        .I1(fdatx[12]),
        .I2(fdatx[13]),
        .O(fdatx_14_sn_1));
  LUT6 #(
    .INIT(64'hFFFFBBFAAAAAAAAA)) 
    fch_issu1_inferred_i_69
       (.I0(fch_issu1_inferred_i_118_n_0),
        .I1(fch_issu1_inferred_i_125_n_0),
        .I2(fdatx[4]),
        .I3(fch_issu1_inferred_i_107_n_0),
        .I4(fch_issu1_inferred_i_117_n_0),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_69_n_0));
  LUT6 #(
    .INIT(64'h0000000002FFFFFF)) 
    fch_issu1_inferred_i_71
       (.I0(fch_issu1_inferred_i_127_n_0),
        .I1(fch_issu1_inferred_i_128_n_0),
        .I2(fch_issu1_inferred_i_129_n_0),
        .I3(fdat[14]),
        .I4(fdat[12]),
        .I5(fch_issu1_inferred_i_130_n_0),
        .O(fch_issu1_inferred_i_71_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFD000000)) 
    fch_issu1_inferred_i_72
       (.I0(fch_issu1_inferred_i_131_n_0),
        .I1(fch_issu1_inferred_i_132_n_0),
        .I2(fch_issu1_inferred_i_133_n_0),
        .I3(fdatx[12]),
        .I4(fdatx[14]),
        .I5(fch_issu1_inferred_i_134_n_0),
        .O(fch_issu1_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    fch_issu1_inferred_i_73
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_86_n_0),
        .I2(fdatx[1]),
        .I3(fdatx[13]),
        .I4(fch_issu1_inferred_i_135_n_0),
        .I5(fch_issu1_inferred_i_136_n_0),
        .O(fch_issu1_inferred_i_73_n_0));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    fch_issu1_inferred_i_76
       (.I0(fch_issu1_inferred_i_137_n_0),
        .I1(fdatx[9]),
        .I2(fdatx[15]),
        .I3(fdatx[8]),
        .I4(fdatx[10]),
        .I5(fdatx[12]),
        .O(fch_issu1_inferred_i_76_n_0));
  LUT6 #(
    .INIT(64'h0000000077FF70FF)) 
    fch_issu1_inferred_i_77
       (.I0(fch_issu1_inferred_i_138_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[11]),
        .I3(fdatx[14]),
        .I4(fch_issu1_inferred_i_139_n_0),
        .I5(fch_issu1_inferred_i_140_n_0),
        .O(fch_issu1_inferred_i_77_n_0));
  LUT6 #(
    .INIT(64'hF4F4F0F0F4FFF0F0)) 
    fch_issu1_inferred_i_78
       (.I0(fch_issu1_inferred_i_141_n_0),
        .I1(fdat[12]),
        .I2(fch_issu1_inferred_i_142_n_0),
        .I3(fdat[11]),
        .I4(fdat[14]),
        .I5(fch_issu1_inferred_i_143_n_0),
        .O(fch_issu1_inferred_i_78_n_0));
  LUT5 #(
    .INIT(32'hFFFF5CCC)) 
    fch_issu1_inferred_i_81
       (.I0(fch_issu1_inferred_i_150_n_0),
        .I1(fdatx[3]),
        .I2(fdatx[11]),
        .I3(fdatx[10]),
        .I4(fch_issu1_inferred_i_88_n_0),
        .O(fch_issu1_inferred_i_81_n_0));
  LUT6 #(
    .INIT(64'h000000000CC4CCCC)) 
    fch_issu1_inferred_i_82
       (.I0(fdatx[11]),
        .I1(fdatx[15]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[13]),
        .I5(fdatx[8]),
        .O(fch_issu1_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'h000000000CC4CCCC)) 
    fch_issu1_inferred_i_83
       (.I0(fdatx[11]),
        .I1(fdatx[15]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[13]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_83_n_0));
  LUT6 #(
    .INIT(64'h00000000080A00FF)) 
    fch_issu1_inferred_i_84
       (.I0(fch_issu1_inferred_i_151_n_0),
        .I1(fdatx[9]),
        .I2(fch_issu1_inferred_i_152_n_0),
        .I3(fdatx[4]),
        .I4(fch_issu1_inferred_i_107_n_0),
        .I5(fch_issu1_inferred_i_88_n_0),
        .O(fch_issu1_inferred_i_84_n_0));
  LUT6 #(
    .INIT(64'h57555555FFFF00FF)) 
    fch_issu1_inferred_i_85
       (.I0(fch_issu1_inferred_i_153_n_0),
        .I1(fch_issu1_inferred_i_154_n_0),
        .I2(fch_issu1_inferred_i_155_n_0),
        .I3(fch_issu1_inferred_i_97_n_0),
        .I4(fdatx[8]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_85_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_86
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .O(fch_issu1_inferred_i_86_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_87
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_87_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    fch_issu1_inferred_i_88
       (.I0(fch_issu1_inferred_i_156_n_0),
        .I1(fdatx[15]),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .I5(fch_issu1_inferred_i_157_n_0),
        .O(fch_issu1_inferred_i_88_n_0));
  LUT6 #(
    .INIT(64'hFF1AFAF0FFFFFFFF)) 
    fch_issu1_inferred_i_89
       (.I0(fdat[8]),
        .I1(\nir_id[18]_i_8_n_0 ),
        .I2(fdat[11]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat_12_sn_1),
        .O(fch_issu1_inferred_i_89_n_0));
  LUT6 #(
    .INIT(64'h04C0C0C800000000)) 
    fch_issu1_inferred_i_90
       (.I0(fdat[0]),
        .I1(fch_issu1_inferred_i_158_n_0),
        .I2(fdat[2]),
        .I3(fdat[3]),
        .I4(fdat[1]),
        .I5(\nir_id[14]_i_8_n_0 ),
        .O(fch_issu1_inferred_i_90_n_0));
  LUT4 #(
    .INIT(16'h0440)) 
    fch_issu1_inferred_i_91
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .I2(fdatx[12]),
        .I3(fdatx[11]),
        .O(fch_issu1_inferred_i_91_n_0));
  LUT6 #(
    .INIT(64'hFFFF1DDDFFFFFFFF)) 
    fch_issu1_inferred_i_92
       (.I0(fch_issu1_inferred_i_159_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[9]),
        .I3(fdatx[7]),
        .I4(fch_issu1_inferred_i_160_n_0),
        .I5(fch_issu1_inferred_i_161_n_0),
        .O(fch_issu1_inferred_i_92_n_0));
  LUT6 #(
    .INIT(64'h00000000830303C3)) 
    fch_issu1_inferred_i_93
       (.I0(fdatx[3]),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_154_n_0),
        .I4(fdatx[6]),
        .I5(fch_issu1_inferred_i_162_n_0),
        .O(fch_issu1_inferred_i_93_n_0));
  LUT6 #(
    .INIT(64'hFFFAFFFF1FA0FFFF)) 
    fch_issu1_inferred_i_94
       (.I0(fdatx[8]),
        .I1(fch_issu1_inferred_i_97_n_0),
        .I2(fdatx[10]),
        .I3(fdatx[11]),
        .I4(fch_issu1_inferred_i_163_n_0),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_94_n_0));
  LUT6 #(
    .INIT(64'hFEEEFEEEFFFEEFFF)) 
    fch_issu1_inferred_i_95
       (.I0(fch_issu1_inferred_i_164_n_0),
        .I1(fch_issu1_inferred_i_165_n_0),
        .I2(fdatx[3]),
        .I3(fdatx[1]),
        .I4(fdatx[0]),
        .I5(fdatx[2]),
        .O(fch_issu1_inferred_i_95_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    fch_issu1_inferred_i_96
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[15]),
        .I4(fadr_1_fl),
        .O(fch_issu1_inferred_i_96_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_97
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .O(fch_issu1_inferred_i_97_n_0));
  LUT6 #(
    .INIT(64'h5000500050005004)) 
    fch_issu1_inferred_i_99
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_49_0),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .I5(fch_issu1_inferred_i_167_n_0),
        .O(fch_issu1_inferred_i_99_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry
       (.CI(\<const0> ),
        .CO({fch_pc_nx2_carry_n_0,fch_pc_nx2_carry_n_1,fch_pc_nx2_carry_n_2,fch_pc_nx2_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\pc0_reg[15]_1 [1],\<const0> }),
        .O(p_2_in_0[3:0]),
        .S({\pc0_reg[15]_1 [3:2],\fadr[3] ,\pc0_reg[15]_1 [0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry__0
       (.CI(fch_pc_nx2_carry_n_0),
        .CO({fch_pc_nx2_carry__0_n_0,fch_pc_nx2_carry__0_n_1,fch_pc_nx2_carry__0_n_2,fch_pc_nx2_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(p_2_in_0[7:4]),
        .S(\pc0_reg[15]_1 [7:4]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry__1
       (.CI(fch_pc_nx2_carry__0_n_0),
        .CO({fch_pc_nx2_carry__1_n_0,fch_pc_nx2_carry__1_n_1,fch_pc_nx2_carry__1_n_2,fch_pc_nx2_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(p_2_in_0[11:8]),
        .S(\pc0_reg[15]_1 [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx2_carry__2
       (.CI(fch_pc_nx2_carry__1_n_0),
        .CO({fch_pc_nx2_carry__2_n_1,fch_pc_nx2_carry__2_n_2,fch_pc_nx2_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\pc_reg[15] ,p_2_in_0[12]}),
        .S(\pc0_reg[15]_1 [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry
       (.CI(\<const0> ),
        .CO({fch_pc_nx4_carry_n_0,fch_pc_nx4_carry_n_1,fch_pc_nx4_carry_n_2,fch_pc_nx4_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\pc0_reg[15]_1 [2],\<const0> }),
        .O({fch_pc_nx4_carry_n_4,fch_pc_nx4_carry_n_5,fch_pc_nx4_carry_n_6,fch_pc_nx4_carry_n_7}),
        .S({\pc0_reg[15]_1 [4:3],S,\pc0_reg[15]_1 [1]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry__0
       (.CI(fch_pc_nx4_carry_n_0),
        .CO({fch_pc_nx4_carry__0_n_0,fch_pc_nx4_carry__0_n_1,fch_pc_nx4_carry__0_n_2,fch_pc_nx4_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({fch_pc_nx4_carry__0_n_4,fch_pc_nx4_carry__0_n_5,fch_pc_nx4_carry__0_n_6,fch_pc_nx4_carry__0_n_7}),
        .S(\pc0_reg[15]_1 [8:5]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry__1
       (.CI(fch_pc_nx4_carry__0_n_0),
        .CO({fch_pc_nx4_carry__1_n_0,fch_pc_nx4_carry__1_n_1,fch_pc_nx4_carry__1_n_2,fch_pc_nx4_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({fch_pc_nx4_carry__1_n_4,fch_pc_nx4_carry__1_n_5,fch_pc_nx4_carry__1_n_6,fch_pc_nx4_carry__1_n_7}),
        .S(\pc0_reg[15]_1 [12:9]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 fch_pc_nx4_carry__2
       (.CI(fch_pc_nx4_carry__1_n_0),
        .CO({fch_pc_nx4_carry__2_n_2,fch_pc_nx4_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(O),
        .S({\<const0> ,\pc0_reg[15]_1 [15:13]}));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(fch_term_fl),
        .R(\<const0> ));
  mcss_fch_fsm fctl
       (.D(fch_pc),
        .E(fch_nir_lir),
        .O({fch_pc_nx4_carry_n_4,fch_pc_nx4_carry_n_5,fch_pc_nx4_carry_n_6,fch_pc_nx4_carry_n_7}),
        .Q(Q),
        .S({fctl_n_85,fctl_n_86,fctl_n_87,fctl_n_88}),
        .alu_sr_flag0({alu_sr_flag0[3],alu_sr_flag0[0]}),
        .alu_sr_flag1(alu_sr_flag1),
        .brdy(brdy),
        .brdy_0(fch_term),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .crdy_0(fctl_n_91),
        .ctl_fetch0(ctl_fetch0),
        .ctl_fetch0_fl(ctl_fetch0_fl),
        .ctl_fetch0_fl_i_15_0(\stat[2]_i_12_n_0 ),
        .ctl_fetch0_fl_i_16_0(ctl_fetch0_fl_i_16),
        .ctl_fetch0_fl_i_16_1(ctl_fetch0_fl_i_16_0),
        .ctl_fetch0_fl_i_27_0(\ccmd[4]_INST_0_i_15_n_0 ),
        .ctl_fetch0_fl_i_2_0(\stat[0]_i_22_n_0 ),
        .ctl_fetch0_fl_i_4_0(\rgf_selc0_wb[1]_i_6_n_0 ),
        .ctl_fetch0_fl_i_4_1(\bdatw[10]_INST_0_i_18_n_0 ),
        .ctl_fetch0_fl_i_8_0(ctl_fetch0_fl_i_8),
        .ctl_fetch0_fl_reg(ir0),
        .ctl_fetch0_fl_reg_0(\rgf_selc0_rn_wb_reg[0] ),
        .ctl_fetch0_fl_reg_1(ctl_fetch0_fl_reg_1),
        .ctl_fetch0_fl_reg_2(ctl_fetch0_fl_reg_2),
        .ctl_fetch0_fl_reg_3(ctl_fetch0_fl_reg_0),
        .ctl_fetch0_fl_reg_4(rst_n_fl_reg_2),
        .ctl_fetch0_fl_reg_5(\bcmd[2]_INST_0_i_9_n_0 ),
        .ctl_fetch1(ctl_fetch1),
        .ctl_fetch1_fl(ctl_fetch1_fl),
        .ctl_fetch1_fl_i_16_0(ctl_fetch1_fl_i_16),
        .ctl_fetch1_fl_i_21_0(ir1),
        .ctl_fetch1_fl_i_25_0(\stat[0]_i_8__1_n_0 ),
        .ctl_fetch1_fl_i_25_1(ctl_fetch1_fl_i_36_n_0),
        .ctl_fetch1_fl_i_27_0(\bdatw[15]_INST_0_i_252_n_0 ),
        .ctl_fetch1_fl_i_27_1(\stat[0]_i_19__0_n_0 ),
        .ctl_fetch1_fl_i_27_2(\stat[2]_i_10__0_n_0 ),
        .ctl_fetch1_fl_i_2_0(\bcmd[0]_INST_0_i_3_n_0 ),
        .ctl_fetch1_fl_i_2_1(\badrx[15]_INST_0_i_5_n_0 ),
        .ctl_fetch1_fl_i_2_2(tout__1_carry_i_22_0),
        .ctl_fetch1_fl_i_2_3(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .ctl_fetch1_fl_i_2_4(rst_n_fl_reg_9),
        .ctl_fetch1_fl_i_2_5(ctl_fetch1_fl_i_20_n_0),
        .ctl_fetch1_fl_i_2_6(\bcmd[1]_0 ),
        .ctl_fetch1_fl_i_34_0(\stat[0]_i_30__0_n_0 ),
        .ctl_fetch1_fl_reg(\rgf_selc1_wb_reg[1] ),
        .ctl_fetch1_fl_reg_0(\bcmd[2]_INST_0_i_7_n_0 ),
        .ctl_fetch1_fl_reg_1(\bcmd[2]_INST_0_i_5_n_0 ),
        .ctl_fetch1_fl_reg_i_6_0(\stat[0]_i_2__1_0 ),
        .ctl_fetch1_fl_reg_i_6_1(\bbus_o[4]_INST_0_i_49_0 ),
        .ctl_fetch1_fl_reg_i_6_2(ctl_fetch1_fl_reg_i_6),
        .ctl_fetch_ext_fl(ctl_fetch_ext_fl),
        .ctl_sr_ldie0(ctl_sr_ldie0),
        .ctl_sr_ldie1(ctl_sr_ldie1),
        .ctl_sr_upd0(ctl_sr_upd0),
        .ctl_sr_upd1(ctl_sr_upd1),
        .eir(eir),
        .\eir_fl_reg[15] (nir),
        .\eir_fl_reg[15]_0 ({\eir_fl_reg_n_0_[15] ,\eir_fl_reg_n_0_[14] ,\eir_fl_reg_n_0_[13] ,\eir_fl_reg_n_0_[12] ,\eir_fl_reg_n_0_[11] ,\eir_fl_reg_n_0_[10] ,\eir_fl_reg_n_0_[9] ,\eir_fl_reg_n_0_[8] ,\eir_fl_reg_n_0_[7] ,\eir_fl_reg_n_0_[6] ,\eir_fl_reg_n_0_[5] ,\eir_fl_reg_n_0_[4] ,\eir_fl_reg_n_0_[3] ,\eir_fl_reg_n_0_[2] ,\eir_fl_reg_n_0_[1] ,\eir_fl_reg_n_0_[0] }),
        .fadr(fadr),
        .\fadr[12] ({fch_pc_nx4_carry__1_n_4,fch_pc_nx4_carry__1_n_5,fch_pc_nx4_carry__1_n_6,fch_pc_nx4_carry__1_n_7}),
        .\fadr[8] ({fch_pc_nx4_carry__0_n_4,fch_pc_nx4_carry__0_n_5,fch_pc_nx4_carry__0_n_6,fch_pc_nx4_carry__0_n_7}),
        .fadr_1_fl(fadr_1_fl),
        .fch_irq_lev(fch_irq_lev),
        .\fch_irq_lev[1]_i_2 (\fadr[15]_INST_0_i_16_n_0 ),
        .\fch_irq_lev[1]_i_2_0 (\rgf_c1bus_wb[14]_i_53_0 ),
        .fch_irq_req(fch_irq_req),
        .fch_irq_req_fl_reg(fch_irq_req_fl_reg_0),
        .fch_issu1(fch_issu1),
        .fch_issu1_fl(fch_issu1_fl),
        .fch_issu1_inferred_i_11_0({nir_id[24],nir_id[21:12]}),
        .fch_issu1_inferred_i_11_1(fch_issu1_inferred_i_94_n_0),
        .fch_issu1_inferred_i_11_2(fch_issu1_inferred_i_95_n_0),
        .fch_issu1_inferred_i_11_3(fch_issu1_inferred_i_89_n_0),
        .fch_issu1_inferred_i_11_4(fch_issu1_inferred_i_90_n_0),
        .fch_issu1_inferred_i_11_5(fch_issu1_inferred_i_91_n_0),
        .fch_issu1_inferred_i_1_0(fch_issu1_inferred_i_25_n_0),
        .fch_issu1_inferred_i_1_1(fch_issu1_inferred_i_26_n_0),
        .fch_issu1_inferred_i_1_2(fch_issu1_inferred_i_27_n_0),
        .fch_issu1_inferred_i_1_3(fch_issu1_inferred_i_14_n_0),
        .fch_issu1_inferred_i_1_4(fch_issu1_inferred_i_15_n_0),
        .fch_issu1_inferred_i_1_5(fch_issu1_inferred_i_16_n_0),
        .fch_issu1_inferred_i_1_6(fch_issu1_inferred_i_17_n_0),
        .fch_issu1_inferred_i_20_0(fch_issu1_inferred_i_102_n_0),
        .fch_issu1_inferred_i_20_1(fch_issu1_inferred_i_103_n_0),
        .fch_issu1_inferred_i_20_2(fch_issu1_inferred_i_99_n_0),
        .fch_issu1_inferred_i_28_0(\nir_id[16]_i_3_n_0 ),
        .fch_issu1_inferred_i_28_1(fch_issu1_inferred_i_109_n_0),
        .fch_issu1_inferred_i_28_2(fch_issu1_inferred_i_110_n_0),
        .fch_issu1_inferred_i_28_3(fch_issu1_inferred_i_111_n_0),
        .fch_issu1_inferred_i_2_0(fch_issu1_inferred_i_39_n_0),
        .fch_issu1_inferred_i_2_1(fch_issu1_inferred_i_36_n_0),
        .fch_issu1_inferred_i_2_2(fch_issu1_inferred_i_37_n_0),
        .fch_issu1_inferred_i_31_0(fch_issu1_inferred_i_126_n_0),
        .fch_issu1_inferred_i_32_0(fch_issu1_inferred_i_145_n_0),
        .fch_issu1_inferred_i_32_1(fch_issu1_inferred_i_146_n_0),
        .fch_issu1_inferred_i_32_2(fch_issu1_inferred_i_147_n_0),
        .fch_issu1_inferred_i_33_0(fch_issu1_inferred_i_148_n_0),
        .fch_issu1_inferred_i_33_1(fch_issu1_inferred_i_88_n_0),
        .fch_issu1_inferred_i_33_2(fch_issu1_inferred_i_149_n_0),
        .fch_issu1_inferred_i_33_3(fdatx_14_sn_1),
        .fch_issu1_inferred_i_41_0(fch_issu1_inferred_i_83_n_0),
        .fch_issu1_inferred_i_41_1(fch_issu1_inferred_i_84_n_0),
        .fch_issu1_inferred_i_41_2(fch_issu1_inferred_i_81_n_0),
        .fch_issu1_inferred_i_41_3(fch_issu1_inferred_i_82_n_0),
        .fch_issu1_inferred_i_5_0(fch_issu1_inferred_i_45_n_0),
        .fch_issu1_inferred_i_5_1(fch_issu1_inferred_i_43_n_0),
        .fch_issu1_inferred_i_6_0(fch_issu1_inferred_i_47_n_0),
        .fch_issu1_inferred_i_6_1(fch_issu1_inferred_i_52_n_0),
        .fch_issu1_inferred_i_6_2(fch_issu1_inferred_i_53_n_0),
        .fch_issu1_inferred_i_6_3(fch_issu1_inferred_i_54_n_0),
        .fch_issu1_inferred_i_6_4(fch_issu1_inferred_i_55_n_0),
        .fch_issu1_inferred_i_7_0(fch_issu1_inferred_i_62_n_0),
        .fch_issu1_inferred_i_7_1(fch_issu1_inferred_i_63_n_0),
        .fch_issu1_inferred_i_7_2(fch_issu1_inferred_i_64_n_0),
        .fch_issu1_inferred_i_7_3(fch_issu1_inferred_i_65_n_0),
        .fch_issu1_inferred_i_7_4(fch_issu1_inferred_i_66_n_0),
        .fch_issu1_inferred_i_7_5(fch_issu1_inferred_i_67_n_0),
        .fch_issu1_inferred_i_7_6(fch_issu1_inferred_i_69_n_0),
        .fch_issu1_inferred_i_8_0(\nir_id[12]_i_2_n_0 ),
        .fch_issu1_inferred_i_8_1(fch_issu1_inferred_i_49_n_0),
        .fch_issu1_inferred_i_8_10(fch_issu1_inferred_i_51_n_0),
        .fch_issu1_inferred_i_8_2(\nir_id[14]_i_2_n_0 ),
        .fch_issu1_inferred_i_8_3(fch_issu1_inferred_i_71_n_0),
        .fch_issu1_inferred_i_8_4(fch_issu1_inferred_i_72_n_0),
        .fch_issu1_inferred_i_8_5(fch_issu1_inferred_i_73_n_0),
        .fch_issu1_inferred_i_8_6(fch_issu1_inferred_i_76_n_0),
        .fch_issu1_inferred_i_8_7(fch_issu1_inferred_i_77_n_0),
        .fch_issu1_inferred_i_8_8(fch_issu1_inferred_i_78_n_0),
        .fch_issu1_inferred_i_8_9(\nir_id[13]_i_2_n_0 ),
        .fch_issu1_ir(fch_issu1_ir),
        .fch_leir_lir_reg_0(\fadr[15]_INST_0_i_11_n_0 ),
        .fch_leir_lir_reg_1(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .fch_leir_nir_reg_0(\stat[2]_i_5__1_n_0 ),
        .fch_leir_nir_reg_1(\stat[2]_i_14_n_0 ),
        .fch_memacc1(fch_memacc1),
        .fch_term_fl(fch_term_fl),
        .fch_wrbufn1(fch_wrbufn1),
        .fdat(fdat),
        .fdatx(fdatx),
        .\grn[15]_i_3__5_0 (\stat_reg[2]_0 ),
        .\grn[15]_i_3__5_1 (\grn[15]_i_3__5 ),
        .\grn_reg[15] (\grn_reg[15] ),
        .\grn_reg[15]_0 (\stat_reg[2] ),
        .\grn_reg[15]_1 (\grn_reg[15]_0 ),
        .in0(ir0),
        .\ir0_fl_reg[0] (fch_irq_req_fl),
        .\ir0_fl_reg[15] (ir0_fl),
        .\ir0_id_fl_reg[20] (\ir0_id_fl[21]_i_4_n_0 ),
        .\ir0_id_fl_reg[21] (ir0_id_fl),
        .ir1(ir1),
        .\ir1_fl_reg[0] (ir1_inferred_i_17_n_0),
        .\ir1_fl_reg[15] (ir1_fl),
        .\ir1_id_fl_reg[20] (\ir1_id_fl_reg[20]_0 ),
        .\ir1_id_fl_reg[21] (ir1_id_fl),
        .\ir1_id_fl_reg[21]_0 ({\nir_id_reg[21]_0 ,lir_id_0[19:16]}),
        .\ir1_id_fl_reg[21]_1 (\ir1_id_fl_reg[21]_0 ),
        .\iv_reg[15] (\iv_reg[15] ),
        .\iv_reg[15]_0 (\iv_reg[15]_0 ),
        .out(fch_issu1),
        .p_2_in(p_2_in),
        .p_2_in_0(p_2_in_0),
        .\pc0_reg[12] (\pc0_reg[15]_1 [12:0]),
        .\pc0_reg[3] (\stat_reg[0] ),
        .\pc_reg[0] (\stat[2]_i_4 ),
        .\pc_reg[11] ({fctl_n_154,fctl_n_155,fctl_n_156,fctl_n_157}),
        .\pc_reg[12] (fctl_n_158),
        .\pc_reg[13] (\pc_reg[13] ),
        .\pc_reg[14] (\pc[14]_i_5_n_0 ),
        .\pc_reg[14]_0 (\rgf_c0bus_wb[14]_i_2_n_0 ),
        .\pc_reg[14]_1 (\pc_reg[14] ),
        .\pc_reg[15] (\bdatr[15] ),
        .\pc_reg[15]_0 ({\cbus_i[15] [15],\cbus_i[15] [13:4],\cbus_i[15] [2:0]}),
        .\pc_reg[15]_1 (\pc_reg[15]_0 ),
        .\pc_reg[15]_2 (\pc_reg[15]_1 ),
        .\pc_reg[7] ({fctl_n_150,fctl_n_151,fctl_n_152,fctl_n_153}),
        .rgf_selc0_stat(rgf_selc0_stat),
        .rgf_selc1_stat(rgf_selc1_stat),
        .rgf_selc1_stat_reg(rgf_selc1_stat_reg),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat_reg_0),
        .rgf_selc1_stat_reg_1(rgf_selc1_stat_reg_1),
        .rgf_selc1_stat_reg_10(rgf_selc1_stat_reg_10),
        .rgf_selc1_stat_reg_11(rgf_selc1_stat_reg_11),
        .rgf_selc1_stat_reg_12(rgf_selc1_stat_reg_12),
        .rgf_selc1_stat_reg_13(rgf_selc1_stat_reg_13),
        .rgf_selc1_stat_reg_14(rgf_selc1_stat_reg_14),
        .rgf_selc1_stat_reg_15(rgf_selc1_stat_reg_15),
        .rgf_selc1_stat_reg_16(rgf_selc1_stat_reg_16),
        .rgf_selc1_stat_reg_17(rgf_selc1_stat_reg_17),
        .rgf_selc1_stat_reg_18(rgf_selc1_stat_reg_18),
        .rgf_selc1_stat_reg_19(rgf_selc1_stat_reg_19),
        .rgf_selc1_stat_reg_2(rgf_selc1_stat_reg_2),
        .rgf_selc1_stat_reg_20(rgf_selc1_stat_reg_20),
        .rgf_selc1_stat_reg_21(rgf_selc1_stat_reg_21),
        .rgf_selc1_stat_reg_22(rgf_selc1_stat_reg_22),
        .rgf_selc1_stat_reg_23(rgf_selc1_stat_reg_23),
        .rgf_selc1_stat_reg_24(rgf_selc1_stat_reg_24),
        .rgf_selc1_stat_reg_25(rgf_selc1_stat_reg_25),
        .rgf_selc1_stat_reg_26(rgf_selc1_stat_reg_26),
        .rgf_selc1_stat_reg_27(rgf_selc1_stat_reg_27),
        .rgf_selc1_stat_reg_28(rgf_selc1_stat_reg_28),
        .rgf_selc1_stat_reg_29(rgf_selc1_stat_reg_29),
        .rgf_selc1_stat_reg_3(rgf_selc1_stat_reg_3),
        .rgf_selc1_stat_reg_30(rgf_selc1_stat_reg_30),
        .rgf_selc1_stat_reg_31(rgf_selc1_stat_reg_31),
        .rgf_selc1_stat_reg_4(rgf_selc1_stat_reg_4),
        .rgf_selc1_stat_reg_5(rgf_selc1_stat_reg_5),
        .rgf_selc1_stat_reg_6(rgf_selc1_stat_reg_6),
        .rgf_selc1_stat_reg_7(rgf_selc1_stat_reg_7),
        .rgf_selc1_stat_reg_8(rgf_selc1_stat_reg_8),
        .rgf_selc1_stat_reg_9(rgf_selc1_stat_reg_9),
        .rst_n(rst_n),
        .rst_n_0(rst_n_0),
        .rst_n_fl(rst_n_fl),
        .rst_n_fl_reg(rst_n_fl_reg_1),
        .rst_n_fl_reg_0(fctl_n_89),
        .rst_n_fl_reg_1(fctl_n_95),
        .rst_n_fl_reg_2(fctl_n_96),
        .rst_n_fl_reg_3({ir0_id,p_0_in_1}),
        .rst_n_fl_reg_4(fctl_n_133),
        .\sp_reg[0] (\sp[0]_i_2_n_0 ),
        .\sp_reg[10] (\sp_reg[10] ),
        .\sp_reg[11] (\sp_reg[11] ),
        .\sp_reg[12] (\sp_reg[12] ),
        .\sp_reg[13] (\sp_reg[13] ),
        .\sp_reg[14] (\sp_reg[14] ),
        .\sp_reg[15] (\sp_reg[15] ),
        .\sp_reg[15]_0 (\sp_reg[15]_0 ),
        .\sp_reg[1] (\sp_reg[1] ),
        .\sp_reg[2] (\sp_reg[2] ),
        .\sp_reg[3] (\sp_reg[3] ),
        .\sp_reg[4] (\sp_reg[4] ),
        .\sp_reg[5] (\sp_reg[5] ),
        .\sp_reg[6] (\sp_reg[6] ),
        .\sp_reg[7] (\sp_reg[7] ),
        .\sp_reg[8] (\sp_reg[8] ),
        .\sp_reg[9] (\sp_reg[9] ),
        .\sr[13]_i_13 (\ccmd[4]_INST_0_i_12_n_0 ),
        .\sr[13]_i_5_0 (\stat_reg[2]_1 ),
        .\sr[13]_i_5_1 (\sr[13]_i_5 ),
        .\sr[13]_i_5_2 (\stat_reg[2]_2 ),
        .\sr[13]_i_5_3 (\sr[13]_i_5_0 ),
        .\sr_reg[0] (\sr_reg[0]_36 ),
        .\sr_reg[0]_0 (\sr_reg[0]_37 ),
        .\sr_reg[0]_1 (\sr_reg[0]_38 ),
        .\sr_reg[0]_10 (\sr_reg[0]_47 ),
        .\sr_reg[0]_11 (\sr_reg[0]_48 ),
        .\sr_reg[0]_12 (\sr_reg[0]_49 ),
        .\sr_reg[0]_13 (\sr_reg[0]_50 ),
        .\sr_reg[0]_14 (\sr_reg[0]_51 ),
        .\sr_reg[0]_15 (\sr_reg[0]_52 ),
        .\sr_reg[0]_16 (\sr_reg[0]_53 ),
        .\sr_reg[0]_17 (\sr_reg[0]_54 ),
        .\sr_reg[0]_18 (\sr_reg[0]_55 ),
        .\sr_reg[0]_19 (\sr_reg[0]_56 ),
        .\sr_reg[0]_2 (\sr_reg[0]_39 ),
        .\sr_reg[0]_20 (\sr_reg[0]_57 ),
        .\sr_reg[0]_21 (\sr_reg[0]_58 ),
        .\sr_reg[0]_22 (\sr_reg[0]_59 ),
        .\sr_reg[0]_3 (\sr_reg[0]_40 ),
        .\sr_reg[0]_4 (\sr_reg[0]_41 ),
        .\sr_reg[0]_5 (\sr_reg[0]_42 ),
        .\sr_reg[0]_6 (\sr_reg[0]_43 ),
        .\sr_reg[0]_7 (\sr_reg[0]_44 ),
        .\sr_reg[0]_8 (\sr_reg[0]_45 ),
        .\sr_reg[0]_9 (\sr_reg[0]_46 ),
        .\sr_reg[15] (\sr_reg[15] ),
        .\sr_reg[15]_0 (\sr_reg[15]_0 ),
        .\sr_reg[1] (\sr_reg[1]_14 ),
        .\sr_reg[1]_0 (\sr_reg[1]_15 ),
        .\sr_reg[1]_1 (\sr_reg[1]_16 ),
        .\sr_reg[1]_2 (\sr_reg[1]_17 ),
        .\sr_reg[1]_3 (\sr_reg[1]_18 ),
        .\sr_reg[1]_4 (\sr_reg[1]_19 ),
        .\sr_reg[1]_5 (\sr_reg[1]_20 ),
        .\sr_reg[1]_6 (\sr_reg[1]_21 ),
        .\sr_reg[3] (\sr[3]_i_7_n_0 ),
        .\sr_reg[3]_0 (\rgf_c0bus_wb[3]_i_2_n_0 ),
        .\sr_reg[4] (\sr_reg[4]_1 ),
        .\sr_reg[5] (\sr_reg[5]_0 ),
        .\sr_reg[5]_0 (\sr[6]_i_6_n_0 ),
        .\sr_reg[5]_1 (\rgf_c1bus_wb[15]_i_4_n_0 ),
        .\sr_reg[5]_2 (\rgf_c1bus_wb[15]_i_5_n_0 ),
        .\sr_reg[5]_3 (\sr[5]_i_7_n_0 ),
        .\sr_reg[5]_4 (\sr[5]_i_8_n_0 ),
        .\sr_reg[5]_5 (\sr[6]_i_7_n_0 ),
        .\sr_reg[5]_6 (\rgf_c0bus_wb[15]_i_4_n_0 ),
        .\sr_reg[5]_7 (\tr_reg[4] ),
        .\sr_reg[5]_8 (\sr[5]_i_9_n_0 ),
        .\sr_reg[5]_9 (\sr[5]_i_10_n_0 ),
        .\sr_reg[6] (\stat_reg[2]_3 ),
        .\sr_reg[6]_0 (\sr_reg[6]_1 ),
        .\sr_reg[6]_1 (\sr[6]_i_8_n_0 ),
        .\sr_reg[7] (tout__1_carry_i_11_0),
        .\sr_reg[7]_0 (\rgf_c1bus_wb[15]_i_3_n_0 ),
        .\sr_reg[7]_1 (\rgf_c1bus_wb_reg[15] [1]),
        .\stat[2]_i_4_0 (\stat[2]_i_9_n_0 ),
        .\stat[2]_i_4_1 (\fadr[15]_INST_0_i_13_n_0 ),
        .\stat[2]_i_4_2 (\fch_irq_lev[1]_i_2_0 ),
        .\stat_reg[0]_0 (\stat_reg[0]_5 ),
        .\stat_reg[0]_1 (\stat_reg[0]_15 ),
        .\stat_reg[0]_2 (\stat_reg[0]_51 ),
        .\stat_reg[0]_3 (\stat_reg[0]_48 ),
        .\stat_reg[0]_4 (\stat[0]_i_2__0_n_0 ),
        .\stat_reg[0]_5 (\stat[0]_i_3__2_n_0 ),
        .\stat_reg[0]_6 (\stat[0]_i_4_n_0 ),
        .\stat_reg[0]_7 (\stat[0]_i_5_n_0 ),
        .\stat_reg[0]_8 (\stat_reg[0]_56 ),
        .\stat_reg[1]_0 (\stat_reg[1] ),
        .\stat_reg[1]_1 (\stat_reg[1]_3 ),
        .\stat_reg[1]_2 (fctl_n_94),
        .\stat_reg[2]_0 (fctl_n_67),
        .\tr_reg[15] (\tr_reg[15]_0 ),
        .\tr_reg[15]_0 (\tr_reg[15]_1 ));
  FDRE \ir0_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[0]),
        .Q(ir0_fl[0]),
        .R(SR));
  FDRE \ir0_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[10]),
        .Q(ir0_fl[10]),
        .R(SR));
  FDRE \ir0_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[11]),
        .Q(ir0_fl[11]),
        .R(SR));
  FDRE \ir0_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[12]),
        .Q(ir0_fl[12]),
        .R(SR));
  FDRE \ir0_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[13]),
        .Q(ir0_fl[13]),
        .R(SR));
  FDRE \ir0_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[14]),
        .Q(ir0_fl[14]),
        .R(SR));
  FDRE \ir0_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[15]),
        .Q(ir0_fl[15]),
        .R(SR));
  FDRE \ir0_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[1]),
        .Q(ir0_fl[1]),
        .R(SR));
  FDRE \ir0_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[2]),
        .Q(ir0_fl[2]),
        .R(SR));
  FDRE \ir0_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[3]),
        .Q(ir0_fl[3]),
        .R(SR));
  FDRE \ir0_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[4]),
        .Q(ir0_fl[4]),
        .R(SR));
  FDRE \ir0_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[5]),
        .Q(ir0_fl[5]),
        .R(SR));
  FDRE \ir0_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[6]),
        .Q(ir0_fl[6]),
        .R(SR));
  FDRE \ir0_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[7]),
        .Q(ir0_fl[7]),
        .R(SR));
  FDRE \ir0_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[8]),
        .Q(ir0_fl[8]),
        .R(SR));
  FDRE \ir0_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0[9]),
        .Q(ir0_fl[9]),
        .R(SR));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[20]_i_8 
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(fdatx_5_sn_1));
  LUT2 #(
    .INIT(4'hB)) 
    \ir0_id_fl[21]_i_4 
       (.I0(fch_irq_req_fl),
        .I1(fch_term_fl),
        .O(\ir0_id_fl[21]_i_4_n_0 ));
  FDRE \ir0_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_0_in_1),
        .Q(ir0_id_fl[20]),
        .R(SR));
  FDRE \ir0_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir0_id),
        .Q(ir0_id_fl[21]),
        .R(SR));
  FDRE \ir1_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[0]),
        .Q(ir1_fl[0]),
        .R(SR));
  FDRE \ir1_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[10]),
        .Q(ir1_fl[10]),
        .R(SR));
  FDRE \ir1_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[11]),
        .Q(ir1_fl[11]),
        .R(SR));
  FDRE \ir1_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[12]),
        .Q(ir1_fl[12]),
        .R(SR));
  FDRE \ir1_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[13]),
        .Q(ir1_fl[13]),
        .R(SR));
  FDRE \ir1_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[14]),
        .Q(ir1_fl[14]),
        .R(SR));
  FDRE \ir1_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[15]),
        .Q(ir1_fl[15]),
        .R(SR));
  FDRE \ir1_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[1]),
        .Q(ir1_fl[1]),
        .R(SR));
  FDRE \ir1_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[2]),
        .Q(ir1_fl[2]),
        .R(SR));
  FDRE \ir1_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[3]),
        .Q(ir1_fl[3]),
        .R(SR));
  FDRE \ir1_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[4]),
        .Q(ir1_fl[4]),
        .R(SR));
  FDRE \ir1_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[5]),
        .Q(ir1_fl[5]),
        .R(SR));
  FDRE \ir1_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[6]),
        .Q(ir1_fl[6]),
        .R(SR));
  FDRE \ir1_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[7]),
        .Q(ir1_fl[7]),
        .R(SR));
  FDRE \ir1_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[8]),
        .Q(ir1_fl[8]),
        .R(SR));
  FDRE \ir1_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir1[9]),
        .Q(ir1_fl[9]),
        .R(SR));
  FDRE \ir1_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_wrbufn1),
        .Q(ir1_id_fl[20]),
        .R(SR));
  FDRE \ir1_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_memacc1),
        .Q(ir1_id_fl[21]),
        .R(SR));
  LUT3 #(
    .INIT(8'h08)) 
    ir1_inferred_i_17
       (.I0(fch_issu1),
        .I1(fch_term_fl),
        .I2(fch_irq_req_fl),
        .O(ir1_inferred_i_17_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[12]_i_1 
       (.I0(\nir_id[12]_i_2_n_0 ),
        .O(lir_id_0[12]));
  LUT5 #(
    .INIT(32'h55551011)) 
    \nir_id[12]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[14]_i_4_n_0 ),
        .I2(\nir_id[12]_i_3_n_0 ),
        .I3(\nir_id[12]_i_4_n_0 ),
        .I4(fdat[15]),
        .O(\nir_id[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h45550505FFFFFFFF)) 
    \nir_id[12]_i_3 
       (.I0(\nir_id[14]_i_10_n_0 ),
        .I1(fdat[8]),
        .I2(fdat[10]),
        .I3(fdat[0]),
        .I4(\nir_id[14]_i_9_n_0 ),
        .I5(fdat[14]),
        .O(\nir_id[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hBAAAAAAA)) 
    \nir_id[12]_i_4 
       (.I0(\nir_id[14]_i_11_n_0 ),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(fdat[10]),
        .I4(fdat[0]),
        .O(\nir_id[12]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[13]_i_1 
       (.I0(\nir_id[13]_i_2_n_0 ),
        .O(lir_id_0[13]));
  LUT6 #(
    .INIT(64'h558F558F0000F000)) 
    \nir_id[13]_i_2 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(\nir_id[13]_i_3_n_0 ),
        .I5(fdat[15]),
        .O(\nir_id[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF08AA)) 
    \nir_id[13]_i_3 
       (.I0(fdat[10]),
        .I1(fdat[1]),
        .I2(fdat[8]),
        .I3(\nir_id[14]_i_9_n_0 ),
        .I4(\nir_id[14]_i_10_n_0 ),
        .I5(\nir_id[13]_i_4_n_0 ),
        .O(\nir_id[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h83B3BFBF00000000)) 
    \nir_id[13]_i_4 
       (.I0(\nir_id[13]_i_5_n_0 ),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[1]),
        .I4(fdat[8]),
        .I5(\nir_id[13]_i_6_n_0 ),
        .O(\nir_id[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0C400C000C00C00C)) 
    \nir_id[13]_i_5 
       (.I0(fdat[3]),
        .I1(fdat[8]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[6]),
        .I5(fdat[4]),
        .O(\nir_id[13]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[13]_i_6 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .O(\nir_id[13]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[14]_i_1 
       (.I0(\nir_id[14]_i_2_n_0 ),
        .O(lir_id_0[14]));
  LUT5 #(
    .INIT(32'hF3F7F3FF)) 
    \nir_id[14]_i_10 
       (.I0(\nir_id[14]_i_12_n_0 ),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .O(\nir_id[14]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h77FFF7F777777777)) 
    \nir_id[14]_i_11 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[8]),
        .I3(\nir_id[14]_i_13_n_0 ),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(\nir_id[14]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \nir_id[14]_i_12 
       (.I0(fdat[6]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .O(\nir_id[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAA0A2000AAA8000A)) 
    \nir_id[14]_i_13 
       (.I0(fdat[8]),
        .I1(fdat[3]),
        .I2(fdat[4]),
        .I3(fdat[6]),
        .I4(fdat[7]),
        .I5(fdat[5]),
        .O(\nir_id[14]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h55551011)) 
    \nir_id[14]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[14]_i_4_n_0 ),
        .I2(\nir_id[14]_i_5_n_0 ),
        .I3(\nir_id[14]_i_6_n_0 ),
        .I4(fdat[15]),
        .O(\nir_id[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h88A82020)) 
    \nir_id[14]_i_3 
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[11]),
        .I4(fdat[12]),
        .O(\nir_id[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h3F3E3F3F3F3F3F3F)) 
    \nir_id[14]_i_4 
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat_0_sn_1),
        .I4(\nir_id[14]_i_7_n_0 ),
        .I5(\nir_id[14]_i_8_n_0 ),
        .O(\nir_id[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000F755FFFFFFFF)) 
    \nir_id[14]_i_5 
       (.I0(fdat[10]),
        .I1(fdat[2]),
        .I2(fdat[8]),
        .I3(\nir_id[14]_i_9_n_0 ),
        .I4(\nir_id[14]_i_10_n_0 ),
        .I5(fdat[14]),
        .O(\nir_id[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAAAAABAAAAA)) 
    \nir_id[14]_i_6 
       (.I0(\nir_id[14]_i_11_n_0 ),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[2]),
        .O(\nir_id[14]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[14]_i_7 
       (.I0(fdat[3]),
        .I1(fdat[2]),
        .O(\nir_id[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \nir_id[14]_i_8 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .I2(fdat_5_sn_1),
        .I3(\nir_id[19]_i_7_n_0 ),
        .I4(fdat[10]),
        .I5(fdat[11]),
        .O(\nir_id[14]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h00B3)) 
    \nir_id[14]_i_9 
       (.I0(fdat[6]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .I3(fdat[9]),
        .O(\nir_id[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF6FFFFFFFFFF)) 
    \nir_id[15]_i_1 
       (.I0(fdat[11]),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(fdat[15]),
        .I5(fdat_12_sn_1),
        .O(lir_id_0[15]));
  LUT3 #(
    .INIT(8'h80)) 
    \nir_id[15]_i_2 
       (.I0(fdat[12]),
        .I1(fdat[14]),
        .I2(fdat[13]),
        .O(fdat_12_sn_1));
  LUT6 #(
    .INIT(64'hE0E0E000EEEEEEEE)) 
    \nir_id[16]_i_1 
       (.I0(\nir_id[18]_i_2_n_0 ),
        .I1(fdat[8]),
        .I2(\nir_id[16]_i_2_n_0 ),
        .I3(\nir_id[16]_i_3_n_0 ),
        .I4(fdat[3]),
        .I5(\nir_id[18]_i_3_n_0 ),
        .O(lir_id_0[16]));
  LUT5 #(
    .INIT(32'hFFFFFB00)) 
    \nir_id[16]_i_2 
       (.I0(fdat[0]),
        .I1(fdat[8]),
        .I2(\nir_id[18]_i_7_n_0 ),
        .I3(fdat[9]),
        .I4(\nir_id[16]_i_4_n_0 ),
        .O(\nir_id[16]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[16]_i_3 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00FF00FFFFFF08FF)) 
    \nir_id[16]_i_4 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[8]),
        .I3(\nir_id[16]_i_3_n_0 ),
        .I4(fdat[3]),
        .I5(fdat[9]),
        .O(\nir_id[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h1500555555405555)) 
    \nir_id[17]_i_1 
       (.I0(\nir_id[17]_i_2_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[4]),
        .I4(\nir_id[18]_i_3_n_0 ),
        .I5(\nir_id[17]_i_3_n_0 ),
        .O(lir_id_0[17]));
  LUT6 #(
    .INIT(64'h000000000AA2AAAA)) 
    \nir_id[17]_i_2 
       (.I0(fdat[15]),
        .I1(fdat[11]),
        .I2(fdat[12]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(fdat[9]),
        .O(\nir_id[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEE0FEE00EE0FEE0F)) 
    \nir_id[17]_i_3 
       (.I0(\nir_id[17]_i_4_n_0 ),
        .I1(\nir_id[17]_i_5_n_0 ),
        .I2(fdat[4]),
        .I3(fdat[9]),
        .I4(fdat[8]),
        .I5(\nir_id[18]_i_8_n_0 ),
        .O(\nir_id[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D0000000)) 
    \nir_id[17]_i_4 
       (.I0(fdat[5]),
        .I1(fdat[3]),
        .I2(fdat[6]),
        .I3(fdat[7]),
        .I4(fdat[8]),
        .I5(fdat[1]),
        .O(\nir_id[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000033)) 
    \nir_id[17]_i_5 
       (.I0(\nir_id[17]_i_6_n_0 ),
        .I1(fdat[7]),
        .I2(fdat[1]),
        .I3(\nir_id[17]_i_7_n_0 ),
        .I4(fdat[3]),
        .I5(fdat[6]),
        .O(\nir_id[17]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[17]_i_6 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(\nir_id[17]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h5F5F5F4F)) 
    \nir_id[17]_i_7 
       (.I0(fdat[6]),
        .I1(fdat[1]),
        .I2(fdat[8]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .O(\nir_id[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h2E00EEEEEEC0EEEE)) 
    \nir_id[18]_i_1 
       (.I0(\nir_id[18]_i_2_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[5]),
        .I4(\nir_id[18]_i_3_n_0 ),
        .I5(\nir_id[18]_i_4_n_0 ),
        .O(lir_id_0[18]));
  LUT5 #(
    .INIT(32'hD5D57555)) 
    \nir_id[18]_i_2 
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .I2(fdat[13]),
        .I3(fdat[11]),
        .I4(fdat[12]),
        .O(\nir_id[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \nir_id[18]_i_3 
       (.I0(\nir_id[18]_i_5_n_0 ),
        .I1(\nir_id[18]_i_6_n_0 ),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[12]),
        .O(\nir_id[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h100010001F001F0F)) 
    \nir_id[18]_i_4 
       (.I0(fdat[2]),
        .I1(\nir_id[18]_i_7_n_0 ),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(\nir_id[18]_i_8_n_0 ),
        .I5(fdat[5]),
        .O(\nir_id[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4400444404440000)) 
    \nir_id[18]_i_5 
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(\nir_id[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h3020103030001000)) 
    \nir_id[18]_i_6 
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[18]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h55FFF57E)) 
    \nir_id[18]_i_7 
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .O(\nir_id[18]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[18]_i_8 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[18]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000A460FFFF)) 
    \nir_id[19]_i_1 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(fdat[15]),
        .I5(\nir_id[19]_i_2_n_0 ),
        .O(lir_id_0[19]));
  LUT6 #(
    .INIT(64'h000000005555F7FF)) 
    \nir_id[19]_i_2 
       (.I0(\nir_id[16]_i_3_n_0 ),
        .I1(\nir_id[19]_i_3_n_0 ),
        .I2(\nir_id[19]_i_4_n_0 ),
        .I3(fdat[9]),
        .I4(\nir_id[19]_i_5_n_0 ),
        .I5(\nir_id[19]_i_6_n_0 ),
        .O(\nir_id[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7FEFFFF)) 
    \nir_id[19]_i_3 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[3]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[7]),
        .O(\nir_id[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h4C0C000000000000)) 
    \nir_id[19]_i_4 
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[3]),
        .I4(fdat[8]),
        .I5(fdat[7]),
        .O(\nir_id[19]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \nir_id[19]_i_5 
       (.I0(fdat[9]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .O(\nir_id[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h555555555555D555)) 
    \nir_id[19]_i_6 
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(\nir_id[19]_i_7_n_0 ),
        .I2(fdat[11]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(\nir_id[19]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[19]_i_7 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[19]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[20]_i_5 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(fdat_5_sn_1));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[21]_i_3 
       (.I0(fdat[0]),
        .I1(fdat[1]),
        .O(fdat_0_sn_1));
  LUT6 #(
    .INIT(64'h0000000301020202)) 
    \nir_id[24]_i_10 
       (.I0(fdat[1]),
        .I1(\nir_id[24]_i_13_n_0 ),
        .I2(fdat[13]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[0]),
        .O(\nir_id[24]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_11 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[24]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_12 
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .O(\nir_id[24]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \nir_id[24]_i_13 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[12]),
        .O(\nir_id[24]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFBBFB)) 
    \nir_id[24]_i_2 
       (.I0(\nir_id[24]_i_5_n_0 ),
        .I1(\nir_id[24]_i_6_n_0 ),
        .I2(\nir_id[24]_i_7_n_0 ),
        .I3(\nir_id[24]_i_8_n_0 ),
        .I4(\nir_id_reg[24]_0 ),
        .I5(fdat[15]),
        .O(lir_id_0[24]));
  LUT4 #(
    .INIT(16'h0060)) 
    \nir_id[24]_i_5 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .O(\nir_id[24]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hCFDFFFDFFFDFFFDF)) 
    \nir_id[24]_i_6 
       (.I0(\nir_id[24]_i_10_n_0 ),
        .I1(\nir_id[24]_i_11_n_0 ),
        .I2(\nir_id[24]_i_12_n_0 ),
        .I3(fdat[9]),
        .I4(fdat[7]),
        .I5(fdat[12]),
        .O(\nir_id[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h950000FF150000FF)) 
    \nir_id[24]_i_7 
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[3]),
        .O(\nir_id[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5EFFFFFFFFFFFFFF)) 
    \nir_id[24]_i_8 
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[10]),
        .I3(fdat[8]),
        .I4(fdat[11]),
        .I5(fdat[12]),
        .O(\nir_id[24]_i_8_n_0 ));
  FDRE \nir_id_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[12]),
        .Q(nir_id[12]),
        .R(SR));
  FDRE \nir_id_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[13]),
        .Q(nir_id[13]),
        .R(SR));
  FDRE \nir_id_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[14]),
        .Q(nir_id[14]),
        .R(SR));
  FDRE \nir_id_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[15]),
        .Q(nir_id[15]),
        .R(SR));
  FDRE \nir_id_reg[16] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[16]),
        .Q(nir_id[16]),
        .R(SR));
  FDRE \nir_id_reg[17] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[17]),
        .Q(nir_id[17]),
        .R(SR));
  FDRE \nir_id_reg[18] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[18]),
        .Q(nir_id[18]),
        .R(SR));
  FDRE \nir_id_reg[19] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[19]),
        .Q(nir_id[19]),
        .R(SR));
  FDRE \nir_id_reg[20] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [0]),
        .Q(nir_id[20]),
        .R(SR));
  FDRE \nir_id_reg[21] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(\nir_id_reg[21]_0 [1]),
        .Q(nir_id[21]),
        .R(SR));
  FDRE \nir_id_reg[24] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(lir_id_0[24]),
        .Q(nir_id[24]),
        .R(SR));
  FDRE \nir_reg[0] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[0]),
        .Q(nir[0]),
        .R(SR));
  FDRE \nir_reg[10] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[10]),
        .Q(nir[10]),
        .R(SR));
  FDRE \nir_reg[11] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[11]),
        .Q(nir[11]),
        .R(SR));
  FDRE \nir_reg[12] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[12]),
        .Q(nir[12]),
        .R(SR));
  FDRE \nir_reg[13] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[13]),
        .Q(nir[13]),
        .R(SR));
  FDRE \nir_reg[14] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[14]),
        .Q(nir[14]),
        .R(SR));
  FDRE \nir_reg[15] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[15]),
        .Q(nir[15]),
        .R(SR));
  FDRE \nir_reg[1] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[1]),
        .Q(nir[1]),
        .R(SR));
  FDRE \nir_reg[2] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[2]),
        .Q(nir[2]),
        .R(SR));
  FDRE \nir_reg[3] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[3]),
        .Q(nir[3]),
        .R(SR));
  FDRE \nir_reg[4] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[4]),
        .Q(nir[4]),
        .R(SR));
  FDRE \nir_reg[5] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[5]),
        .Q(nir[5]),
        .R(SR));
  FDRE \nir_reg[6] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[6]),
        .Q(nir[6]),
        .R(SR));
  FDRE \nir_reg[7] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[7]),
        .Q(nir[7]),
        .R(SR));
  FDRE \nir_reg[8] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[8]),
        .Q(nir[8]),
        .R(SR));
  FDRE \nir_reg[9] 
       (.C(clk),
        .CE(fch_nir_lir),
        .D(fdat[9]),
        .Q(nir[9]),
        .R(SR));
  LUT2 #(
    .INIT(4'h2)) 
    \pc0[15]_i_2 
       (.I0(fch_issu1),
        .I1(\stat_reg[0]_51 ),
        .O(\stat_reg[0] ));
  FDRE \pc0_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[0]),
        .Q(\pc0_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc0_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[10]),
        .Q(\pc0_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc0_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[11]),
        .Q(\pc0_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc0_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[12]),
        .Q(\pc0_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc0_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(D[0]),
        .Q(\pc0_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc0_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(D[1]),
        .Q(\pc0_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc0_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(D[2]),
        .Q(\pc0_reg[15]_0 [15]),
        .R(SR));
  FDRE \pc0_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[1]),
        .Q(\pc0_reg[15]_0 [1]),
        .R(SR));
  FDRE \pc0_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[2]),
        .Q(\pc0_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc0_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[3]),
        .Q(\pc0_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc0_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[4]),
        .Q(\pc0_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc0_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[5]),
        .Q(\pc0_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc0_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[6]),
        .Q(\pc0_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc0_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[7]),
        .Q(\pc0_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc0_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[8]),
        .Q(\pc0_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc0_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[9]),
        .Q(\pc0_reg[15]_0 [9]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry
       (.CI(\<const0> ),
        .CO({pc10_carry_n_0,pc10_carry_n_1,pc10_carry_n_2,pc10_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,fch_pc[1],\<const0> }),
        .O({pc10_carry_n_4,pc10_carry_n_5,pc10_carry_n_6,pc10_carry_n_7}),
        .S({fctl_n_85,fctl_n_86,fctl_n_87,fctl_n_88}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry__0
       (.CI(pc10_carry_n_0),
        .CO({pc10_carry__0_n_0,pc10_carry__0_n_1,pc10_carry__0_n_2,pc10_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({pc10_carry__0_n_4,pc10_carry__0_n_5,pc10_carry__0_n_6,pc10_carry__0_n_7}),
        .S({fctl_n_150,fctl_n_151,fctl_n_152,fctl_n_153}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry__1
       (.CI(pc10_carry__0_n_0),
        .CO({pc10_carry__1_n_0,pc10_carry__1_n_1,pc10_carry__1_n_2,pc10_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({pc10_carry__1_n_4,pc10_carry__1_n_5,pc10_carry__1_n_6,pc10_carry__1_n_7}),
        .S({fctl_n_154,fctl_n_155,fctl_n_156,fctl_n_157}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 pc10_carry__2
       (.CI(pc10_carry__1_n_0),
        .CO({pc10_carry__2_n_1,pc10_carry__2_n_2,pc10_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({pc10_carry__2_n_4,pc10_carry__2_n_5,pc10_carry__2_n_6,pc10_carry__2_n_7}),
        .S({\pc1_reg[15]_1 ,fctl_n_158}));
  FDRE \pc1_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_7),
        .Q(\pc1_reg[15]_0 [0]),
        .R(SR));
  FDRE \pc1_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_5),
        .Q(\pc1_reg[15]_0 [10]),
        .R(SR));
  FDRE \pc1_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_4),
        .Q(\pc1_reg[15]_0 [11]),
        .R(SR));
  FDRE \pc1_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_7),
        .Q(\pc1_reg[15]_0 [12]),
        .R(SR));
  FDRE \pc1_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_6),
        .Q(\pc1_reg[15]_0 [13]),
        .R(SR));
  FDRE \pc1_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_5),
        .Q(\pc1_reg[15]_0 [14]),
        .R(SR));
  FDRE \pc1_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__2_n_4),
        .Q(\pc1_reg[15]_0 [15]),
        .R(SR));
  FDSE \pc1_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_6),
        .Q(\pc1_reg[15]_0 [1]),
        .S(SR));
  FDRE \pc1_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_5),
        .Q(\pc1_reg[15]_0 [2]),
        .R(SR));
  FDRE \pc1_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry_n_4),
        .Q(\pc1_reg[15]_0 [3]),
        .R(SR));
  FDRE \pc1_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_7),
        .Q(\pc1_reg[15]_0 [4]),
        .R(SR));
  FDRE \pc1_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_6),
        .Q(\pc1_reg[15]_0 [5]),
        .R(SR));
  FDRE \pc1_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_5),
        .Q(\pc1_reg[15]_0 [6]),
        .R(SR));
  FDRE \pc1_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__0_n_4),
        .Q(\pc1_reg[15]_0 [7]),
        .R(SR));
  FDRE \pc1_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_7),
        .Q(\pc1_reg[15]_0 [8]),
        .R(SR));
  FDRE \pc1_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(pc10_carry__1_n_6),
        .Q(\pc1_reg[15]_0 [9]),
        .R(SR));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \pc[14]_i_5 
       (.I0(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb_reg[14] ),
        .I2(\rgf_c0bus_wb_reg[15] [2]),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\pc[14]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \pc[15]_i_7 
       (.I0(fch_term),
        .I1(fctl_n_67),
        .O(\stat[2]_i_4 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[0]_i_1 
       (.I0(\rgf_c0bus_wb[0]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb_reg[3] [0]),
        .I3(\rgf_c0bus_wb_reg[0] ),
        .I4(\rgf_c0bus_wb_reg[0]_i_4_n_0 ),
        .O(\cbus_i[15] [0]));
  LUT6 #(
    .INIT(64'hF00070F000002000)) 
    \rgf_c0bus_wb[0]_i_11 
       (.I0(\stat_reg[2]_10 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .I2(\stat_reg[0]_2 ),
        .I3(a0bus_0[0]),
        .I4(\tr_reg[0]_0 ),
        .I5(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h3333744700007447)) 
    \rgf_c0bus_wb[0]_i_12 
       (.I0(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(a0bus_0[0]),
        .I3(\stat_reg[2]_10 ),
        .I4(\stat_reg[1]_1 ),
        .I5(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rgf_c0bus_wb[0]_i_14 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\tr_reg[0]_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\bbus_o[3]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \rgf_c0bus_wb[0]_i_15 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\tr_reg[0]_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_3_0 ),
        .I5(a0bus_0[0]),
        .O(\rgf_c0bus_wb[0]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c0bus_wb[0]_i_16 
       (.I0(\tr_reg[0]_0 ),
        .I1(\stat_reg[1]_2 ),
        .I2(a0bus_0[0]),
        .O(\rgf_c0bus_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE000000AE00)) 
    \rgf_c0bus_wb[0]_i_2 
       (.I0(\rgf_c0bus_wb[0]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_7_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFBBBBBBB)) 
    \rgf_c0bus_wb[0]_i_5 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[0]_i_2_0 ),
        .I2(\stat_reg[1]_1 ),
        .I3(a0bus_0[15]),
        .I4(\ccmd[0]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[3]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAEBF)) 
    \rgf_c0bus_wb[0]_i_6 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[13]_i_2_2 ),
        .I3(\rgf_c0bus_wb[0]_i_2_1 ),
        .O(\rgf_c0bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFAEEAAAA)) 
    \rgf_c0bus_wb[0]_i_7 
       (.I0(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_3_0 ),
        .I2(\rgf_c0bus_wb[13]_i_2_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFBFFBBB)) 
    \rgf_c0bus_wb[0]_i_8 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[8]_2 ),
        .I4(\rgf_c0bus_wb_reg[8]_1 ),
        .O(\rgf_c0bus_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDDDFFF)) 
    \rgf_c0bus_wb[0]_i_9 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I2(\sr[4]_i_66_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[5]_i_2_0 ),
        .I5(\rgf_c0bus_wb[11]_i_11_0 ),
        .O(\rgf_c0bus_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA8808FFFFFFFF)) 
    \rgf_c0bus_wb[10]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_7_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\rgf_c0bus_wb[10]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_5_n_0 ),
        .O(\cbus_i[15] [10]));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[10]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_3_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_58_0 ),
        .O(\rgf_c0bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF0F1F0F0F0F1F1F1)) 
    \rgf_c0bus_wb[10]_i_12 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\badr[15]_INST_0_i_2 ),
        .I3(\rgf_c0bus_wb[10]_i_4_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .I5(\rgf_c0bus_wb[10]_i_4_1 ),
        .O(\rgf_c0bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0400044404440444)) 
    \rgf_c0bus_wb[10]_i_13 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\rgf_c0bus_wb[10]_i_4_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I5(\sr[4]_i_60_2 ),
        .O(\rgf_c0bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0001110155555555)) 
    \rgf_c0bus_wb[10]_i_15 
       (.I0(\tr_reg[4] ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[10]_i_4_0 ),
        .I5(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[10]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[10]_i_16 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(a0bus_0[9]),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\rgf_c0bus_wb[10]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c0bus_wb[10]_i_23 
       (.I0(\bbus_o[0]_INST_0_i_1_0 ),
        .I1(a0bus_0[15]),
        .I2(\tr_reg[0]_0 ),
        .I3(a0bus_0[14]),
        .O(\rgf_c0bus_wb[10]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h82880808)) 
    \rgf_c0bus_wb[10]_i_25 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\bdatw[10]_0 ),
        .I3(\stat_reg[2]_10 ),
        .I4(a0bus_0[10]),
        .O(\rgf_c0bus_wb[10]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00550055030003FF)) 
    \rgf_c0bus_wb[10]_i_26 
       (.I0(\rgf_c0bus_wb[2]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_i_17_0 ),
        .I2(\rgf_c0bus_wb_reg[10]_i_17_1 ),
        .I3(\stat_reg[1]_1 ),
        .I4(\rgf_c0bus_wb_reg[10]_i_17_2 ),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[10]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h5101)) 
    \rgf_c0bus_wb[10]_i_3 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[10]_3 ),
        .O(\rgf_c0bus_wb[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \rgf_c0bus_wb[10]_i_4 
       (.I0(\rgf_c0bus_wb[10]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb_reg[10]_1 ),
        .I4(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h1101)) 
    \rgf_c0bus_wb[10]_i_5 
       (.I0(\rgf_c0bus_wb_reg[10]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_0 ),
        .I2(\rgf_c0bus_wb_reg[11]_0 [2]),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00B00000)) 
    \rgf_c0bus_wb[11]_i_1 
       (.I0(\rgf_c0bus_wb[11]_i_2_n_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\rgf_c0bus_wb[11]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_6_n_0 ),
        .O(\cbus_i[15] [11]));
  LUT5 #(
    .INIT(32'h56666666)) 
    \rgf_c0bus_wb[11]_i_11 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\tr_reg[0]_0 ),
        .I4(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\bbus_o[2]_INST_0_i_1_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[11]_i_12 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c0bus_wb[11]_i_14 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_3 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[11]_i_4_0 ),
        .O(\rgf_c0bus_wb[11]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h55FFD5F7)) 
    \rgf_c0bus_wb[11]_i_15 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb_reg[11]_2 ),
        .I3(a0bus_0[15]),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[11]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c0bus_wb[11]_i_16 
       (.I0(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I1(\sr[4]_i_60_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_65_0 ),
        .I4(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00011101)) 
    \rgf_c0bus_wb[11]_i_17 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[11]_i_5_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb_reg[11]_2 ),
        .O(\rgf_c0bus_wb[11]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[11]_i_18 
       (.I0(a0bus_0[10]),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1D110000)) 
    \rgf_c0bus_wb[11]_i_19 
       (.I0(\sr[4]_i_72_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\stat_reg[1]_1 ),
        .I3(\rgf_c0bus_wb[3]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000F000F3F5F3F5)) 
    \rgf_c0bus_wb[11]_i_2 
       (.I0(\rgf_c0bus_wb[11]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_2 ),
        .I2(\tr_reg[4] ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb_reg[11]_1 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[11]_i_21 
       (.I0(\tr_reg[0]_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\bbus_o[1]_INST_0_i_1_2 ));
  LUT3 #(
    .INIT(8'h56)) 
    \rgf_c0bus_wb[11]_i_22 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\tr_reg[0]_0 ),
        .O(\bbus_o[0]_INST_0_i_1_0 ));
  LUT5 #(
    .INIT(32'h0000A708)) 
    \rgf_c0bus_wb[11]_i_27 
       (.I0(a0bus_0[11]),
        .I1(\stat_reg[2]_10 ),
        .I2(bdatw_11_sn_1),
        .I3(\stat_reg[1]_1 ),
        .I4(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[11]_i_3 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(\stat_reg[2]_10 ));
  LUT6 #(
    .INIT(64'h88888880AAAAAAAA)) 
    \rgf_c0bus_wb[11]_i_4 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I2(\stat_reg[1]_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb_reg[11]_3 ),
        .I5(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFBAAAA)) 
    \rgf_c0bus_wb[11]_i_5 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[11]_i_6 
       (.I0(\rgf_c0bus_wb[11]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11] ),
        .I2(\rgf_c0bus_wb_reg[11]_0 [3]),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[11]_i_7 
       (.I0(\bbus_o[1]_INST_0_i_1_2 ),
        .I1(a0bus_0[15]),
        .O(\rgf_c0bus_wb[11]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hA999)) 
    \rgf_c0bus_wb[11]_i_9 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\tr_reg[0]_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\bbus_o[1]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4440)) 
    \rgf_c0bus_wb[12]_i_1 
       (.I0(\rgf_c0bus_wb[12]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_7_0 ),
        .I2(\tr_reg[4] ),
        .I3(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .O(\cbus_i[15] [12]));
  LUT6 #(
    .INIT(64'hF0F1F0F1F0F0F1F1)) 
    \rgf_c0bus_wb[12]_i_10 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_3_0 ),
        .I4(\rgf_c0bus_wb[12]_i_3_1 ),
        .I5(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[12]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h08FBFFFF)) 
    \rgf_c0bus_wb[12]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_3_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_0 ),
        .I3(a0bus_0[15]),
        .I4(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[12]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2EFF)) 
    \rgf_c0bus_wb[12]_i_12 
       (.I0(\tr_reg[4] ),
        .I1(\stat_reg[1]_2 ),
        .I2(a0bus_0[12]),
        .I3(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFF14)) 
    \rgf_c0bus_wb[12]_i_13 
       (.I0(\stat_reg[1]_1 ),
        .I1(a0bus_0[12]),
        .I2(\stat_reg[2]_10 ),
        .I3(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000882A88EA)) 
    \rgf_c0bus_wb[12]_i_15 
       (.I0(\stat_reg[1]_1 ),
        .I1(a0bus_0[12]),
        .I2(\stat_reg[2]_10 ),
        .I3(bdatw_12_sn_1),
        .I4(\ccmd[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h1555)) 
    \rgf_c0bus_wb[12]_i_18 
       (.I0(\bbus_o[1]_INST_0_i_1_0 ),
        .I1(a0bus_0[0]),
        .I2(\tr_reg[0]_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\bbus_o[1]_INST_0_i_1_1 ));
  LUT6 #(
    .INIT(64'h3400F4F43400F400)) 
    \rgf_c0bus_wb[12]_i_2 
       (.I0(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(\tr_reg[4] ),
        .I3(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb_reg[12]_0 ),
        .I5(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hD5D5D500D5D5D5D5)) 
    \rgf_c0bus_wb[12]_i_3 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(a0bus_0[11]),
        .I3(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF444F444FFFFF444)) 
    \rgf_c0bus_wb[12]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [0]),
        .I2(cbus_i[8]),
        .I3(\stat_reg[0]_3 ),
        .I4(bdatr[3]),
        .I5(\rgf_c0bus_wb_reg[9]_2 ),
        .O(\rgf_c0bus_wb[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF7500)) 
    \rgf_c0bus_wb[12]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb_reg[12] ),
        .I3(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c0bus_wb[12]_i_6 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[12]_i_3_0 ),
        .O(\rgf_c0bus_wb[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF111F000)) 
    \rgf_c0bus_wb[12]_i_7 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb_reg[4]_1 ),
        .I3(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_2_0 ),
        .I5(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[12]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[12]_i_9 
       (.I0(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I1(\sr[4]_i_68_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_68_0 ),
        .O(\rgf_c0bus_wb[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hE000FFFFFFFFFFFF)) 
    \rgf_c0bus_wb[13]_i_1 
       (.I0(\rgf_c0bus_wb[13]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_6_n_0 ),
        .O(\cbus_i[15] [13]));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[13]_i_10 
       (.I0(\stat_reg[1]_1 ),
        .I1(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[11]_i_3_0 ));
  LUT4 #(
    .INIT(16'h2AAA)) 
    \rgf_c0bus_wb[13]_i_11 
       (.I0(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(a0bus_0[15]),
        .I3(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[13]_i_12 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[5]_i_3_0 ),
        .O(\rgf_c0bus_wb[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF111F000)) 
    \rgf_c0bus_wb[13]_i_13 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_4_0 ),
        .I4(\rgf_c0bus_wb_reg[4]_2 ),
        .I5(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[13]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h1141004155414441)) 
    \rgf_c0bus_wb[13]_i_16 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[13]),
        .I3(\stat_reg[1]_1 ),
        .I4(a0bus_0[5]),
        .I5(bbus_o_7_sn_1),
        .O(\rgf_c0bus_wb[13]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    \rgf_c0bus_wb[13]_i_17 
       (.I0(\stat_reg[1]_2 ),
        .I1(\rgf_c0bus_wb_reg[5] ),
        .I2(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I3(a0bus_0[13]),
        .I4(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[13]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0000C60C)) 
    \rgf_c0bus_wb[13]_i_18 
       (.I0(\stat_reg[2]_10 ),
        .I1(\stat_reg[1]_1 ),
        .I2(bbus_o_13_sn_1),
        .I3(a0bus_0[13]),
        .I4(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFE000000FEFEFEFE)) 
    \rgf_c0bus_wb[13]_i_2 
       (.I0(\rgf_c0bus_wb[13]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_3_0 ),
        .I4(a0bus_0[12]),
        .I5(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hEAAA)) 
    \rgf_c0bus_wb[13]_i_23 
       (.I0(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\stat_reg[1]_1 ),
        .I3(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h40000000)) 
    \rgf_c0bus_wb[13]_i_25 
       (.I0(\tr_reg[4] ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\tr_reg[0]_0 ),
        .I4(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h2023)) 
    \rgf_c0bus_wb[13]_i_3 
       (.I0(\stat_reg[1]_1 ),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\stat_reg[0]_2 ),
        .I3(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_7_0 ));
  LUT6 #(
    .INIT(64'hADFF0D0DADFF0DFF)) 
    \rgf_c0bus_wb[13]_i_4 
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I2(\tr_reg[4] ),
        .I3(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb_reg[13] ),
        .I5(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0BBB0BBB00000BBB)) 
    \rgf_c0bus_wb[13]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [1]),
        .I2(cbus_i[9]),
        .I3(\stat_reg[0]_3 ),
        .I4(bdatr[4]),
        .I5(\rgf_c0bus_wb_reg[9]_2 ),
        .O(\rgf_c0bus_wb[13]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h001F)) 
    \rgf_c0bus_wb[13]_i_6 
       (.I0(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00011101)) 
    \rgf_c0bus_wb[13]_i_7 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[13]_i_2_2 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[13]_i_2_1 ),
        .O(\rgf_c0bus_wb[13]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[13]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_2_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[0]_i_2_1 ),
        .O(\rgf_c0bus_wb[13]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \rgf_c0bus_wb[13]_i_9 
       (.I0(\badr[15]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[5]_i_3_1 ),
        .I2(\stat_reg[1]_1 ),
        .I3(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[14]_i_1 
       (.I0(\rgf_c0bus_wb[14]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb_reg[15] [2]),
        .I3(\rgf_c0bus_wb_reg[14] ),
        .I4(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .O(\cbus_i[15] [14]));
  LUT5 #(
    .INIT(32'hD0D0D000)) 
    \rgf_c0bus_wb[14]_i_10 
       (.I0(bbus_o_6_sn_1),
        .I1(\stat_reg[1]_2 ),
        .I2(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I3(a0bus_0[14]),
        .I4(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[14]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h0000A708)) 
    \rgf_c0bus_wb[14]_i_11 
       (.I0(a0bus_0[14]),
        .I1(\stat_reg[2]_10 ),
        .I2(bbus_o_14_sn_1),
        .I3(\stat_reg[1]_1 ),
        .I4(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF0F1F0F0F0F1F1F1)) 
    \rgf_c0bus_wb[14]_i_13 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\stat_reg[2]_10 ),
        .I3(\rgf_c0bus_wb[14]_i_5_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .I5(\rgf_c0bus_wb_reg[10]_3 ),
        .O(\rgf_c0bus_wb[14]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \rgf_c0bus_wb[14]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I1(\sr[4]_i_64_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[10]_2 ),
        .O(\rgf_c0bus_wb[14]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF47FFFF)) 
    \rgf_c0bus_wb[14]_i_15 
       (.I0(a0bus_0[14]),
        .I1(\tr_reg[0]_0 ),
        .I2(a0bus_0[15]),
        .I3(\bbus_o[0]_INST_0_i_1_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[14]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00004747FF000000)) 
    \rgf_c0bus_wb[14]_i_16 
       (.I0(\rgf_c0bus_wb[5]_i_3_2 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[9]_i_3_0 ),
        .I3(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .I4(\stat_reg[1]_1 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[14]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFFFEEE)) 
    \rgf_c0bus_wb[14]_i_17 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[10]_i_4_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\sr[4]_i_58_0 ),
        .I5(\badr[15]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[14]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hD0)) 
    \rgf_c0bus_wb[14]_i_18 
       (.I0(\stat_reg[2]_10 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .I2(\stat_reg[0]_2 ),
        .O(\stat_reg[1]_2 ));
  LUT6 #(
    .INIT(64'hEE00FA00EE000000)) 
    \rgf_c0bus_wb[14]_i_2 
       (.I0(\rgf_c0bus_wb[14]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb_reg[14]_0 ),
        .I2(\rgf_c0bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_7_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c0bus_wb[14]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[14]_i_4 
       (.I0(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h000D)) 
    \rgf_c0bus_wb[14]_i_5 
       (.I0(\stat_reg[1]_1 ),
        .I1(\sr[4]_i_16_0 ),
        .I2(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_c0bus_wb[14]_i_7 
       (.I0(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[14]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hD500D5D5)) 
    \rgf_c0bus_wb[14]_i_8 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(a0bus_0[13]),
        .I3(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hEEBEFFBEAABEBBBE)) 
    \rgf_c0bus_wb[14]_i_9 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[14]),
        .I3(\stat_reg[1]_1 ),
        .I4(a0bus_0[6]),
        .I5(bbus_o_7_sn_1),
        .O(\rgf_c0bus_wb[14]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[15]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15] [3]),
        .I2(\rgf_c0bus_wb_reg[15]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb_reg[15]_0 ),
        .O(\cbus_i[15] [15]));
  LUT5 #(
    .INIT(32'hA02A0080)) 
    \rgf_c0bus_wb[15]_i_10 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[15]),
        .I3(\bdatw[15] ),
        .I4(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00545555)) 
    \rgf_c0bus_wb[15]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I1(a0bus_0[7]),
        .I2(\stat_reg[2]_10 ),
        .I3(\rgf_c0bus_wb_reg[10]_i_17_0 ),
        .I4(\stat_reg[1]_1 ),
        .I5(\rgf_c0bus_wb[15]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[15]_i_12 
       (.I0(a0bus_0[14]),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF0F0000EE0E)) 
    \rgf_c0bus_wb[15]_i_13 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_4_1 ),
        .I4(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_4_2 ),
        .O(\rgf_c0bus_wb[15]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_c0bus_wb[15]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_4_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .O(\rgf_c0bus_wb[15]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c0bus_wb[15]_i_15 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[7]_3 ),
        .O(\rgf_c0bus_wb[15]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c0bus_wb[15]_i_16 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[11]_i_4_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[2]_i_2_0 ),
        .O(\rgf_c0bus_wb[15]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hAABE)) 
    \rgf_c0bus_wb[15]_i_17 
       (.I0(\stat_reg[0]_2 ),
        .I1(a0bus_0[15]),
        .I2(\stat_reg[2]_10 ),
        .I3(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[15]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hD0D0D000)) 
    \rgf_c0bus_wb[15]_i_19 
       (.I0(bbus_o_7_sn_1),
        .I1(\stat_reg[1]_2 ),
        .I2(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I3(a0bus_0[15]),
        .I4(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFAAFFFFD0DDDDDD)) 
    \rgf_c0bus_wb[15]_i_2 
       (.I0(\stat_reg[1]_1 ),
        .I1(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I2(\ccmd[1]_INST_0_i_1_n_0 ),
        .I3(\stat_reg[2]_10 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_20 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[15]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \rgf_c0bus_wb[15]_i_22 
       (.I0(a0bus_0[15]),
        .I1(\stat_reg[1]_1 ),
        .I2(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[15]_i_24 
       (.I0(\tr_reg[4] ),
        .I1(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F02020F000202)) 
    \rgf_c0bus_wb[15]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_6 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .O(\stat_reg[1]_1 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[15]_i_7 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_8 
       (.I0(\sr[5]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[15]_i_9 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(\stat_reg[0]_2 ));
  LUT5 #(
    .INIT(32'hFFFFB080)) 
    \rgf_c0bus_wb[1]_i_1 
       (.I0(\rgf_c0bus_wb[1]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_4_n_0 ),
        .O(\cbus_i[15] [1]));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[1]_i_10 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[1]_i_3_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[9]_i_3_0 ),
        .O(\rgf_c0bus_wb[1]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1011)) 
    \rgf_c0bus_wb[1]_i_11 
       (.I0(\rgf_c0bus_wb[1]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .I3(\stat_reg[1]_1 ),
        .I4(\rgf_c0bus_wb[1]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAAABE)) 
    \rgf_c0bus_wb[1]_i_13 
       (.I0(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\stat_reg[2]_10 ),
        .I3(\stat_reg[1]_1 ),
        .I4(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[1]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hD100)) 
    \rgf_c0bus_wb[1]_i_14 
       (.I0(a0bus_0[1]),
        .I1(\stat_reg[1]_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h41044500)) 
    \rgf_c0bus_wb[1]_i_15 
       (.I0(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\stat_reg[1]_1 ),
        .I4(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[1]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h00FB)) 
    \rgf_c0bus_wb[1]_i_2 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb_reg[9]_0 ),
        .I3(\rgf_c0bus_wb[1]_i_5_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F0E0E0F0F000E)) 
    \rgf_c0bus_wb[1]_i_3 
       (.I0(\rgf_c0bus_wb_reg[1] ),
        .I1(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_8_n_0 ),
        .I3(\stat_reg[2]_10 ),
        .I4(\rgf_c0bus_wb[1]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFEA)) 
    \rgf_c0bus_wb[1]_i_4 
       (.I0(\rgf_c0bus_wb[1]_i_11_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(cbus_i[0]),
        .I3(\rgf_c0bus_wb_reg[1]_0 ),
        .I4(\rgf_c0bus_wb_reg[3] [1]),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5F5FCFCF0F000F0F)) 
    \rgf_c0bus_wb[1]_i_5 
       (.I0(\rgf_c0bus_wb_reg[10]_3 ),
        .I1(\rgf_c0bus_wb_reg[10]_2 ),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .I3(\badr[1]_INST_0_i_2 ),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEAAAAAAA)) 
    \rgf_c0bus_wb[1]_i_7 
       (.I0(\stat_reg[2]_10 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\tr_reg[0]_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I5(\tr_reg[4] ),
        .O(\rgf_c0bus_wb[1]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[1]_i_8 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\rgf_c0bus_wb[1]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c0bus_wb[1]_i_9 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[5]_i_3_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_58_0 ),
        .O(\rgf_c0bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4440)) 
    \rgf_c0bus_wb[2]_i_1 
       (.I0(\rgf_c0bus_wb[2]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_7_0 ),
        .I2(\tr_reg[4] ),
        .I3(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .O(\cbus_i[15] [2]));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[2]_i_10 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[10]_i_4_0 ),
        .O(\rgf_c0bus_wb[2]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c0bus_wb[2]_i_11 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\sr[4]_i_65_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_60_0 ),
        .O(\rgf_c0bus_wb[2]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[2]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\rgf_c0bus_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0D0F0000)) 
    \rgf_c0bus_wb[2]_i_13 
       (.I0(\stat_reg[1]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c0bus_wb[2]_i_15 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAEAAAEAABFBB)) 
    \rgf_c0bus_wb[2]_i_16 
       (.I0(\stat_reg[1]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(\ccmd[0]_INST_0_i_1_n_0 ),
        .I4(\stat_reg[2]_10 ),
        .I5(a0bus_0[2]),
        .O(\rgf_c0bus_wb[2]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000A708)) 
    \rgf_c0bus_wb[2]_i_17 
       (.I0(a0bus_0[2]),
        .I1(\stat_reg[2]_10 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(\stat_reg[1]_1 ),
        .I4(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA8AAA8AAA8A8)) 
    \rgf_c0bus_wb[2]_i_2 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb_reg[2] ),
        .I2(\rgf_c0bus_wb[2]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_3_0 ),
        .I4(\rgf_c0bus_wb_reg[2]_0 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFEE0E)) 
    \rgf_c0bus_wb[2]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .I2(\stat_reg[2]_10 ),
        .I3(\rgf_c0bus_wb[2]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFEA)) 
    \rgf_c0bus_wb[2]_i_4 
       (.I0(\rgf_c0bus_wb[2]_i_13_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(cbus_i[1]),
        .I3(\rgf_c0bus_wb_reg[2]_1 ),
        .I4(\rgf_c0bus_wb_reg[3] [2]),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    \rgf_c0bus_wb[2]_i_6 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb[2]_i_2_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\sr[4]_i_64_1 ),
        .O(\rgf_c0bus_wb[2]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c0bus_wb[2]_i_8 
       (.I0(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_4_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[10]_i_4_1 ),
        .I4(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4777000000000000)) 
    \rgf_c0bus_wb[2]_i_9 
       (.I0(\rgf_c0bus_wb[10]_i_4_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I3(\sr[4]_i_60_2 ),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .I5(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[3]_i_1 
       (.I0(\rgf_c0bus_wb[3]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb_reg[3] [3]),
        .I3(\rgf_c0bus_wb_reg[3]_0 ),
        .I4(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .O(\cbus_i[15] [3]));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[3]_i_10 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c0bus_wb[3]_i_11 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[3]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hF8F9FDF9)) 
    \rgf_c0bus_wb[3]_i_12 
       (.I0(\stat_reg[2]_10 ),
        .I1(a0bus_0[3]),
        .I2(\stat_reg[1]_1 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h41044500)) 
    \rgf_c0bus_wb[3]_i_13 
       (.I0(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I1(a0bus_0[3]),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(\stat_reg[1]_1 ),
        .I4(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[3]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[3]_i_14 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\sr[4]_i_68_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_68_0 ),
        .O(\rgf_c0bus_wb[3]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h45405555)) 
    \rgf_c0bus_wb[3]_i_15 
       (.I0(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[11]_i_5_0 ),
        .I4(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h2E000000)) 
    \rgf_c0bus_wb[3]_i_16 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb_reg[11]_2 ),
        .I3(\bbus_o[2]_INST_0_i_1_0 ),
        .I4(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h47440000FFFFFFFF)) 
    \rgf_c0bus_wb[3]_i_17 
       (.I0(\rgf_c0bus_wb_reg[11]_2 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_2 ),
        .I3(a0bus_0[15]),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .I5(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[3]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[3]_i_18 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(\rgf_c0bus_wb_reg[8]_4 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[7]_2 ),
        .O(\rgf_c0bus_wb[3]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF0200020)) 
    \rgf_c0bus_wb[3]_i_2 
       (.I0(\rgf_c0bus_wb[3]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\tr_reg[4] ),
        .I4(\rgf_c0bus_wb[3]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0F0D0000)) 
    \rgf_c0bus_wb[3]_i_4 
       (.I0(\stat_reg[1]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[3]_i_5 
       (.I0(a0bus_0[2]),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h08AA)) 
    \rgf_c0bus_wb[3]_i_6 
       (.I0(\rgf_c0bus_wb[3]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2000022722272)) 
    \rgf_c0bus_wb[3]_i_7 
       (.I0(\bbus_o[1]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_1 ),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .I3(\rgf_c0bus_wb_reg[11]_3 ),
        .I4(\rgf_c0bus_wb[3]_i_18_n_0 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF80B08080)) 
    \rgf_c0bus_wb[4]_i_1 
       (.I0(\rgf_c0bus_wb[4]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\rgf_c0bus_wb[4]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_5_n_0 ),
        .O(\cbus_i[15] [4]));
  LUT6 #(
    .INIT(64'h0000000004000444)) 
    \rgf_c0bus_wb[4]_i_10 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[4]_i_3_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[4]_i_3_1 ),
        .I5(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h50001540)) 
    \rgf_c0bus_wb[4]_i_13 
       (.I0(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[4]),
        .I3(\stat_reg[1]_1 ),
        .I4(\tr_reg[4] ),
        .O(\rgf_c0bus_wb[4]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hD5FF)) 
    \rgf_c0bus_wb[4]_i_14 
       (.I0(\stat_reg[1]_1 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hAABE)) 
    \rgf_c0bus_wb[4]_i_15 
       (.I0(\stat_reg[0]_2 ),
        .I1(a0bus_0[4]),
        .I2(\stat_reg[2]_10 ),
        .I3(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c0bus_wb[4]_i_16 
       (.I0(a0bus_0[4]),
        .I1(\stat_reg[1]_2 ),
        .I2(\tr_reg[4] ),
        .I3(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFF4F4F4)) 
    \rgf_c0bus_wb[4]_i_17 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_0 [0]),
        .I2(\rgf_c0bus_wb[4]_i_5_0 ),
        .I3(cbus_i[3]),
        .I4(\stat_reg[0]_3 ),
        .O(\rgf_c0bus_wb[4]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0035F035)) 
    \rgf_c0bus_wb[4]_i_2 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb_reg[4]_1 ),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb_reg[4]_2 ),
        .O(\rgf_c0bus_wb[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \rgf_c0bus_wb[4]_i_20 
       (.I0(\rgf_c0bus_wb[4]_i_6_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_1 ),
        .I2(p_0_in),
        .I3(p_1_in),
        .I4(\tr_reg[0]_1 ),
        .I5(\tr_reg[0]_0 ),
        .O(\rgf_c0bus_wb[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F20000F20000)) 
    \rgf_c0bus_wb[4]_i_3 
       (.I0(\rgf_c0bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_10_n_0 ),
        .I2(\stat_reg[2]_10 ),
        .I3(\bbus_o[2]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb_reg[4] ),
        .I5(\rgf_c0bus_wb_reg[4]_0 ),
        .O(\rgf_c0bus_wb[4]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[4]_i_4 
       (.I0(a0bus_0[3]),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAEEEE)) 
    \rgf_c0bus_wb[4]_i_5 
       (.I0(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FFFF00FF)) 
    \rgf_c0bus_wb[4]_i_6 
       (.I0(\rgf_c0bus_wb[4]_i_2_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[4]_i_2_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_20_n_0 ),
        .I5(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[4]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h55551555)) 
    \rgf_c0bus_wb[4]_i_9 
       (.I0(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\bbus_o[2]_INST_0_i_1_0 ),
        .I3(a0bus_0[15]),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF54)) 
    \rgf_c0bus_wb[5]_i_1 
       (.I0(\rgf_c0bus_wb[5]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_5_n_0 ),
        .O(\cbus_i[15] [5]));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c0bus_wb[5]_i_10 
       (.I0(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_2_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[13]_i_2_2 ),
        .I4(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[5]_i_11 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(a0bus_0[4]),
        .O(\rgf_c0bus_wb[5]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[5]_i_12 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[9]_i_3_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[5]_i_3_2 ),
        .O(\rgf_c0bus_wb[5]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c0bus_wb[5]_i_13 
       (.I0(\rgf_c0bus_wb[5]_i_3_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h2222220202022202)) 
    \rgf_c0bus_wb[5]_i_15 
       (.I0(\rgf_c0bus_wb[5]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I2(\stat_reg[1]_1 ),
        .I3(a0bus_0[13]),
        .I4(\stat_reg[2]_10 ),
        .I5(\rgf_c0bus_wb_reg[5] ),
        .O(\rgf_c0bus_wb[5]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[5]_i_16 
       (.I0(\ccmd[3]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[5]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFF9F8F9F8F9F8F9)) 
    \rgf_c0bus_wb[5]_i_17 
       (.I0(\stat_reg[2]_10 ),
        .I1(a0bus_0[5]),
        .I2(\stat_reg[1]_1 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\stat_reg[1]_2 ),
        .I5(\rgf_c0bus_wb_reg[5] ),
        .O(\rgf_c0bus_wb[5]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFD00FFFF)) 
    \rgf_c0bus_wb[5]_i_2 
       (.I0(\rgf_c0bus_wb[5]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb_reg[5]_1 ),
        .I2(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I3(\tr_reg[4] ),
        .I4(\rgf_c0bus_wb[15]_i_7_0 ),
        .O(\rgf_c0bus_wb[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hDD0DFF0F0000FF0F)) 
    \rgf_c0bus_wb[5]_i_3 
       (.I0(\rgf_c0bus_wb[5]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFF4F4F4)) 
    \rgf_c0bus_wb[5]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_0 [1]),
        .I2(\rgf_c0bus_wb_reg[5]_0 ),
        .I3(cbus_i[4]),
        .I4(\stat_reg[0]_3 ),
        .O(\rgf_c0bus_wb[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAABEFAFAAA)) 
    \rgf_c0bus_wb[5]_i_5 
       (.I0(\rgf_c0bus_wb[5]_i_15_n_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(\stat_reg[1]_1 ),
        .I3(a0bus_0[5]),
        .I4(\rgf_c0bus_wb_reg[5] ),
        .I5(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c0bus_wb[5]_i_6 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(\rgf_c0bus_wb[5]_i_2_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\badr[1]_INST_0_i_2 ),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[5]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    \rgf_c0bus_wb[5]_i_8 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb[5]_i_2_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[5]_i_2_0 ),
        .O(\rgf_c0bus_wb[5]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c0bus_wb[5]_i_9 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\rgf_c0bus_wb[5]_i_3_1 ),
        .O(\rgf_c0bus_wb[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFB080)) 
    \rgf_c0bus_wb[6]_i_1 
       (.I0(\rgf_c0bus_wb[6]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .O(\cbus_i[15] [6]));
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \rgf_c0bus_wb[6]_i_10 
       (.I0(\sr[4]_i_65_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[10]_i_4_0 ),
        .I3(\stat_reg[2]_10 ),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .I5(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[6]_i_11 
       (.I0(\sr[4]_i_70_0 ),
        .I1(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hF2F0D0F0)) 
    \rgf_c0bus_wb[6]_i_13 
       (.I0(\bbus_o[1]_INST_0_i_1_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_0 ),
        .I2(a0bus_0[15]),
        .I3(\tr_reg[0]_0 ),
        .I4(a0bus_0[14]),
        .O(\rgf_c0bus_wb[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hEEBEFFBEAABEBBBE)) 
    \rgf_c0bus_wb[6]_i_15 
       (.I0(\stat_reg[1]_2 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[6]),
        .I3(\stat_reg[1]_1 ),
        .I4(a0bus_0[14]),
        .I5(bbus_o_6_sn_1),
        .O(\rgf_c0bus_wb[6]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h41044500)) 
    \rgf_c0bus_wb[6]_i_16 
       (.I0(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I1(a0bus_0[6]),
        .I2(bbus_o_6_sn_1),
        .I3(\stat_reg[1]_1 ),
        .I4(\stat_reg[2]_10 ),
        .O(\rgf_c0bus_wb[6]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00003F05)) 
    \rgf_c0bus_wb[6]_i_2 
       (.I0(\rgf_c0bus_wb_reg[6]_0 ),
        .I1(\rgf_c0bus_wb_reg[6]_1 ),
        .I2(\bbus_o[2]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[11]_i_3_0 ),
        .I4(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EE0E0E0E)) 
    \rgf_c0bus_wb[6]_i_3 
       (.I0(\rgf_c0bus_wb[6]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I3(a0bus_0[5]),
        .I4(\rgf_c0bus_wb[11]_i_3_0 ),
        .I5(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFEA)) 
    \rgf_c0bus_wb[6]_i_4 
       (.I0(\rgf_c0bus_wb[6]_i_11_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(cbus_i[5]),
        .I3(\rgf_c0bus_wb_reg[6] ),
        .I4(\rgf_c0bus_wb_reg[7]_0 [2]),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    \rgf_c0bus_wb[6]_i_7 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\sr[4]_i_64_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb_reg[10]_2 ),
        .O(\rgf_c0bus_wb[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h888888880F000FFF)) 
    \rgf_c0bus_wb[6]_i_8 
       (.I0(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\sr[4]_i_65_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[10]_i_4_0 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[6]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c0bus_wb[6]_i_9 
       (.I0(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_4_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_58_0 ),
        .I4(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBF008C00)) 
    \rgf_c0bus_wb[7]_i_1 
       (.I0(\rgf_c0bus_wb[7]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_7_0 ),
        .I4(\rgf_c0bus_wb[7]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_5_n_0 ),
        .O(\cbus_i[15] [7]));
  LUT6 #(
    .INIT(64'hFF00FF007F00FF00)) 
    \rgf_c0bus_wb[7]_i_13 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\tr_reg[0]_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(\stat_reg[2]_10 ),
        .I4(a0bus_0[15]),
        .I5(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[7]_i_14 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[1]_1 ),
        .I2(a0bus_0[7]),
        .I3(\stat_reg[2]_10 ),
        .I4(bbus_o_7_sn_1),
        .O(\rgf_c0bus_wb[7]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c0bus_wb[7]_i_2 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[7]_3 ),
        .O(\rgf_c0bus_wb[7]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[7]_i_3 
       (.I0(\rgf_c0bus_wb[11]_i_11_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[11]_3 ),
        .O(\rgf_c0bus_wb[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAB000000ABABABAB)) 
    \rgf_c0bus_wb[7]_i_4 
       (.I0(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb_reg[7]_1 ),
        .I3(\rgf_c0bus_wb[11]_i_3_0 ),
        .I4(a0bus_0[6]),
        .I5(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFEA)) 
    \rgf_c0bus_wb[7]_i_5 
       (.I0(\rgf_c0bus_wb_reg[7]_i_11_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(cbus_i[6]),
        .I3(\rgf_c0bus_wb_reg[7] ),
        .I4(\rgf_c0bus_wb_reg[7]_0 [3]),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[7]_i_7 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[11]_i_11_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF02A2)) 
    \rgf_c0bus_wb[7]_i_9 
       (.I0(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I1(\sr[4]_i_60_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[11]_i_5_0 ),
        .I4(\badr[15]_INST_0_i_2 ),
        .I5(\rgf_c0bus_wb[7]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBF008C00)) 
    \rgf_c0bus_wb[8]_i_1 
       (.I0(\rgf_c0bus_wb[8]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[8]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_7_0 ),
        .I4(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_5_n_0 ),
        .O(\cbus_i[15] [8]));
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \rgf_c0bus_wb[8]_i_10 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\tr_reg[0]_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[0]),
        .I4(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\rgf_c0bus_wb[8]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0047FFFF00470047)) 
    \rgf_c0bus_wb[8]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_3_1 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\sr[4]_i_68_0 ),
        .I3(\rgf_c0bus_wb[11]_i_11_0 ),
        .I4(\stat_reg[2]_10 ),
        .I5(\badr[15]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8F88FFFF8F880000)) 
    \rgf_c0bus_wb[8]_i_13 
       (.I0(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I3(\sr[4]_i_71_0 ),
        .I4(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c0bus_wb[8]_i_15 
       (.I0(\tr_reg[0]_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[8]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFF14)) 
    \rgf_c0bus_wb[8]_i_16 
       (.I0(\stat_reg[1]_1 ),
        .I1(a0bus_0[8]),
        .I2(\stat_reg[2]_10 ),
        .I3(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[8]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h82880808)) 
    \rgf_c0bus_wb[8]_i_18 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\bdatw[8]_0 ),
        .I3(\stat_reg[2]_10 ),
        .I4(a0bus_0[8]),
        .O(\rgf_c0bus_wb[8]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[8]_i_2 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb_reg[8]_3 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb_reg[8]_4 ),
        .O(\rgf_c0bus_wb[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hCAFF0000FFFFFFFF)) 
    \rgf_c0bus_wb[8]_i_3 
       (.I0(\rgf_c0bus_wb_reg[8]_1 ),
        .I1(\rgf_c0bus_wb_reg[8]_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[11]_i_3_0 ),
        .I4(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAE000000AEAEAEAE)) 
    \rgf_c0bus_wb[8]_i_4 
       (.I0(\rgf_c0bus_wb[8]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb_reg[8]_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[11]_i_3_0 ),
        .I4(a0bus_0[7]),
        .I5(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[8]_i_5 
       (.I0(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb_reg[8] ),
        .I2(\rgf_c0bus_wb_reg[11]_0 [0]),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFB080)) 
    \rgf_c0bus_wb[9]_i_1 
       (.I0(\rgf_c0bus_wb[9]_i_2_n_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\rgf_c0bus_wb[9]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_5_n_0 ),
        .O(\cbus_i[15] [9]));
  LUT4 #(
    .INIT(16'h2700)) 
    \rgf_c0bus_wb[9]_i_10 
       (.I0(\bbus_o[1]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[13]_i_2_2 ),
        .I2(\rgf_c0bus_wb[0]_i_2_1 ),
        .I3(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAABABFAAAA)) 
    \rgf_c0bus_wb[9]_i_11 
       (.I0(\badr[15]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[9]_i_3_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[9]_i_3_1 ),
        .I4(\stat_reg[1]_1 ),
        .I5(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[9]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA8A80)) 
    \rgf_c0bus_wb[9]_i_12 
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[9]_i_3_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\rgf_c0bus_wb[1]_i_3_0 ),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\rgf_c0bus_wb[9]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[9]_i_13 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(a0bus_0[8]),
        .O(\rgf_c0bus_wb[9]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c0bus_wb[9]_i_14 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_10 ),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[9]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[9]_i_15 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[1]_1 ),
        .O(\rgf_c0bus_wb[9]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFF14)) 
    \rgf_c0bus_wb[9]_i_16 
       (.I0(\stat_reg[1]_1 ),
        .I1(a0bus_0[9]),
        .I2(\stat_reg[2]_10 ),
        .I3(\stat_reg[0]_2 ),
        .O(\rgf_c0bus_wb[9]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h41440404)) 
    \rgf_c0bus_wb[9]_i_18 
       (.I0(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(bdatw_9_sn_1),
        .I3(\stat_reg[2]_10 ),
        .I4(a0bus_0[9]),
        .O(\rgf_c0bus_wb[9]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hA3A3A3A30303F303)) 
    \rgf_c0bus_wb[9]_i_2 
       (.I0(\rgf_c0bus_wb_reg[9]_0 ),
        .I1(\rgf_c0bus_wb_reg[9]_1 ),
        .I2(\bbus_o[2]_INST_0_i_1_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\badr[1]_INST_0_i_2 ),
        .I5(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\rgf_c0bus_wb[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00FE00FE000000FE)) 
    \rgf_c0bus_wb[9]_i_3 
       (.I0(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF444F444FFFFF444)) 
    \rgf_c0bus_wb[9]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_0 [1]),
        .I2(cbus_i[7]),
        .I3(\stat_reg[0]_3 ),
        .I4(bdatr[0]),
        .I5(\rgf_c0bus_wb_reg[9]_2 ),
        .O(\rgf_c0bus_wb[9]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8F880000)) 
    \rgf_c0bus_wb[9]_i_5 
       (.I0(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb_reg[9] ),
        .I4(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c0bus_wb[9]_i_8 
       (.I0(\bbus_o[0]_INST_0_i_1_0 ),
        .I1(a0bus_0[0]),
        .I2(\tr_reg[0]_0 ),
        .I3(a0bus_0[1]),
        .O(\badr[1]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h00011101)) 
    \rgf_c0bus_wb[9]_i_9 
       (.I0(\stat_reg[1]_1 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[13]_i_2_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[9]_i_3_0 ),
        .O(\rgf_c0bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[0]_i_4 
       (.I0(\rgf_c0bus_wb[0]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_12_n_0 ),
        .O(\rgf_c0bus_wb_reg[0]_i_4_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_7_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[10]_i_17 
       (.I0(\rgf_c0bus_wb[10]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_26_n_0 ),
        .O(\rgf_c0bus_wb_reg[10]_i_17_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_7_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[15]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c0bus_wb_reg[15]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_7_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[7]_i_11 
       (.I0(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I1(\sr[4]_i_69_0 ),
        .O(\rgf_c0bus_wb_reg[7]_i_11_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFEFE)) 
    \rgf_c1bus_wb[0]_i_1 
       (.I0(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_4_n_0 ),
        .I3(tout__1_carry_i_11_0),
        .I4(\rgf_c1bus_wb_reg[3]_2 [0]),
        .I5(\rgf_c1bus_wb_reg[0]_0 ),
        .O(\bdatr[15] [0]));
  LUT4 #(
    .INIT(16'hAEBF)) 
    \rgf_c1bus_wb[0]_i_10 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\sr[4]_i_36_0 ),
        .I3(\sr[4]_i_25_0 ),
        .O(\rgf_c1bus_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFAEEAAAA)) 
    \rgf_c1bus_wb[0]_i_11 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\sr[4]_i_39_0 ),
        .I2(\rgf_c1bus_wb[0]_i_4_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF808A0000)) 
    \rgf_c1bus_wb[0]_i_13 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_37_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[0]_i_4_1 ),
        .I4(\stat_reg[2]_8 ),
        .I5(\rgf_c1bus_wb[0]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0500053005000500)) 
    \rgf_c1bus_wb[0]_i_14 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\rgf_c1bus_wb[0]_i_18_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[15]),
        .I4(\rgf_c1bus_wb[0]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hAA8A)) 
    \rgf_c1bus_wb[0]_i_15 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[15]),
        .I3(ir1[11]),
        .O(\rgf_c1bus_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA88AA88AAAA8A)) 
    \rgf_c1bus_wb[0]_i_16 
       (.I0(\rgf_c1bus_wb[0]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_22_n_0 ),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .I4(ir1[3]),
        .I5(ir1[1]),
        .O(\rgf_c1bus_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0400FFFF)) 
    \rgf_c1bus_wb[0]_i_17 
       (.I0(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\stat_reg[2]_8 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[4]_0 ),
        .O(\rgf_c1bus_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FDD0FDDD)) 
    \rgf_c1bus_wb[0]_i_18 
       (.I0(rst_n_fl_reg_9),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h11000015)) 
    \rgf_c1bus_wb[0]_i_19 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .O(\rgf_c1bus_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hCB000800CF000000)) 
    \rgf_c1bus_wb[0]_i_2 
       (.I0(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\tr_reg[0] ),
        .I3(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0400)) 
    \rgf_c1bus_wb[0]_i_20 
       (.I0(\bdatw[15]_INST_0_i_188_n_0 ),
        .I1(ir1[9]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_c1bus_wb[0]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_24_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBF3BBF3A)) 
    \rgf_c1bus_wb[0]_i_21 
       (.I0(ir1[14]),
        .I1(ir1[15]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(tout__1_carry_i_15_n_0),
        .I5(\rgf_c1bus_wb[0]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF77F)) 
    \rgf_c1bus_wb[0]_i_22 
       (.I0(\fadr[15]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_16_0 ),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(ir1[2]),
        .I4(\badr[15]_INST_0_i_153_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_61_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h52501000)) 
    \rgf_c1bus_wb[0]_i_23 
       (.I0(ir1[5]),
        .I1(ir1[3]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .O(\rgf_c1bus_wb[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00FE000000051111)) 
    \rgf_c1bus_wb[0]_i_24 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\rgf_c1bus_wb[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h00400000FFFFFFFF)) 
    \rgf_c1bus_wb[0]_i_25 
       (.I0(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I1(ir1[6]),
        .I2(ir1[8]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[7]),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0090)) 
    \rgf_c1bus_wb[0]_i_26 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(\rgf_c1bus_wb[0]_i_27_n_0 ),
        .I3(ir1[15]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\rgf_selc1_wb_reg[1] [2]),
        .O(\rgf_c1bus_wb[0]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[0]_i_27 
       (.I0(ir1[11]),
        .I1(ir1[13]),
        .O(\rgf_c1bus_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h00C0CCC000440044)) 
    \rgf_c1bus_wb[0]_i_3 
       (.I0(\rgf_c1bus_wb[0]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\stat_reg[2]_6 ),
        .I4(\tr_reg[0] ),
        .I5(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAE00AE)) 
    \rgf_c1bus_wb[0]_i_4 
       (.I0(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb_reg[0] ),
        .I4(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFFFFABAFAFA)) 
    \rgf_c1bus_wb[0]_i_6 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_c1bus_wb[0]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [2]),
        .I4(ir1[14]),
        .I5(\rgf_c1bus_wb[0]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hA0AF3F30)) 
    \rgf_c1bus_wb[0]_i_7 
       (.I0(\tr_reg[0] ),
        .I1(a1bus_0[8]),
        .I2(\stat_reg[1]_0 ),
        .I3(a1bus_0[0]),
        .I4(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0111)) 
    \rgf_c1bus_wb[0]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I3(\stat_reg[2]_4 ),
        .O(\stat_reg[2]_6 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAFEAE)) 
    \rgf_c1bus_wb[0]_i_9 
       (.I0(\tr_reg[4]_0 ),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\stat_reg[1]_0 ),
        .I3(a1bus_0[15]),
        .I4(\stat_reg[2]_4 ),
        .I5(\bdatw[11]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h10111010FFFFFFFF)) 
    \rgf_c1bus_wb[10]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[10] ),
        .I2(\tr_reg[4]_0 ),
        .I3(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .O(\bdatr[15] [10]));
  LUT4 #(
    .INIT(16'h5404)) 
    \rgf_c1bus_wb[10]_i_10 
       (.I0(\bdatw[8]_INST_0_i_16_1 ),
        .I1(a1bus_0[15]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[14]),
        .O(\badr[14]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hFF07000700000000)) 
    \rgf_c1bus_wb[10]_i_12 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[8]_INST_0_i_16_1 ),
        .I2(\badr[14]_INST_0_i_1 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb_reg[10]_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[10]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h5140)) 
    \rgf_c1bus_wb[10]_i_13 
       (.I0(\stat_reg[1]_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb_reg[10]_0 ),
        .I3(\sr[4]_i_44_0 ),
        .O(\rgf_c1bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF0D0000)) 
    \rgf_c1bus_wb[10]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\sr[4]_i_52_0 ),
        .I2(\rgf_c1bus_wb[10]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h11111FF1)) 
    \rgf_c1bus_wb[10]_i_16 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(a1bus_0[10]),
        .I3(\stat_reg[2]_4 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[10]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hE200)) 
    \rgf_c1bus_wb[10]_i_17 
       (.I0(\bdatw[10]_INST_0_i_16_n_0 ),
        .I1(\stat_reg[2]_6 ),
        .I2(a1bus_0[10]),
        .I3(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hC0007800)) 
    \rgf_c1bus_wb[10]_i_18 
       (.I0(\stat_reg[2]_4 ),
        .I1(a1bus_0[10]),
        .I2(\stat_reg[1]_0 ),
        .I3(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I4(bdatw_10_sn_1),
        .O(\rgf_c1bus_wb[10]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFBBBFAAAAAAAA)) 
    \rgf_c1bus_wb[10]_i_3 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\bdatw[9]_INST_0_i_16_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\badr[14]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb_reg[10]_0 ),
        .I5(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF101F1010)) 
    \rgf_c1bus_wb[10]_i_4 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\rgf_c1bus_wb_reg[1] ),
        .I5(\rgf_c1bus_wb[15]_i_14_1 ),
        .O(\rgf_c1bus_wb[10]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h51510051)) 
    \rgf_c1bus_wb[10]_i_5 
       (.I0(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I1(bdatr[1]),
        .I2(\rgf_c1bus_wb_reg[12] ),
        .I3(\rgf_c1bus_wb_reg[11] [0]),
        .I4(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[10]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hCCCC440C)) 
    \rgf_c1bus_wb[10]_i_9 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(a1bus_0[9]),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[10]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAABBABAAAAAAAA)) 
    \rgf_c1bus_wb[11]_i_1 
       (.I0(\rgf_c1bus_wb[11]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_6_n_0 ),
        .O(\bdatr[15] [11]));
  LUT4 #(
    .INIT(16'h6566)) 
    \rgf_c1bus_wb[11]_i_10 
       (.I0(\bdatw[10]_INST_0_i_16_n_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\bdatw[9]_INST_0_i_16_n_0 ),
        .I3(\tr_reg[0] ),
        .O(\bdatw[8]_INST_0_i_16_0 ));
  LUT4 #(
    .INIT(16'hFD5D)) 
    \rgf_c1bus_wb[11]_i_11 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_3 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[11]_i_3_0 ),
        .O(\rgf_c1bus_wb[11]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[11]_i_12 
       (.I0(\bdatw[9]_INST_0_i_16_n_0 ),
        .I1(\tr_reg[0] ),
        .O(\bdatw[8]_INST_0_i_16_2 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[11]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(a1bus_0[10]),
        .I2(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[11]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF88FFA0FF88)) 
    \rgf_c1bus_wb[11]_i_16 
       (.I0(\stat_reg[1]_0 ),
        .I1(a1bus_0[15]),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[15]_i_14_1 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\rgf_c1bus_wb_reg[11]_0 ),
        .O(\rgf_c1bus_wb[11]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00022202)) 
    \rgf_c1bus_wb[11]_i_17 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\rgf_c1bus_wb[11]_i_6_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb_reg[11]_0 ),
        .O(\rgf_c1bus_wb[11]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00011101)) 
    \rgf_c1bus_wb[11]_i_18 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\sr[4]_i_33_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[15]_i_4_0 ),
        .O(\rgf_c1bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1100011100001000)) 
    \rgf_c1bus_wb[11]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(a1bus_0[11]),
        .I4(\bdatw[11]_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[11]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[11]_i_2 
       (.I0(\rgf_c1bus_wb_reg[11]_i_7_n_0 ),
        .I1(bdatr[2]),
        .I2(\rgf_c1bus_wb_reg[12] ),
        .I3(\rgf_c1bus_wb_reg[11] [1]),
        .I4(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1151)) 
    \rgf_c1bus_wb[11]_i_20 
       (.I0(\rgf_c1bus_wb[11]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(a1bus_0[3]),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb[11]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h11111FF1)) 
    \rgf_c1bus_wb[11]_i_21 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(a1bus_0[11]),
        .I3(\stat_reg[2]_4 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[11]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hA202)) 
    \rgf_c1bus_wb[11]_i_22 
       (.I0(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\stat_reg[2]_6 ),
        .I3(a1bus_0[11]),
        .O(\rgf_c1bus_wb[11]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h88888808AAAAAAAA)) 
    \rgf_c1bus_wb[11]_i_3 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[11]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb_reg[3]_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFF755F7)) 
    \rgf_c1bus_wb[11]_i_4 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(a1bus_0[15]),
        .I2(\bdatw[8]_INST_0_i_16_2 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb_reg[11]_0 ),
        .O(\rgf_c1bus_wb[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hF200FFFF)) 
    \rgf_c1bus_wb[11]_i_5 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_1 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hBBBBBBBA)) 
    \rgf_c1bus_wb[11]_i_6 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[11]_i_8 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_1 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45454500)) 
    \rgf_c1bus_wb[12]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\rgf_c1bus_wb[12]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .O(\bdatr[15] [12]));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[12]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(a1bus_0[11]),
        .O(\rgf_c1bus_wb[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000554555550010)) 
    \rgf_c1bus_wb[12]_i_12 
       (.I0(\stat_reg[1]_0 ),
        .I1(\bdatw[9]_INST_0_i_16_n_0 ),
        .I2(\tr_reg[0] ),
        .I3(\bdatw[10]_INST_0_i_16_n_0 ),
        .I4(\tr_reg[4]_0 ),
        .I5(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \rgf_c1bus_wb[12]_i_13 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\sr[6]_i_6_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[12]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hDFCCCCCC)) 
    \rgf_c1bus_wb[12]_i_14 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[2]_7 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(a1bus_0[15]),
        .O(\rgf_c1bus_wb[12]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h20202022)) 
    \rgf_c1bus_wb[12]_i_2 
       (.I0(\rgf_c1bus_wb[12]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\stat_reg[2]_8 ),
        .I4(\rgf_c1bus_wb_reg[12]_1 ),
        .O(\rgf_c1bus_wb[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h1100011100001000)) 
    \rgf_c1bus_wb[12]_i_22 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(a1bus_0[12]),
        .I4(\bdatw[12]_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[12]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1151)) 
    \rgf_c1bus_wb[12]_i_23 
       (.I0(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(a1bus_0[4]),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h11111FF1)) 
    \rgf_c1bus_wb[12]_i_24 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\stat_reg[2]_4 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[12]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hA202)) 
    \rgf_c1bus_wb[12]_i_25 
       (.I0(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\stat_reg[2]_6 ),
        .I3(a1bus_0[12]),
        .O(\rgf_c1bus_wb[12]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h00F2)) 
    \rgf_c1bus_wb[12]_i_3 
       (.I0(\stat_reg[2]_4 ),
        .I1(\rgf_c1bus_wb[12]_i_8_n_0 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\rgf_c1bus_wb[12]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAA20)) 
    \rgf_c1bus_wb[12]_i_4 
       (.I0(\rgf_c1bus_wb[12]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[12]_0 ),
        .I2(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[12]_i_5 
       (.I0(\rgf_c1bus_wb_reg[12]_i_15_n_0 ),
        .I1(bdatr[3]),
        .I2(\rgf_c1bus_wb_reg[12] ),
        .I3(\rgf_c1bus_wb_reg[15] [0]),
        .I4(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[12]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFD5D)) 
    \rgf_c1bus_wb[12]_i_6 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[6]_i_6_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[6]_i_9_0 ),
        .O(\rgf_c1bus_wb[12]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h20)) 
    \rgf_c1bus_wb[12]_i_8 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_25_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[12]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \rgf_c1bus_wb[12]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_14_0 ),
        .I1(\sr[4]_i_37_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb_reg[4]_1 ),
        .O(\rgf_c1bus_wb[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4540)) 
    \rgf_c1bus_wb[13]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_2_n_0 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb_reg[13] ),
        .I5(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .O(\bdatr[15] [13]));
  LUT6 #(
    .INIT(64'hAAABAAAAAAABABAB)) 
    \rgf_c1bus_wb[13]_i_11 
       (.I0(\rgf_c1bus_wb[15]_i_14_1 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_39_0 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\sr[4]_i_36_0 ),
        .O(\rgf_c1bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hD0FFFFFFD0D0D0D0)) 
    \rgf_c1bus_wb[13]_i_12 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(\stat_reg[2]_8 ),
        .I4(a1bus_0[12]),
        .I5(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c1bus_wb[13]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(a1bus_0[13]),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb[13]_i_5_0 ),
        .O(\rgf_c1bus_wb[13]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h06FF)) 
    \rgf_c1bus_wb[13]_i_14 
       (.I0(a1bus_0[13]),
        .I1(\stat_reg[2]_4 ),
        .I2(\stat_reg[1]_0 ),
        .I3(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h00007F4C)) 
    \rgf_c1bus_wb[13]_i_15 
       (.I0(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(tout__1_carry__0),
        .I3(a1bus_0[13]),
        .I4(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c1bus_wb[13]_i_17 
       (.I0(\bdatw[8]_INST_0_i_16_1 ),
        .I1(a1bus_0[0]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[1]),
        .O(\rgf_c1bus_wb[13]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h5F535053)) 
    \rgf_c1bus_wb[13]_i_2 
       (.I0(\rgf_c1bus_wb_reg[13]_1 ),
        .I1(\rgf_c1bus_wb[13]_i_7_n_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\stat_reg[2]_8 ),
        .I4(\rgf_c1bus_wb_reg[13]_2 ),
        .O(\rgf_c1bus_wb[13]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[13]_i_23 
       (.I0(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF880A)) 
    \rgf_c1bus_wb[13]_i_3 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[13]_6 ),
        .I2(\rgf_c1bus_wb_reg[13]_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\rgf_c1bus_wb[13]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAABAFF)) 
    \rgf_c1bus_wb[13]_i_5 
       (.I0(\rgf_c1bus_wb[13]_i_13_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(a1bus_0[5]),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c1bus_wb[13]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_2_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEFFFFEEEF)) 
    \rgf_c1bus_wb[14]_i_1 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_6_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\bdatr[15] [14]));
  LUT4 #(
    .INIT(16'hA202)) 
    \rgf_c1bus_wb[14]_i_11 
       (.I0(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_3_1 ),
        .I2(\stat_reg[2]_6 ),
        .I3(a1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[14]_i_12 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(tout__1_carry_i_13_n_0),
        .I2(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h9A220000)) 
    \rgf_c1bus_wb[14]_i_13 
       (.I0(\stat_reg[1]_0 ),
        .I1(\rgf_c1bus_wb[14]_i_3_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(a1bus_0[14]),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF757F)) 
    \rgf_c1bus_wb[14]_i_14 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(a1bus_0[14]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[15]),
        .I4(\bdatw[8]_INST_0_i_16_1 ),
        .O(\rgf_c1bus_wb[14]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[14]_i_15 
       (.I0(\stat_reg[2]_8 ),
        .I1(a1bus_0[13]),
        .O(\rgf_c1bus_wb[14]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF0F8)) 
    \rgf_c1bus_wb[14]_i_16 
       (.I0(\stat_reg[1]_0 ),
        .I1(a1bus_0[15]),
        .I2(\stat_reg[2]_7 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[15]_i_14_1 ));
  LUT5 #(
    .INIT(32'hDC8CCCCC)) 
    \rgf_c1bus_wb[14]_i_19 
       (.I0(\bdatw[8]_INST_0_i_16_1 ),
        .I1(a1bus_0[15]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[14]),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[14]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h0000002E)) 
    \rgf_c1bus_wb[14]_i_21 
       (.I0(\sr[4]_i_34_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\sr[4]_i_43_1 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[14]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDDFDD)) 
    \rgf_c1bus_wb[14]_i_22 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_43_0 ),
        .I4(\rgf_c1bus_wb[1]_i_2_0 ),
        .O(\rgf_c1bus_wb[14]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[14]_i_23 
       (.I0(tout__1_carry_i_13_n_0),
        .I1(\stat_reg[1]_6 ),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .O(\rgf_c1bus_wb[14]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000FB)) 
    \rgf_c1bus_wb[14]_i_24 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\bcmd[2]_INST_0_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_34_n_0 ),
        .I3(\stat_reg[1]_6 ),
        .I4(\rgf_c1bus_wb[14]_i_35_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[14]_i_25 
       (.I0(tout__1_carry_i_13_n_0),
        .I1(\rgf_c1bus_wb[14]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \rgf_c1bus_wb[14]_i_26 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAAAABABABAB)) 
    \rgf_c1bus_wb[14]_i_27 
       (.I0(\rgf_c1bus_wb[14]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_39_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_40_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_41_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_42_n_0 ),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[14]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hA9)) 
    \rgf_c1bus_wb[14]_i_28 
       (.I0(\bdatw[9]_INST_0_i_16_n_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\tr_reg[0] ),
        .O(\bdatw[8]_INST_0_i_16_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF510000)) 
    \rgf_c1bus_wb[14]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb_reg[14]_0 ),
        .I3(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h1F1F1F1F00001F0F)) 
    \rgf_c1bus_wb[14]_i_34 
       (.I0(ir1[8]),
        .I1(\rgf_c1bus_wb[14]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_44_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_45_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_46_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_c1bus_wb[14]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0200020000000200)) 
    \rgf_c1bus_wb[14]_i_35 
       (.I0(ir1[15]),
        .I1(ir1[13]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\read_cyc_reg[1] ),
        .I4(ir1[11]),
        .I5(ir1[14]),
        .O(\rgf_c1bus_wb[14]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000222F)) 
    \rgf_c1bus_wb[14]_i_36 
       (.I0(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_47_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\rgf_c1bus_wb[14]_i_48_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(ir1[12]),
        .O(\rgf_c1bus_wb[14]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF3AA)) 
    \rgf_c1bus_wb[14]_i_37 
       (.I0(\rgf_c1bus_wb[14]_i_49_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_50_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[11]),
        .I4(\rgf_c1bus_wb[14]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_52_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h82A2AAAA8222AAAA)) 
    \rgf_c1bus_wb[14]_i_38 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(\rgf_c1bus_wb[14]_i_53_0 ),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[14]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0057000000000000)) 
    \rgf_c1bus_wb[14]_i_39 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(rst_n_fl_reg_9),
        .I3(\rgf_selc1_rn_wb[1]_i_12_n_0 ),
        .I4(ir1[7]),
        .I5(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0D0FFD0)) 
    \rgf_c1bus_wb[14]_i_4 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I5(\tr_reg[4]_0 ),
        .O(\rgf_c1bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF5554)) 
    \rgf_c1bus_wb[14]_i_40 
       (.I0(\rgf_c1bus_wb[14]_i_53_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_54_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I3(ir1[6]),
        .I4(\rgf_c1bus_wb[14]_i_55_n_0 ),
        .I5(ir1[15]),
        .O(\rgf_c1bus_wb[14]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000880)) 
    \rgf_c1bus_wb[14]_i_41 
       (.I0(\rgf_c1bus_wb[14]_i_53_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[10]),
        .I4(ir1[7]),
        .I5(ir1[9]),
        .O(\rgf_c1bus_wb[14]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF5F1D551)) 
    \rgf_c1bus_wb[14]_i_42 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(ir1[9]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\rgf_c1bus_wb[14]_i_56_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_57_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0A0A0A0A22000000)) 
    \rgf_c1bus_wb[14]_i_43 
       (.I0(\rgf_c1bus_wb[14]_i_58_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[9]),
        .I3(ir1[6]),
        .I4(rst_n_fl_reg_9),
        .I5(ir1[10]),
        .O(\rgf_c1bus_wb[14]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0000EF2F00000000)) 
    \rgf_c1bus_wb[14]_i_44 
       (.I0(\rgf_c1bus_wb[14]_i_59_n_0 ),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .I3(\rgf_c1bus_wb[14]_i_60_n_0 ),
        .I4(ir1[15]),
        .I5(ir1[14]),
        .O(\rgf_c1bus_wb[14]_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hBBFFE0FF)) 
    \rgf_c1bus_wb[14]_i_45 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[11]),
        .I4(ir1[9]),
        .O(\rgf_c1bus_wb[14]_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[14]_i_46 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .O(\rgf_c1bus_wb[14]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    \rgf_c1bus_wb[14]_i_47 
       (.I0(\rgf_c1bus_wb[14]_i_61_n_0 ),
        .I1(\fadr[15]_INST_0_i_16_n_0 ),
        .I2(\rgf_selc1_wb_reg[1]_0 ),
        .I3(\rgf_c1bus_wb[14]_i_62_n_0 ),
        .I4(ir1[6]),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[14]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EFAFEFEF)) 
    \rgf_c1bus_wb[14]_i_48 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[13]),
        .I2(ir1[15]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .I5(\rgf_c1bus_wb[14]_i_63_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FFDF)) 
    \rgf_c1bus_wb[14]_i_49 
       (.I0(ir1[14]),
        .I1(ir1[15]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(\rgf_c1bus_wb[14]_i_64_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0545054055455540)) 
    \rgf_c1bus_wb[14]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_14_1 ),
        .I1(\rgf_c1bus_wb_reg[14]_1 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\rgf_c1bus_wb_reg[14]_2 ),
        .I5(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[14]_i_50 
       (.I0(ir1[12]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_c1bus_wb[14]_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hDFDFDFFF)) 
    \rgf_c1bus_wb[14]_i_51 
       (.I0(ir1[14]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(ir1[13]),
        .I3(ir1[15]),
        .I4(ir1[12]),
        .O(\rgf_c1bus_wb[14]_i_51_n_0 ));
  LUT5 #(
    .INIT(32'h0000BF00)) 
    \rgf_c1bus_wb[14]_i_52 
       (.I0(ir1[15]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(ir1[12]),
        .I4(rst_n_fl_reg_9),
        .O(\rgf_c1bus_wb[14]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1FF1FFFF)) 
    \rgf_c1bus_wb[14]_i_53 
       (.I0(ctl_fetch1_fl_i_20_n_0),
        .I1(rst_n_fl_reg_9),
        .I2(ir1[6]),
        .I3(ir1[7]),
        .I4(\stat[2]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_65_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0100010001000000)) 
    \rgf_c1bus_wb[14]_i_54 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[3]),
        .I2(ir1[1]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ir1[0]),
        .I5(ir1[2]),
        .O(\rgf_c1bus_wb[14]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \rgf_c1bus_wb[14]_i_55 
       (.I0(\rgf_c1bus_wb[14]_i_53_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I2(ir1[9]),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .I5(ir1[8]),
        .O(\rgf_c1bus_wb[14]_i_55_n_0 ));
  LUT5 #(
    .INIT(32'hF3F3F1FE)) 
    \rgf_c1bus_wb[14]_i_56 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[3]),
        .I4(ir1[4]),
        .O(\rgf_c1bus_wb[14]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFBEFFBEFFBEBFBE)) 
    \rgf_c1bus_wb[14]_i_57 
       (.I0(\rgf_c1bus_wb[14]_i_66_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[9]),
        .O(\rgf_c1bus_wb[14]_i_57_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[14]_i_58 
       (.I0(ir1[7]),
        .I1(ir1[11]),
        .O(\rgf_c1bus_wb[14]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hF000F00001050000)) 
    \rgf_c1bus_wb[14]_i_59 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(ir1[6]),
        .I2(ir1[10]),
        .I3(ir1[7]),
        .I4(rst_n_fl_reg_9),
        .I5(ir1[11]),
        .O(\rgf_c1bus_wb[14]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hD000D0D0D000D000)) 
    \rgf_c1bus_wb[14]_i_6 
       (.I0(\rgf_c1bus_wb_reg[14]_3 ),
        .I1(\stat_reg[2]_8 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb[14]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000800040)) 
    \rgf_c1bus_wb[14]_i_60 
       (.I0(ir1[7]),
        .I1(\stat[0]_i_22__0_n_0 ),
        .I2(ir1[11]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ir1[4]),
        .I5(ir1[5]),
        .O(\rgf_c1bus_wb[14]_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_c1bus_wb[14]_i_61 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .I3(ir1[4]),
        .O(\rgf_c1bus_wb[14]_i_61_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[14]_i_62 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .O(\rgf_c1bus_wb[14]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h0002020200000002)) 
    \rgf_c1bus_wb[14]_i_63 
       (.I0(\rgf_c1bus_wb[14]_i_67_n_0 ),
        .I1(ir1[14]),
        .I2(ir1[15]),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .I5(ir1[0]),
        .O(\rgf_c1bus_wb[14]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFE0F0FFFF)) 
    \rgf_c1bus_wb[14]_i_64 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[10]),
        .I3(ir1[6]),
        .I4(ir1[12]),
        .I5(\rgf_c1bus_wb[14]_i_68_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h77FF77FFFFFFFFFC)) 
    \rgf_c1bus_wb[14]_i_65 
       (.I0(\rgf_c1bus_wb[14]_i_53_0 ),
        .I1(ir1[7]),
        .I2(ir1[5]),
        .I3(ir1[8]),
        .I4(ir1[4]),
        .I5(ir1[12]),
        .O(\rgf_c1bus_wb[14]_i_65_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rgf_c1bus_wb[14]_i_66 
       (.I0(ir1[7]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .O(\rgf_c1bus_wb[14]_i_66_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[14]_i_67 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(ir1[2]),
        .I3(ir1[6]),
        .I4(ctl_fetch1_fl_i_36_n_0),
        .O(\rgf_c1bus_wb[14]_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFAA00C0)) 
    \rgf_c1bus_wb[14]_i_68 
       (.I0(ir1[10]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_c1bus_wb[14]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEF111F)) 
    \rgf_c1bus_wb[14]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h11111FF1)) 
    \rgf_c1bus_wb[14]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(a1bus_0[14]),
        .I3(\stat_reg[2]_4 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[14]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c1bus_wb[14]_i_9 
       (.I0(\stat_reg[1]_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_0 ),
        .I2(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4F4FFF4)) 
    \rgf_c1bus_wb[15]_i_1 
       (.I0(tout__1_carry_i_11_0),
        .I1(\rgf_c1bus_wb_reg[15] [1]),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I5(\rgf_c1bus_wb_reg[15]_0 ),
        .O(\bdatr[15] [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFF9020B000)) 
    \rgf_c1bus_wb[15]_i_10 
       (.I0(a1bus_0[15]),
        .I1(fch_leir_nir_reg),
        .I2(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[2]_4 ),
        .I5(\rgf_c1bus_wb[15]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFDFFDDD)) 
    \rgf_c1bus_wb[15]_i_11 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[11]_i_6_0 ),
        .I4(\rgf_c1bus_wb[15]_i_4_0 ),
        .O(\rgf_c1bus_wb[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000047)) 
    \rgf_c1bus_wb[15]_i_12 
       (.I0(\sr[4]_i_33_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb_reg[10]_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .I5(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hAA2A)) 
    \rgf_c1bus_wb[15]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(a1bus_0[15]),
        .I3(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[15]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h99999A99)) 
    \rgf_c1bus_wb[15]_i_14 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\bdatw[10]_INST_0_i_16_n_0 ),
        .I3(\tr_reg[0] ),
        .I4(\bdatw[9]_INST_0_i_16_n_0 ),
        .O(\bdatw[9]_INST_0_i_16_0 ));
  LUT5 #(
    .INIT(32'hAAAA2A20)) 
    \rgf_c1bus_wb[15]_i_16 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_3 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb_reg[3]_1 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_17 
       (.I0(\stat_reg[2]_4 ),
        .I1(\tr_reg[4]_0 ),
        .O(\rgf_c1bus_wb[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF0F00008808)) 
    \rgf_c1bus_wb[15]_i_19 
       (.I0(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(\rgf_c1bus_wb[15]_i_10_0 ),
        .I3(\stat_reg[2]_6 ),
        .I4(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[15]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(tout__1_carry_i_11_n_0),
        .O(tout__1_carry_i_11_0));
  LUT3 #(
    .INIT(8'hF8)) 
    \rgf_c1bus_wb[15]_i_23 
       (.I0(a1bus_0[15]),
        .I1(\stat_reg[1]_0 ),
        .I2(\stat_reg[2]_7 ),
        .O(\rgf_c1bus_wb[15]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \rgf_c1bus_wb[15]_i_24 
       (.I0(\tr_reg[4]_0 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\bdatw[10]_INST_0_i_16_n_0 ),
        .I3(\tr_reg[0] ),
        .I4(\bdatw[9]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFBFF)) 
    \rgf_c1bus_wb[15]_i_27 
       (.I0(\bdatw[9]_INST_0_i_16_n_0 ),
        .I1(\tr_reg[0] ),
        .I2(\bdatw[10]_INST_0_i_16_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\bdatw[11]_INST_0_i_16_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[15]_i_3 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBAAFBAAFBAAFB)) 
    \rgf_c1bus_wb[15]_i_4 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I4(\stat_reg[2]_8 ),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0D0FFD0)) 
    \rgf_c1bus_wb[15]_i_5 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[6]_2 ),
        .I2(\rgf_c1bus_wb[15]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb_reg[15]_1 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[15]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[15]_i_8 
       (.I0(\stat_reg[1]_0 ),
        .I1(\stat_reg[2]_4 ),
        .O(\stat_reg[2]_8 ));
  LUT6 #(
    .INIT(64'h22820082AA828882)) 
    \rgf_c1bus_wb[15]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(a1bus_0[15]),
        .I3(\stat_reg[1]_0 ),
        .I4(a1bus_0[7]),
        .I5(\rgf_c1bus_wb[15]_i_10_0 ),
        .O(\rgf_c1bus_wb[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55554454)) 
    \rgf_c1bus_wb[1]_i_1 
       (.I0(\rgf_c1bus_wb[1]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb_reg[1] ),
        .I3(\rgf_c1bus_wb[1]_i_5_n_0 ),
        .I4(\tr_reg[4]_0 ),
        .I5(\rgf_c1bus_wb[1]_i_6_n_0 ),
        .O(\bdatr[15] [1]));
  LUT5 #(
    .INIT(32'h00004E00)) 
    \rgf_c1bus_wb[1]_i_10 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[9]_i_3_0 ),
        .I2(\rgf_c1bus_wb[9]_i_3_1 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[1]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hCCCC440C)) 
    \rgf_c1bus_wb[1]_i_12 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[1]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hEFAAEAAA)) 
    \rgf_c1bus_wb[1]_i_15 
       (.I0(\rgf_c1bus_wb[1]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h2A888000)) 
    \rgf_c1bus_wb[1]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(\bdatw[9]_INST_0_i_16_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(a1bus_0[1]),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[1]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[1]_i_18 
       (.I0(\bdatw[9]_INST_0_i_16_n_0 ),
        .I1(\stat_reg[2]_6 ),
        .I2(a1bus_0[1]),
        .O(\rgf_c1bus_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFC0A0CF)) 
    \rgf_c1bus_wb[1]_i_19 
       (.I0(\bdatw[9]_INST_0_i_16_n_0 ),
        .I1(a1bus_0[9]),
        .I2(\stat_reg[1]_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(a1bus_0[1]),
        .I5(\stat_reg[2]_6 ),
        .O(\rgf_c1bus_wb[1]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hFBAA)) 
    \rgf_c1bus_wb[1]_i_2 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_8_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .O(\rgf_c1bus_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000FC54FC)) 
    \rgf_c1bus_wb[1]_i_3 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb_reg[1]_1 ),
        .I5(\rgf_c1bus_wb[1]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h7F55)) 
    \rgf_c1bus_wb[1]_i_5 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(a1bus_0[0]),
        .I3(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c1bus_wb[1]_i_6 
       (.I0(\rgf_c1bus_wb[1]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb_reg[1]_0 ),
        .I2(\rgf_c1bus_wb_reg[3]_2 [1]),
        .I3(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFAFCFAFC0000F000)) 
    \rgf_c1bus_wb[1]_i_7 
       (.I0(\sr[4]_i_43_0 ),
        .I1(\sr[4]_i_43_1 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I5(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[1]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h028A0000)) 
    \rgf_c1bus_wb[1]_i_8 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb[1]_i_2_0 ),
        .I3(\rgf_c1bus_wb[1]_i_2_1 ),
        .I4(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAABABF)) 
    \rgf_c1bus_wb[1]_i_9 
       (.I0(\stat_reg[2]_7 ),
        .I1(\rgf_c1bus_wb[9]_i_3_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[9]_i_3_2 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1110)) 
    \rgf_c1bus_wb[2]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_2_n_0 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\rgf_c1bus_wb[2]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb_reg[2] ),
        .I5(\rgf_c1bus_wb[2]_i_5_n_0 ),
        .O(\bdatr[15] [2]));
  LUT4 #(
    .INIT(16'h1054)) 
    \rgf_c1bus_wb[2]_i_10 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\badr[14]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb_reg[10]_0 ),
        .O(\rgf_c1bus_wb[2]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[2]_i_11 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_33_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[15]_i_4_0 ),
        .O(\rgf_c1bus_wb[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hCCCC440C)) 
    \rgf_c1bus_wb[2]_i_12 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(a1bus_0[1]),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h2A888000)) 
    \rgf_c1bus_wb[2]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(\bdatw[10]_INST_0_i_16_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(a1bus_0[2]),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[2]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[2]_i_15 
       (.I0(\bdatw[10]_INST_0_i_16_n_0 ),
        .I1(\stat_reg[2]_6 ),
        .I2(a1bus_0[2]),
        .O(\rgf_c1bus_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFC0A0CF)) 
    \rgf_c1bus_wb[2]_i_16 
       (.I0(\bdatw[10]_INST_0_i_16_n_0 ),
        .I1(a1bus_0[10]),
        .I2(\stat_reg[1]_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(a1bus_0[2]),
        .I5(\stat_reg[2]_6 ),
        .O(\rgf_c1bus_wb[2]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFDC8C)) 
    \rgf_c1bus_wb[2]_i_17 
       (.I0(\bdatw[8]_INST_0_i_16_1 ),
        .I1(a1bus_0[15]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[14]),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA2022AAAA)) 
    \rgf_c1bus_wb[2]_i_2 
       (.I0(\tr_reg[4]_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(\rgf_c1bus_wb_reg[2]_0 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[2]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFEE0E)) 
    \rgf_c1bus_wb[2]_i_3 
       (.I0(\stat_reg[2]_7 ),
        .I1(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(\rgf_c1bus_wb[2]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEFAAEAAA)) 
    \rgf_c1bus_wb[2]_i_5 
       (.I0(\rgf_c1bus_wb[2]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h777FFF7F)) 
    \rgf_c1bus_wb[2]_i_7 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(\sr[4]_i_45_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\sr[4]_i_34_0 ),
        .O(\rgf_c1bus_wb[2]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[2]_i_8 
       (.I0(\rgf_c1bus_wb[15]_i_14_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_3 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[11]_i_3_0 ),
        .O(\rgf_c1bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0055515100050101)) 
    \rgf_c1bus_wb[2]_i_9 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_44_0 ),
        .I2(\stat_reg[1]_0 ),
        .I3(\rgf_c1bus_wb_reg[10]_0 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\rgf_c1bus_wb[2]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04550400)) 
    \rgf_c1bus_wb[3]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[3] ),
        .I2(\rgf_c1bus_wb[3]_i_3_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\rgf_c1bus_wb[3]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_5_n_0 ),
        .O(\bdatr[15] [3]));
  LUT6 #(
    .INIT(64'h0F0F0B010F0F0F0F)) 
    \rgf_c1bus_wb[3]_i_10 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(a1bus_0[15]),
        .I2(\stat_reg[2]_7 ),
        .I3(\rgf_c1bus_wb_reg[11]_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[3]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h90B02000)) 
    \rgf_c1bus_wb[3]_i_11 
       (.I0(a1bus_0[3]),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h22820082AA828882)) 
    \rgf_c1bus_wb[3]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(a1bus_0[3]),
        .I3(\stat_reg[1]_0 ),
        .I4(a1bus_0[11]),
        .I5(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FFF0777)) 
    \rgf_c1bus_wb[3]_i_13 
       (.I0(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(\stat_reg[2]_6 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(a1bus_0[3]),
        .I5(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFF3FFF3FFF3FC404)) 
    \rgf_c1bus_wb[3]_i_3 
       (.I0(\rgf_c1bus_wb_reg[3]_0 ),
        .I1(\bdatw[9]_INST_0_i_16_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb_reg[3]_1 ),
        .I4(\stat_reg[2]_4 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hC000C0C0C888C8C8)) 
    \rgf_c1bus_wb[3]_i_4 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb_reg[12]_0 ),
        .O(\rgf_c1bus_wb[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFEFFFFFFFE)) 
    \rgf_c1bus_wb[3]_i_5 
       (.I0(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb_reg[3]_3 ),
        .I4(\rgf_c1bus_wb_reg[3]_2 [2]),
        .I5(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[3]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[3]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(a1bus_0[2]),
        .O(\rgf_c1bus_wb[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h10151010FFFFFFFF)) 
    \rgf_c1bus_wb[3]_i_8 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\bdatw[8]_INST_0_i_16_2 ),
        .I4(a1bus_0[15]),
        .I5(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00011101)) 
    \rgf_c1bus_wb[3]_i_9 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\rgf_c1bus_wb[11]_i_6_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb_reg[11]_0 ),
        .O(\rgf_c1bus_wb[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04550400)) 
    \rgf_c1bus_wb[4]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb_reg[4] ),
        .I3(\tr_reg[4]_0 ),
        .I4(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .O(\bdatr[15] [4]));
  LUT5 #(
    .INIT(32'h33BF33B3)) 
    \rgf_c1bus_wb[4]_i_10 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(\stat_reg[1]_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(a1bus_0[3]),
        .O(\rgf_c1bus_wb[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2E222EEE)) 
    \rgf_c1bus_wb[4]_i_11 
       (.I0(\rgf_c1bus_wb[4]_i_22_n_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb[4]_i_4_2 ),
        .I3(\bdatw[8]_INST_0_i_16_1 ),
        .I4(\rgf_c1bus_wb[4]_i_4_3 ),
        .I5(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FDFFFDDD)) 
    \rgf_c1bus_wb[4]_i_13 
       (.I0(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb[4]_i_4_0 ),
        .I3(\bdatw[8]_INST_0_i_16_1 ),
        .I4(\rgf_c1bus_wb[4]_i_4_1 ),
        .I5(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_135 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [4]),
        .O(\sr_reg[0]_31 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_137 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [4]),
        .O(\sr_reg[0]_15 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_139 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [3]),
        .O(\sr_reg[1]_10 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[4]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(a1bus_0[4]),
        .I2(\stat_reg[2]_4 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[4]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_141 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [3]),
        .O(\sr_reg[0]_32 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_143 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [3]),
        .O(\sr_reg[0]_16 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_145 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [2]),
        .O(\sr_reg[0]_33 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_147 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [2]),
        .O(\sr_reg[0]_17 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_149 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [1]),
        .O(\sr_reg[1]_12 ));
  LUT6 #(
    .INIT(64'h22820082AA828882)) 
    \rgf_c1bus_wb[4]_i_15 
       (.I0(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(a1bus_0[4]),
        .I3(\stat_reg[1]_0 ),
        .I4(a1bus_0[12]),
        .I5(\tr_reg[4]_0 ),
        .O(\rgf_c1bus_wb[4]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_151 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [1]),
        .O(\sr_reg[0]_34 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_153 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [1]),
        .O(\sr_reg[0]_18 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_155 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [15]),
        .O(\sr_reg[0]_20 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_157 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [15]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_159 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [13]),
        .O(\sr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h000000000FFF0777)) 
    \rgf_c1bus_wb[4]_i_16 
       (.I0(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(\stat_reg[2]_6 ),
        .I3(\tr_reg[4]_0 ),
        .I4(a1bus_0[4]),
        .I5(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_161 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [14]),
        .O(\sr_reg[0]_21 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_163 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [14]),
        .O(\sr_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_165 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [0]),
        .O(\sr_reg[0]_19 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_167 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [14]),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_169 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [12]),
        .O(\sr_reg[0]_23 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_171 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [12]),
        .O(\sr_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_173 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [13]),
        .O(\sr_reg[0]_22 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_175 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [13]),
        .O(\sr_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_177 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [12]),
        .O(\sr_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_179 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [5]),
        .O(\sr_reg[0]_30 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_181 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [5]),
        .O(\sr_reg[0]_14 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_183 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [5]),
        .O(\sr_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_185 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [6]),
        .O(\sr_reg[0]_29 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_187 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [6]),
        .O(\sr_reg[0]_13 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_189 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [7]),
        .O(\sr_reg[0]_28 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_191 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [7]),
        .O(\sr_reg[0]_12 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_193 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [7]),
        .O(\sr_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_195 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [8]),
        .O(\sr_reg[0]_27 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_197 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [8]),
        .O(\sr_reg[0]_11 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_199 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [9]),
        .O(\sr_reg[0]_26 ));
  LUT6 #(
    .INIT(64'hEAEFEAEAAAAAAAAA)) 
    \rgf_c1bus_wb[4]_i_2 
       (.I0(\stat_reg[2]_8 ),
        .I1(\rgf_c1bus_wb_reg[4]_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\bdatw[8]_INST_0_i_16_2 ),
        .I4(a1bus_0[0]),
        .I5(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_201 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [9]),
        .O(\sr_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_203 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [8]),
        .O(\sr_reg[1]_5 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_205 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [10]),
        .O(\sr_reg[0]_25 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_207 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [10]),
        .O(\sr_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_209 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [11]),
        .O(\sr_reg[0]_24 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \rgf_c1bus_wb[4]_i_211 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_87 [11]),
        .O(\sr_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_213 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [10]),
        .O(\sr_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \rgf_c1bus_wb[4]_i_215 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [2]),
        .O(\sr_reg[1]_11 ));
  LUT6 #(
    .INIT(64'h5555555400000000)) 
    \rgf_c1bus_wb[4]_i_22 
       (.I0(\stat_reg[2]_4 ),
        .I1(\rgf_c1bus_wb[4]_i_11_0 ),
        .I2(a1bus_b02),
        .I3(\rgf_c1bus_wb[4]_i_11_1 ),
        .I4(\rgf_c1bus_wb[4]_i_11_2 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h808880888088AAAA)) 
    \rgf_c1bus_wb[4]_i_4 
       (.I0(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb_reg[4]_0 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\stat_reg[2]_4 ),
        .I5(\rgf_c1bus_wb[4]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFEFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb_reg[4]_2 ),
        .I4(\rgf_c1bus_wb_reg[7]_1 [0]),
        .I5(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40454040)) 
    \rgf_c1bus_wb[5]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\rgf_c1bus_wb[5]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb_reg[5] ),
        .I5(\rgf_c1bus_wb[5]_i_5_n_0 ),
        .O(\bdatr[15] [5]));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c1bus_wb[5]_i_10 
       (.I0(\rgf_c1bus_wb[5]_i_12_n_0 ),
        .I1(\sr[4]_i_53_0 ),
        .I2(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I3(\sr[4]_i_53_1 ),
        .I4(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[5]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(a1bus_0[5]),
        .I2(\stat_reg[2]_4 ),
        .I3(tout__1_carry__0),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[5]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h33100310)) 
    \rgf_c1bus_wb[5]_i_2 
       (.I0(\rgf_c1bus_wb[13]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\stat_reg[2]_8 ),
        .I4(\rgf_c1bus_wb_reg[13]_2 ),
        .O(\rgf_c1bus_wb[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFE040)) 
    \rgf_c1bus_wb[5]_i_3 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(\rgf_c1bus_wb_reg[14]_2 ),
        .I4(\rgf_c1bus_wb[5]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c1bus_wb[5]_i_5 
       (.I0(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[5]_0 ),
        .I2(\rgf_c1bus_wb_reg[7]_1 [1]),
        .I3(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[5]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h1B00)) 
    \rgf_c1bus_wb[5]_i_6 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_43_0 ),
        .I2(\rgf_c1bus_wb[1]_i_2_0 ),
        .I3(\rgf_c1bus_wb[15]_i_14_0 ),
        .O(\rgf_c1bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2A3B6E7FFFFFFFFF)) 
    \rgf_c1bus_wb[5]_i_7 
       (.I0(\bdatw[8]_INST_0_i_16_1 ),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[15]),
        .I3(a1bus_0[14]),
        .I4(a1bus_0[13]),
        .I5(\bdatw[8]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[5]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[5]_i_8 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(a1bus_0[4]),
        .I2(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAABAAAAA)) 
    \rgf_c1bus_wb[5]_i_9 
       (.I0(\stat_reg[2]_4 ),
        .I1(\bdatw[9]_INST_0_i_16_n_0 ),
        .I2(\tr_reg[0] ),
        .I3(\bdatw[10]_INST_0_i_16_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\tr_reg[4]_0 ),
        .O(\stat_reg[2]_7 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4540)) 
    \rgf_c1bus_wb[6]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb_reg[6] ),
        .I5(\rgf_c1bus_wb[6]_i_5_n_0 ),
        .O(\bdatr[15] [6]));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[6]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(a1bus_0[5]),
        .I2(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[6]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFD5D)) 
    \rgf_c1bus_wb[6]_i_11 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[10]_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_33_0 ),
        .O(\rgf_c1bus_wb[6]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_c1bus_wb[6]_i_12 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[6]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[6]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\stat_reg[2]_4 ),
        .I3(\rgf_c1bus_wb[14]_i_3_1 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[6]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[6]_i_16 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[6]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000F350)) 
    \rgf_c1bus_wb[6]_i_2 
       (.I0(\rgf_c1bus_wb_reg[6]_3 ),
        .I1(\rgf_c1bus_wb_reg[6]_2 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\stat_reg[2]_8 ),
        .I4(\rgf_c1bus_wb[6]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h0D0F000F)) 
    \rgf_c1bus_wb[6]_i_3 
       (.I0(\rgf_c1bus_wb[6]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hBFAAAEAA)) 
    \rgf_c1bus_wb[6]_i_5 
       (.I0(\rgf_c1bus_wb[6]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb_reg[6]_0 ),
        .I3(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb_reg[6]_1 ),
        .O(\rgf_c1bus_wb[6]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h08A80000)) 
    \rgf_c1bus_wb[6]_i_7 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_34_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_43_1 ),
        .I4(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[6]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[6]_i_8 
       (.I0(\stat_reg[1]_0 ),
        .I1(\bdatw[9]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAABABF)) 
    \rgf_c1bus_wb[6]_i_9 
       (.I0(\stat_reg[2]_7 ),
        .I1(\sr[4]_i_44_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_46_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45440000)) 
    \rgf_c1bus_wb[7]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .I3(\rgf_c1bus_wb[15]_i_14_0 ),
        .I4(\rgf_c1bus_wb[7]_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .O(\bdatr[15] [7]));
  LUT4 #(
    .INIT(16'hAA8A)) 
    \rgf_c1bus_wb[7]_i_11 
       (.I0(\stat_reg[2]_4 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABABAAABAAAB)) 
    \rgf_c1bus_wb[7]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_14_1 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[15]_i_4_0 ),
        .I4(\rgf_c1bus_wb[11]_i_6_0 ),
        .I5(\bdatw[8]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[7]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0F0FFF2)) 
    \rgf_c1bus_wb[7]_i_13 
       (.I0(\stat_reg[2]_4 ),
        .I1(\rgf_c1bus_wb[15]_i_10_0 ),
        .I2(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c1bus_wb[7]_i_15 
       (.I0(a1bus_0[7]),
        .I1(\rgf_c1bus_wb[15]_i_10_0 ),
        .I2(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[2]_4 ),
        .O(\rgf_c1bus_wb[7]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[7]_i_16 
       (.I0(\stat_reg[2]_4 ),
        .I1(a1bus_0[15]),
        .I2(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[7]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h06FF)) 
    \rgf_c1bus_wb[7]_i_17 
       (.I0(a1bus_0[7]),
        .I1(\stat_reg[2]_4 ),
        .I2(\stat_reg[1]_0 ),
        .I3(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FFF0777)) 
    \rgf_c1bus_wb[7]_i_18 
       (.I0(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I1(\stat_reg[2]_4 ),
        .I2(\stat_reg[2]_6 ),
        .I3(\rgf_c1bus_wb[15]_i_10_0 ),
        .I4(a1bus_0[7]),
        .I5(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h8B00FFFF)) 
    \rgf_c1bus_wb[7]_i_2 
       (.I0(\rgf_c1bus_wb_reg[7]_3 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb_reg[3]_1 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\tr_reg[4]_0 ),
        .O(\rgf_c1bus_wb[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_4 
       (.I0(\stat_reg[2]_8 ),
        .I1(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[15]_i_14_0 ));
  LUT6 #(
    .INIT(64'hABAABBBBABAAABAA)) 
    \rgf_c1bus_wb[7]_i_5 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[7]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb_reg[7]_2 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c1bus_wb[7]_i_6 
       (.I0(\rgf_c1bus_wb[7]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_0 ),
        .I2(\rgf_c1bus_wb_reg[7]_1 [2]),
        .I3(tout__1_carry_i_11_0),
        .O(\rgf_c1bus_wb[7]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[7]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[7]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF54)) 
    \rgf_c1bus_wb[8]_i_1 
       (.I0(\rgf_c1bus_wb[8]_i_2_n_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\rgf_c1bus_wb[8]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[8] ),
        .I4(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .O(\bdatr[15] [8]));
  LUT4 #(
    .INIT(16'h2EFF)) 
    \rgf_c1bus_wb[8]_i_12 
       (.I0(\tr_reg[0] ),
        .I1(\stat_reg[2]_6 ),
        .I2(a1bus_0[8]),
        .I3(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h11111FF1)) 
    \rgf_c1bus_wb[8]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(a1bus_0[8]),
        .I3(\stat_reg[2]_4 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[8]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[8]_i_14 
       (.I0(\stat_reg[2]_4 ),
        .I1(a1bus_0[0]),
        .O(\rgf_c1bus_wb[8]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[8]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(a1bus_0[8]),
        .I2(\stat_reg[2]_4 ),
        .I3(bdatw_8_sn_1),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[8]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[8]_i_16 
       (.I0(\bdatw[10]_INST_0_i_16_n_0 ),
        .I1(\tr_reg[0] ),
        .I2(\bdatw[9]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCFCCCECCCCCCCCCC)) 
    \rgf_c1bus_wb[8]_i_2 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb_reg[8]_1 ),
        .O(\rgf_c1bus_wb[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h80CC8080CCCCCCCC)) 
    \rgf_c1bus_wb[8]_i_3 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb_reg[8]_2 ),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb[15]_i_14_1 ),
        .I5(\rgf_c1bus_wb_reg[8]_0 ),
        .O(\rgf_c1bus_wb[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF57770000)) 
    \rgf_c1bus_wb[8]_i_5 
       (.I0(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA820)) 
    \rgf_c1bus_wb[8]_i_6 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb_reg[4]_1 ),
        .I3(\sr[6]_i_6_1 ),
        .O(\rgf_c1bus_wb[8]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[8]_i_7 
       (.I0(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\stat_reg[2]_8 ),
        .O(\rgf_c1bus_wb[8]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[8]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(a1bus_0[7]),
        .O(\rgf_c1bus_wb[8]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF54)) 
    \rgf_c1bus_wb[9]_i_1 
       (.I0(\rgf_c1bus_wb[9]_i_2_n_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\rgf_c1bus_wb[9]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb_reg[9] ),
        .I4(\rgf_c1bus_wb_reg[9]_i_5_n_0 ),
        .O(\bdatr[15] [9]));
  LUT6 #(
    .INIT(64'hCECEEECCCCCCCCCC)) 
    \rgf_c1bus_wb[9]_i_10 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[15]_i_14_1 ),
        .I2(\rgf_c1bus_wb[9]_i_3_1 ),
        .I3(\rgf_c1bus_wb[9]_i_3_0 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[9]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h8A80AAAA)) 
    \rgf_c1bus_wb[9]_i_11 
       (.I0(\stat_reg[2]_4 ),
        .I1(\rgf_c1bus_wb[9]_i_3_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_29_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .O(\rgf_c1bus_wb[9]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[9]_i_12 
       (.I0(\stat_reg[2]_8 ),
        .I1(a1bus_0[8]),
        .O(\rgf_c1bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h1100011100001000)) 
    \rgf_c1bus_wb[9]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .I3(a1bus_0[9]),
        .I4(\bdatw[9]_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[9]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1151)) 
    \rgf_c1bus_wb[9]_i_14 
       (.I0(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(a1bus_0[1]),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h757F)) 
    \rgf_c1bus_wb[9]_i_15 
       (.I0(\bdatw[8]_INST_0_i_16_1 ),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[15]),
        .O(\rgf_c1bus_wb[9]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h11111FF1)) 
    \rgf_c1bus_wb[9]_i_18 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(a1bus_0[9]),
        .I3(\stat_reg[2]_4 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[9]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hE200)) 
    \rgf_c1bus_wb[9]_i_19 
       (.I0(\bdatw[9]_INST_0_i_16_n_0 ),
        .I1(\stat_reg[2]_6 ),
        .I2(a1bus_0[9]),
        .I3(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hEFAAAAAA)) 
    \rgf_c1bus_wb[9]_i_2 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[9]_0 ),
        .I2(\bdatw[11]_INST_0_i_16_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00FE00FE000000FE)) 
    \rgf_c1bus_wb[9]_i_3 
       (.I0(\rgf_c1bus_wb[9]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEAFBFBFBAAFBBBFB)) 
    \rgf_c1bus_wb[9]_i_7 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I3(\stat_reg[2]_8 ),
        .I4(\rgf_c1bus_wb[1]_i_2_0 ),
        .I5(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00022202)) 
    \rgf_c1bus_wb[9]_i_8 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\rgf_c1bus_wb[9]_i_3_2 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[9]_i_3_1 ),
        .O(\rgf_c1bus_wb[9]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000027)) 
    \rgf_c1bus_wb[9]_i_9 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[0]_i_4_0 ),
        .I2(\sr[4]_i_39_0 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\stat_reg[1]_0 ),
        .O(\rgf_c1bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[11]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_20_n_0 ),
        .O(\rgf_c1bus_wb_reg[11]_i_7_n_0 ),
        .S(\rgf_c1bus_wb[14]_i_12_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[12]_i_15 
       (.I0(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_23_n_0 ),
        .O(\rgf_c1bus_wb_reg[12]_i_15_n_0 ),
        .S(\rgf_c1bus_wb[14]_i_12_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[9]_i_5 
       (.I0(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .O(\rgf_c1bus_wb_reg[9]_i_5_n_0 ),
        .S(\rgf_c1bus_wb[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hD500D5D5D500D500)) 
    \rgf_selc0_rn_wb[0]_i_1 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_4_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_5_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0]_0 ),
        .O(\stat_reg[2] [0]));
  LUT6 #(
    .INIT(64'h000D0000000D000D)) 
    \rgf_selc0_rn_wb[0]_i_10 
       (.I0(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_19_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_20_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAAAAA)) 
    \rgf_selc0_rn_wb[0]_i_11 
       (.I0(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_23_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(ir0[15]),
        .I4(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(\rgf_selc0_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0031001100110011)) 
    \rgf_selc0_rn_wb[0]_i_12 
       (.I0(\rgf_selc0_rn_wb[0]_i_24_n_0 ),
        .I1(rst_n_fl_reg_2),
        .I2(ir0[12]),
        .I3(\ccmd[4]_INST_0_i_20_n_0 ),
        .I4(ir0[11]),
        .I5(\rgf_selc0_rn_wb[0]_i_25_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hDD0DFF0FDD0D0000)) 
    \rgf_selc0_rn_wb[0]_i_13 
       (.I0(ir0[10]),
        .I1(\rgf_selc0_rn_wb[0]_i_26_n_0 ),
        .I2(ir0[3]),
        .I3(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I4(ir0[11]),
        .I5(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0111100010000111)) 
    \rgf_selc0_rn_wb[0]_i_14 
       (.I0(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(\sr_reg[15]_0 [7]),
        .I4(\sr_reg[15]_0 [5]),
        .I5(ir0[11]),
        .O(\rgf_selc0_rn_wb[0]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h08888888)) 
    \rgf_selc0_rn_wb[0]_i_15 
       (.I0(ir0[8]),
        .I1(ir0[15]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .I4(ir0[13]),
        .O(\rgf_selc0_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00008808AAAAAAAA)) 
    \rgf_selc0_rn_wb[0]_i_16 
       (.I0(\ccmd[0]_INST_0_i_11_n_0 ),
        .I1(ir0[11]),
        .I2(ir0[12]),
        .I3(\sr_reg[15]_0 [4]),
        .I4(ir0[13]),
        .I5(\rgf_selc0_rn_wb[0]_i_5_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h5F1F5F1F00005F1F)) 
    \rgf_selc0_rn_wb[0]_i_17 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(ir0[10]),
        .I2(ir0[3]),
        .I3(\stat[0]_i_17_n_0 ),
        .I4(\ccmd[4]_INST_0_i_18_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_29_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0200000003F003F0)) 
    \rgf_selc0_rn_wb[0]_i_18 
       (.I0(\rgf_selc0_rn_wb[0]_i_30_n_0 ),
        .I1(crdy),
        .I2(ir0[11]),
        .I3(ir0[10]),
        .I4(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_31_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8000C0C080000000)) 
    \rgf_selc0_rn_wb[0]_i_19 
       (.I0(ir0[3]),
        .I1(\rgf_selc0_rn_wb[0]_i_32_n_0 ),
        .I2(\stat[0]_i_7_n_0 ),
        .I3(crdy),
        .I4(ir0[7]),
        .I5(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \rgf_selc0_rn_wb[0]_i_2 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h3FFFFFFFFFFFBBBB)) 
    \rgf_selc0_rn_wb[0]_i_20 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(brdy),
        .I3(ir0[0]),
        .I4(ir0[6]),
        .I5(ir0[5]),
        .O(\rgf_selc0_rn_wb[0]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \rgf_selc0_rn_wb[0]_i_21 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .O(\rgf_selc0_rn_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0020220000202000)) 
    \rgf_selc0_rn_wb[0]_i_22 
       (.I0(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .I1(ir0[0]),
        .I2(ir0[2]),
        .I3(ir0[1]),
        .I4(ir0[3]),
        .I5(brdy),
        .O(\rgf_selc0_rn_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h000C00C000002F00)) 
    \rgf_selc0_rn_wb[0]_i_23 
       (.I0(brdy),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ir0[3]),
        .I5(ir0[2]),
        .O(\rgf_selc0_rn_wb[0]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFDFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_24 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .I2(ir0[0]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA00000C000000)) 
    \rgf_selc0_rn_wb[0]_i_25 
       (.I0(ir0[0]),
        .I1(ir0[3]),
        .I2(ir0[6]),
        .I3(brdy),
        .I4(ir0[7]),
        .I5(ir0[8]),
        .O(\rgf_selc0_rn_wb[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFFFFFAFAF33F3)) 
    \rgf_selc0_rn_wb[0]_i_26 
       (.I0(\rgf_selc0_rn_wb[0]_i_33_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[9]),
        .I5(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF77FFFF5F)) 
    \rgf_selc0_rn_wb[0]_i_27 
       (.I0(ir0[3]),
        .I1(ir0[6]),
        .I2(crdy),
        .I3(ir0[7]),
        .I4(ir0[8]),
        .I5(\ccmd[4]_INST_0_i_20_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[0]_i_28 
       (.I0(ir0[15]),
        .I1(ir0[14]),
        .O(\rgf_selc0_rn_wb[0]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_selc0_rn_wb[0]_i_29 
       (.I0(ir0[3]),
        .I1(ir0[7]),
        .I2(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc0_rn_wb[0]_i_3 
       (.I0(ir0[3]),
        .I1(ir0[0]),
        .I2(ir0[1]),
        .I3(ir0[2]),
        .O(\rgf_selc0_rn_wb[0]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_30 
       (.I0(ir0[0]),
        .I1(ir0[7]),
        .O(\rgf_selc0_rn_wb[0]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hDFFFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_31 
       (.I0(brdy),
        .I1(ir0[6]),
        .I2(ir0[9]),
        .I3(ir0[8]),
        .I4(ir0[3]),
        .O(\rgf_selc0_rn_wb[0]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_32 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .O(\rgf_selc0_rn_wb[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hEFFF33FAFFFFFFFB)) 
    \rgf_selc0_rn_wb[0]_i_33 
       (.I0(ir0[3]),
        .I1(ir0[7]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(ir0[0]),
        .O(\rgf_selc0_rn_wb[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_selc0_rn_wb[0]_i_4 
       (.I0(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0]_1 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\rgf_selc0_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000000000E000E0E)) 
    \rgf_selc0_rn_wb[0]_i_5 
       (.I0(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_12_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_15_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc0_rn_wb[0]_i_6 
       (.I0(ir0[7]),
        .I1(ir0[5]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .O(\rgf_selc0_rn_wb[0]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[0]_i_7 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .O(\rgf_selc0_rn_wb[0]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[0]_i_8 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\rgf_selc0_rn_wb[0]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc0_rn_wb[0]_i_9 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[15]),
        .I3(ir0[14]),
        .O(\rgf_selc0_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0055005700550055)) 
    \rgf_selc0_rn_wb[1]_i_1 
       (.I0(\rgf_selc0_rn_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(\rgf_selc0_rn_wb_reg[0] [2]),
        .I4(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .O(\stat_reg[2] [1]));
  LUT4 #(
    .INIT(16'h0440)) 
    \rgf_selc0_rn_wb[1]_i_10 
       (.I0(ir0[0]),
        .I1(ir0[2]),
        .I2(ir0[1]),
        .I3(ir0[3]),
        .O(\rgf_selc0_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \rgf_selc0_rn_wb[1]_i_11 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[9]),
        .I3(\rgf_selc0_rn_wb[2]_i_12_n_0 ),
        .I4(ir0[15]),
        .I5(\bcmd[0]_INST_0_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[1]_i_12 
       (.I0(crdy),
        .I1(ir0[11]),
        .O(\rgf_selc0_rn_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hE0E04040FFE04040)) 
    \rgf_selc0_rn_wb[1]_i_13 
       (.I0(ir0[7]),
        .I1(ir0[1]),
        .I2(\ccmd[4]_INST_0_i_18_n_0 ),
        .I3(ir0[10]),
        .I4(ir0[4]),
        .I5(\stat[0]_i_17_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF04FF04FF04FF)) 
    \rgf_selc0_rn_wb[1]_i_14 
       (.I0(\rgf_selc0_rn_wb[1]_i_22_n_0 ),
        .I1(ir0[1]),
        .I2(ir0[7]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\rgf_selc0_rn_wb[1]_i_23_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_24_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA808880888088)) 
    \rgf_selc0_rn_wb[1]_i_15 
       (.I0(\stat[0]_i_7_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_25_n_0 ),
        .I2(crdy),
        .I3(ir0[7]),
        .I4(\bdatw[10]_INST_0_i_18_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_19_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h8A88888888888888)) 
    \rgf_selc0_rn_wb[1]_i_16 
       (.I0(\stat[0]_i_7_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_26_n_0 ),
        .I2(ir0[5]),
        .I3(\rgf_selc0_rn_wb[1]_i_27_n_0 ),
        .I4(ir0[1]),
        .I5(\stat[2]_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \rgf_selc0_rn_wb[1]_i_17 
       (.I0(crdy),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .O(\rgf_selc0_rn_wb[1]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h40000000)) 
    \rgf_selc0_rn_wb[1]_i_18 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .I3(ir0[8]),
        .I4(ir0[7]),
        .O(\rgf_selc0_rn_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8AAAAAAAAA8AAA8A)) 
    \rgf_selc0_rn_wb[1]_i_19 
       (.I0(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I1(\ccmd[4]_INST_0_i_20_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I3(ir0[7]),
        .I4(ir0[6]),
        .I5(ir0[8]),
        .O(\rgf_selc0_rn_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000000BFFBBFF)) 
    \rgf_selc0_rn_wb[1]_i_2 
       (.I0(\rgf_selc0_rn_wb[1]_i_6_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0]_1 ),
        .I4(\rgf_selc0_rn_wb[1]_i_10_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_11_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h80808C8080808080)) 
    \rgf_selc0_rn_wb[1]_i_20 
       (.I0(ir0[1]),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(brdy),
        .I4(ir0[6]),
        .I5(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF040004)) 
    \rgf_selc0_rn_wb[1]_i_21 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(\ccmd[4]_INST_0_i_20_n_0 ),
        .I3(\ccmd[4]_INST_0_i_12_n_0 ),
        .I4(crdy),
        .I5(ir0[11]),
        .O(\rgf_selc0_rn_wb[1]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \rgf_selc0_rn_wb[1]_i_22 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[10]),
        .I3(ir0[11]),
        .I4(crdy),
        .O(\rgf_selc0_rn_wb[1]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h08000000)) 
    \rgf_selc0_rn_wb[1]_i_23 
       (.I0(ir0[4]),
        .I1(brdy),
        .I2(ir0[6]),
        .I3(ir0[9]),
        .I4(ir0[8]),
        .O(\rgf_selc0_rn_wb[1]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h46)) 
    \rgf_selc0_rn_wb[1]_i_24 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(crdy),
        .O(\rgf_selc0_rn_wb[1]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    \rgf_selc0_rn_wb[1]_i_25 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[1]),
        .I3(ir0[7]),
        .I4(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000404000FF)) 
    \rgf_selc0_rn_wb[1]_i_26 
       (.I0(\rgf_selc0_rn_wb[1]_i_28_n_0 ),
        .I1(ir0[8]),
        .I2(\bcmd[0]_INST_0_i_21_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_29_n_0 ),
        .I4(ir0[9]),
        .I5(ir0[7]),
        .O(\rgf_selc0_rn_wb[1]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_rn_wb[1]_i_27 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .O(\rgf_selc0_rn_wb[1]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \rgf_selc0_rn_wb[1]_i_28 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[4]),
        .O(\rgf_selc0_rn_wb[1]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \rgf_selc0_rn_wb[1]_i_29 
       (.I0(ir0[4]),
        .I1(ir0[8]),
        .I2(crdy),
        .O(\rgf_selc0_rn_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000557F)) 
    \rgf_selc0_rn_wb[1]_i_3 
       (.I0(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I1(\ccmd[4]_INST_0_i_12_n_0 ),
        .I2(ir0[4]),
        .I3(\rgf_selc0_rn_wb[1]_i_13_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_14_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \rgf_selc0_rn_wb[1]_i_4 
       (.I0(ir0[12]),
        .I1(ir0[13]),
        .I2(ir0[14]),
        .I3(ir0[15]),
        .O(\rgf_selc0_rn_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEFEEEFFFFFEEE)) 
    \rgf_selc0_rn_wb[1]_i_5 
       (.I0(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I4(ir0[4]),
        .I5(\rgf_selc0_rn_wb[1]_i_19_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000F7F7F7F7F7)) 
    \rgf_selc0_rn_wb[1]_i_6 
       (.I0(\rgf_selc0_rn_wb[1]_i_20_n_0 ),
        .I1(ir0[11]),
        .I2(\ccmd[4]_INST_0_i_20_n_0 ),
        .I3(ir0[1]),
        .I4(\ccmd[4]_INST_0_i_12_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc0_rn_wb[1]_i_7 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\rgf_selc0_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \rgf_selc0_rn_wb[1]_i_8 
       (.I0(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_18_n_0 ),
        .I3(ir0[4]),
        .I4(ir0[6]),
        .I5(\ccmd[4]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000075FF7575)) 
    \rgf_selc0_rn_wb[2]_i_1 
       (.I0(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I5(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(\stat_reg[2] [2]));
  LUT4 #(
    .INIT(16'h6000)) 
    \rgf_selc0_rn_wb[2]_i_10 
       (.I0(ir0[10]),
        .I1(ir0[11]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .O(\rgf_selc0_rn_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEEEEEEEEEEEEE)) 
    \rgf_selc0_rn_wb[2]_i_11 
       (.I0(\rgf_selc0_rn_wb[2]_i_17_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_18_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_19_n_0 ),
        .I3(\stat[0]_i_7_n_0 ),
        .I4(ir0[3]),
        .I5(ir0[2]),
        .O(\rgf_selc0_rn_wb[2]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_selc0_rn_wb[2]_i_12 
       (.I0(ir0[11]),
        .I1(ir0[13]),
        .I2(ir0[12]),
        .I3(ir0[14]),
        .O(\rgf_selc0_rn_wb[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hD555FFFF)) 
    \rgf_selc0_rn_wb[2]_i_13 
       (.I0(ir0[15]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(ir0[13]),
        .I4(ir0[10]),
        .O(\rgf_selc0_rn_wb[2]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFE0FFFF)) 
    \rgf_selc0_rn_wb[2]_i_14 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[11]),
        .O(\rgf_selc0_rn_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hE0EEE0E0E0E0E0E0)) 
    \rgf_selc0_rn_wb[2]_i_15 
       (.I0(\rgf_selc0_rn_wb[2]_i_20_n_0 ),
        .I1(\stat[0]_i_7_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_21_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_22_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_23_n_0 ),
        .I5(ir0[9]),
        .O(\rgf_selc0_rn_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \rgf_selc0_rn_wb[2]_i_16 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(brdy),
        .I5(\ccmd[4]_INST_0_i_20_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h3370007000500050)) 
    \rgf_selc0_rn_wb[2]_i_17 
       (.I0(\rgf_selc0_rn_wb[1]_i_22_n_0 ),
        .I1(\stat[0]_i_16_n_0 ),
        .I2(ir0[2]),
        .I3(ir0[7]),
        .I4(ir0[5]),
        .I5(\badr[15]_INST_0_i_205_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hA000C0000000C000)) 
    \rgf_selc0_rn_wb[2]_i_18 
       (.I0(ir0[5]),
        .I1(ir0[2]),
        .I2(ir0[8]),
        .I3(\bdatw[15]_INST_0_i_61_n_0 ),
        .I4(ir0[7]),
        .I5(crdy),
        .O(\rgf_selc0_rn_wb[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \rgf_selc0_rn_wb[2]_i_19 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .I3(brdy),
        .I4(ir0[5]),
        .I5(ir0[7]),
        .O(\rgf_selc0_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0007)) 
    \rgf_selc0_rn_wb[2]_i_2 
       (.I0(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[11]),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4040100000001000)) 
    \rgf_selc0_rn_wb[2]_i_20 
       (.I0(\ccmd[4]_INST_0_i_20_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(crdy),
        .I4(ir0[8]),
        .I5(ir0[6]),
        .O(\rgf_selc0_rn_wb[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h030B0300FFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_21 
       (.I0(crdy),
        .I1(ir0[8]),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(ir0[5]),
        .I5(ir0[11]),
        .O(\rgf_selc0_rn_wb[2]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hF0FFDFFE)) 
    \rgf_selc0_rn_wb[2]_i_22 
       (.I0(ir0[4]),
        .I1(ir0[3]),
        .I2(ir0[5]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .O(\rgf_selc0_rn_wb[2]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_rn_wb[2]_i_23 
       (.I0(ir0[8]),
        .I1(ir0[2]),
        .O(\rgf_selc0_rn_wb[2]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555F7FF)) 
    \rgf_selc0_rn_wb[2]_i_3 
       (.I0(ir0[5]),
        .I1(brdy),
        .I2(ir0[6]),
        .I3(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I4(\ccmd[3]_INST_0_i_14_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_selc0_rn_wb[2]_i_4 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[12]),
        .I3(ir0[15]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\rgf_selc0_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEE0000EE0E)) 
    \rgf_selc0_rn_wb[2]_i_5 
       (.I0(\rgf_selc0_rn_wb[2]_i_12_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_13_n_0 ),
        .I2(ir0[5]),
        .I3(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_15_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \rgf_selc0_rn_wb[2]_i_7 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .O(\rgf_selc0_rn_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF7F0000)) 
    \rgf_selc0_rn_wb[2]_i_8 
       (.I0(ir0[8]),
        .I1(ir0[2]),
        .I2(ir0[7]),
        .I3(\ccmd[4]_INST_0_i_20_n_0 ),
        .I4(ir0[11]),
        .I5(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_9 
       (.I0(ir0[15]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[12]),
        .I4(ir0[14]),
        .I5(ir0[13]),
        .O(\rgf_selc0_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc0_stat_i_2
       (.I0(\stat_reg[2]_0 [1]),
        .I1(\stat_reg[2]_0 [0]),
        .O(E));
  LUT6 #(
    .INIT(64'h4445444455555555)) 
    \rgf_selc0_wb[0]_i_1 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_4_n_0 ),
        .I4(\rgf_selc0_wb[0]_i_5_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_6_n_0 ),
        .O(\stat_reg[2]_0 [0]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[0]_i_10 
       (.I0(ir0[11]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\rgf_selc0_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hC00AFFFFC00A0000)) 
    \rgf_selc0_wb[0]_i_11 
       (.I0(\rgf_selc0_rn_wb[1]_i_27_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_16_n_0 ),
        .I2(ir0[9]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[8]),
        .I5(\rgf_selc0_wb[0]_i_17_n_0 ),
        .O(\rgf_selc0_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h88880080888822A2)) 
    \rgf_selc0_wb[0]_i_12 
       (.I0(\ccmd[0]_INST_0_i_17_n_0 ),
        .I1(ir0[11]),
        .I2(brdy),
        .I3(ir0[6]),
        .I4(ir0[8]),
        .I5(\ccmd[4]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h7F7FF0F05757F0FF)) 
    \rgf_selc0_wb[0]_i_13 
       (.I0(ir0[8]),
        .I1(crdy),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[6]),
        .I4(ir0[10]),
        .I5(ir0[7]),
        .O(\rgf_selc0_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF7FF77FFF7FF)) 
    \rgf_selc0_wb[0]_i_14 
       (.I0(ir0[8]),
        .I1(brdy),
        .I2(ir0[10]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[6]),
        .I5(ir0[4]),
        .O(\rgf_selc0_wb[0]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hAAA8)) 
    \rgf_selc0_wb[0]_i_15 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .O(\rgf_selc0_wb[0]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[0]_i_16 
       (.I0(brdy),
        .I1(ir0[6]),
        .O(\rgf_selc0_wb[0]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h4504)) 
    \rgf_selc0_wb[0]_i_17 
       (.I0(ir0[9]),
        .I1(crdy),
        .I2(ir0[7]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\rgf_selc0_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h282200008AAA0000)) 
    \rgf_selc0_wb[0]_i_2 
       (.I0(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .I4(ir0[15]),
        .I5(ir0[14]),
        .O(\rgf_selc0_wb[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h8888888F)) 
    \rgf_selc0_wb[0]_i_3 
       (.I0(ir0[1]),
        .I1(ir0[3]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(crdy),
        .O(\rgf_selc0_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    \rgf_selc0_wb[0]_i_4 
       (.I0(ir0[2]),
        .I1(ir0[0]),
        .I2(\ccmd[4]_INST_0_i_13_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I4(ir0[9]),
        .I5(ir0[4]),
        .O(\rgf_selc0_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \rgf_selc0_wb[0]_i_5 
       (.I0(\bcmd[0]_INST_0_i_19_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[7]),
        .I3(\ccmd[0]_INST_0_i_11_n_0 ),
        .I4(ir0[13]),
        .I5(ir0[12]),
        .O(\rgf_selc0_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBABBBBBBBB)) 
    \rgf_selc0_wb[0]_i_6 
       (.I0(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_7_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_9_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(ir0[11]),
        .O(\rgf_selc0_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF404040)) 
    \rgf_selc0_wb[0]_i_7 
       (.I0(\rgf_selc0_wb[0]_i_10_n_0 ),
        .I1(ir0[10]),
        .I2(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I3(\ccmd[3]_INST_0_i_14_n_0 ),
        .I4(\ccmd[2]_INST_0_i_3_0 ),
        .I5(\rgf_selc0_wb[0]_i_12_n_0 ),
        .O(\rgf_selc0_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000AAA80200AAA8)) 
    \rgf_selc0_wb[0]_i_8 
       (.I0(\rgf_selc0_wb[0]_i_13_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[9]),
        .I5(ir0[10]),
        .O(\rgf_selc0_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFB00FBFB00000000)) 
    \rgf_selc0_wb[0]_i_9 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\ccmd[1]_INST_0_i_18_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_22_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I4(\stat[0]_i_25_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_15_n_0 ),
        .O(\rgf_selc0_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00F1FFFF00F100F1)) 
    \rgf_selc0_wb[1]_i_1 
       (.I0(\rgf_selc0_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_4_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [2]),
        .I4(\rgf_selc0_wb[1]_i_5_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_6_n_0 ),
        .O(\stat_reg[2]_0 [1]));
  LUT5 #(
    .INIT(32'h70000000)) 
    \rgf_selc0_wb[1]_i_10 
       (.I0(\stat[0]_i_25_n_0 ),
        .I1(\stat[0]_i_27_n_0 ),
        .I2(ir0[11]),
        .I3(ir0[9]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\rgf_selc0_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AA8AAAAA)) 
    \rgf_selc0_wb[1]_i_11 
       (.I0(\rgf_selc0_wb[1]_i_20_n_0 ),
        .I1(ir0[9]),
        .I2(ir0[7]),
        .I3(ir0[11]),
        .I4(ir0[6]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\rgf_selc0_wb[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_selc0_wb[1]_i_12 
       (.I0(ir0[10]),
        .I1(ir0[9]),
        .I2(ir0[8]),
        .O(\rgf_selc0_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFAFBFF0F)) 
    \rgf_selc0_wb[1]_i_13 
       (.I0(ir0[9]),
        .I1(crdy),
        .I2(ir0[11]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[10]),
        .I5(ir0[7]),
        .O(\rgf_selc0_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCECECCCCCECEFCCF)) 
    \rgf_selc0_wb[1]_i_14 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_21_n_0 ),
        .I2(ir0[11]),
        .I3(\rgf_selc0_wb[1]_i_22_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(ir0[14]),
        .O(\rgf_selc0_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FFFFFFB0)) 
    \rgf_selc0_wb[1]_i_15 
       (.I0(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_24_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_4_1 ),
        .I3(\rgf_selc0_wb[1]_i_26_n_0 ),
        .I4(ir0[15]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\rgf_selc0_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFF5F00C000550000)) 
    \rgf_selc0_wb[1]_i_16 
       (.I0(\rgf_selc0_wb[1]_i_4_0 ),
        .I1(\sr_reg[15]_0 [6]),
        .I2(ir0[11]),
        .I3(ir0[14]),
        .I4(ir0[15]),
        .I5(\ccmd[0]_INST_0_i_1_0 ),
        .O(\rgf_selc0_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h5555554555555555)) 
    \rgf_selc0_wb[1]_i_17 
       (.I0(\rgf_selc0_wb[1]_i_28_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_29_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I3(ir0[11]),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\ccmd[4]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_wb[1]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc0_wb[1]_i_18 
       (.I0(ir0[15]),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .O(\rgf_selc0_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABABABABABABA)) 
    \rgf_selc0_wb[1]_i_19 
       (.I0(\rgf_selc0_wb[1]_i_30_n_0 ),
        .I1(ir0[11]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[6]),
        .I4(ir0[10]),
        .I5(ir0[9]),
        .O(\rgf_selc0_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h37FF35FFFFFFFFFF)) 
    \rgf_selc0_wb[1]_i_2 
       (.I0(\rgf_selc0_wb[1]_i_7_n_0 ),
        .I1(ir0[12]),
        .I2(ir0[14]),
        .I3(\rgf_selc0_wb[1]_i_8_n_0 ),
        .I4(\sr_reg[15]_0 [6]),
        .I5(ir0[13]),
        .O(\rgf_selc0_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFF5DFFF555DFFFD)) 
    \rgf_selc0_wb[1]_i_20 
       (.I0(\stat[0]_i_23__0_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[4]),
        .I3(ir0[6]),
        .I4(ir0[7]),
        .I5(ir0[5]),
        .O(\rgf_selc0_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00040000000F0000)) 
    \rgf_selc0_wb[1]_i_21 
       (.I0(ir0[7]),
        .I1(crdy),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[9]),
        .I4(ir0[11]),
        .I5(\ccmd[1]_INST_0_i_18_n_0 ),
        .O(\rgf_selc0_wb[1]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_wb[1]_i_22 
       (.I0(ir0[12]),
        .I1(\sr_reg[15]_0 [7]),
        .O(\rgf_selc0_wb[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \rgf_selc0_wb[1]_i_23 
       (.I0(ir0[2]),
        .I1(\ccmd[1]_INST_0_i_10_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_31_n_0 ),
        .I3(\bcmd[0]_INST_0_i_22_n_0 ),
        .I4(ir0[0]),
        .I5(ir0[14]),
        .O(\rgf_selc0_wb[1]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0451)) 
    \rgf_selc0_wb[1]_i_24 
       (.I0(ir0[12]),
        .I1(ir0[14]),
        .I2(\sr_reg[15]_0 [5]),
        .I3(ir0[11]),
        .O(\rgf_selc0_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h082008A008000880)) 
    \rgf_selc0_wb[1]_i_26 
       (.I0(\rgf_selc0_wb[1]_i_32_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[1]),
        .I3(ir0[3]),
        .I4(ir0[0]),
        .I5(brdy),
        .O(\rgf_selc0_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h4044404040404040)) 
    \rgf_selc0_wb[1]_i_28 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .I3(\ccmd[4]_INST_0_i_20_n_0 ),
        .I4(ir0[7]),
        .I5(\rgf_selc0_wb[1]_i_33_n_0 ),
        .O(\rgf_selc0_wb[1]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAA55F300FFFF)) 
    \rgf_selc0_wb[1]_i_29 
       (.I0(ir0[3]),
        .I1(brdy),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[1]),
        .I4(ir0[0]),
        .I5(ir0[2]),
        .O(\rgf_selc0_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFE00FE)) 
    \rgf_selc0_wb[1]_i_3 
       (.I0(\rgf_selc0_wb[1]_i_9_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_10_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_11_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_12_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_13_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_14_n_0 ),
        .O(\rgf_selc0_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7000000)) 
    \rgf_selc0_wb[1]_i_30 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .I2(ir0[5]),
        .I3(ir0[9]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(brdy),
        .O(\rgf_selc0_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \rgf_selc0_wb[1]_i_31 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(ir0[8]),
        .I3(crdy),
        .I4(ir0[9]),
        .I5(ir0[10]),
        .O(\rgf_selc0_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf_selc0_wb[1]_i_32 
       (.I0(ir0[9]),
        .I1(\bdatw[15]_INST_0_i_19_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(ir0[11]),
        .I5(\rgf_selc0_wb[1]_i_34_n_0 ),
        .O(\rgf_selc0_wb[1]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hAA08)) 
    \rgf_selc0_wb[1]_i_33 
       (.I0(ir0[11]),
        .I1(brdy),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .O(\rgf_selc0_wb[1]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc0_wb[1]_i_34 
       (.I0(ir0[5]),
        .I1(ir0[4]),
        .I2(ir0[6]),
        .I3(ir0[8]),
        .I4(ir0[10]),
        .I5(ir0[7]),
        .O(\rgf_selc0_wb[1]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0F4F4F0FFF4F4)) 
    \rgf_selc0_wb[1]_i_4 
       (.I0(ir0[13]),
        .I1(\rgf_selc0_wb[1]_i_15_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I3(ir0[15]),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(\rgf_selc0_wb[1]_i_17_n_0 ),
        .O(\rgf_selc0_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFFFF)) 
    \rgf_selc0_wb[1]_i_5 
       (.I0(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I1(\ccmd[1]_INST_0_i_9_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I3(\rgf_selc0_rn_wb_reg[0] [2]),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\rgf_selc0_wb[1]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \rgf_selc0_wb[1]_i_6 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(\rgf_selc0_wb[1]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h4015)) 
    \rgf_selc0_wb[1]_i_7 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[12]),
        .I2(\sr_reg[15]_0 [7]),
        .I3(ir0[11]),
        .O(\rgf_selc0_wb[1]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_wb[1]_i_8 
       (.I0(ir0[15]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\rgf_selc0_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000E00)) 
    \rgf_selc0_wb[1]_i_9 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\ccmd[4]_INST_0_i_12_n_0 ),
        .I2(ir0[9]),
        .I3(ir0[7]),
        .I4(crdy),
        .I5(\rgf_selc0_wb[1]_i_19_n_0 ),
        .O(\rgf_selc0_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5555100055555555)) 
    \rgf_selc1_rn_wb[0]_i_1 
       (.I0(\rgf_selc1_rn_wb_reg[0] ),
        .I1(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I2(\rgf_selc1_wb_reg[1]_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\stat_reg[2]_1 [0]));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[0]_i_10 
       (.I0(ir1[9]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .O(\rgf_selc1_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \rgf_selc1_rn_wb[0]_i_11 
       (.I0(ir1[8]),
        .I1(\rgf_selc1_rn_wb[1]_i_9_n_0 ),
        .I2(ir1[0]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(ir1[10]),
        .O(\rgf_selc1_rn_wb[0]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc1_rn_wb[0]_i_12 
       (.I0(ir1[12]),
        .I1(ir1[13]),
        .I2(ir1[14]),
        .O(\rgf_selc1_rn_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040F00000)) 
    \rgf_selc1_rn_wb[0]_i_13 
       (.I0(\stat_reg[0]_48 ),
        .I1(brdy),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hEF00EFEF00000000)) 
    \rgf_selc1_rn_wb[0]_i_14 
       (.I0(\rgf_selc1_rn_wb[0]_i_21_n_0 ),
        .I1(ir1[15]),
        .I2(ir1[14]),
        .I3(\rgf_selc1_rn_wb[2]_i_7_n_0 ),
        .I4(ir1[8]),
        .I5(\sr_reg[4] ),
        .O(\rgf_selc1_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF00FFDFF)) 
    \rgf_selc1_rn_wb[0]_i_15 
       (.I0(brdy),
        .I1(\stat_reg[0]_48 ),
        .I2(ir1[3]),
        .I3(ir1[1]),
        .I4(ir1[2]),
        .I5(ir1[0]),
        .O(\rgf_selc1_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_16 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_rn_wb[0]_i_22_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I3(ir1[8]),
        .I4(ir1[7]),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_selc1_rn_wb[0]_i_17 
       (.I0(ir1[0]),
        .I1(ir1[3]),
        .I2(ir1[7]),
        .O(\rgf_selc1_rn_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hD5DDDDDDDDDDDDDD)) 
    \rgf_selc1_rn_wb[0]_i_18 
       (.I0(\rgf_selc1_rn_wb[0]_i_24_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .I2(\stat_reg[0]_48 ),
        .I3(brdy),
        .I4(\rgf_selc1_rn_wb[0]_i_26_n_0 ),
        .I5(\bdatw[11]_INST_0_i_28_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h33337FFF00005555)) 
    \rgf_selc1_rn_wb[0]_i_19 
       (.I0(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I1(ir1[3]),
        .I2(\stat_reg[0]_55 ),
        .I3(\rgf_selc1_wb[0]_i_18_n_0 ),
        .I4(rst_n_fl_reg_9),
        .I5(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_20 
       (.I0(ir1[3]),
        .I1(ir1[2]),
        .O(\rgf_selc1_rn_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hA200A2A2AAAAAAAA)) 
    \rgf_selc1_rn_wb[0]_i_21 
       (.I0(\stat[1]_i_6__0_n_0 ),
        .I1(ir1[3]),
        .I2(\rgf_selc1_rn_wb[1]_i_21_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_28_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc1_rn_wb[0]_i_22 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[15]),
        .I3(ir1[14]),
        .O(\rgf_selc1_rn_wb[0]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_23 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\rgf_selc1_rn_wb[0]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc1_rn_wb[0]_i_24 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .O(\rgf_selc1_rn_wb[0]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \rgf_selc1_rn_wb[0]_i_25 
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .O(\rgf_selc1_rn_wb[0]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[0]_i_26 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .O(\rgf_selc1_rn_wb[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF27FFFFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_27 
       (.I0(ir1[7]),
        .I1(ir1[3]),
        .I2(ir1[0]),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .I5(\bdatw[15]_INST_0_i_197_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h70FFFFFF77FFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_28 
       (.I0(ir1[7]),
        .I1(\rgf_selc1_rn_wb[0]_i_29_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_20_n_0 ),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .I5(ir1[0]),
        .O(\rgf_selc1_rn_wb[0]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc1_rn_wb[0]_i_29 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .I2(ir1[3]),
        .I3(ir1[4]),
        .O(\rgf_selc1_rn_wb[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAAA882AAAAAAAAAA)) 
    \rgf_selc1_rn_wb[0]_i_3 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .I3(ir1[2]),
        .I4(ir1[0]),
        .I5(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF800)) 
    \rgf_selc1_rn_wb[0]_i_5 
       (.I0(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_11_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_13_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_rn_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCCCDDCCCFCCDD)) 
    \rgf_selc1_rn_wb[0]_i_6 
       (.I0(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF7550000FFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_7 
       (.I0(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_17_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_18_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf_selc1_rn_wb[0]_i_8 
       (.I0(ir1[14]),
        .I1(ir1[12]),
        .I2(\bcmd[0]_INST_0_i_14_n_0 ),
        .I3(\bcmd[0]_INST_0_i_7_n_0 ),
        .I4(ir1[13]),
        .I5(ir1[11]),
        .O(\rgf_selc1_rn_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF00404000000000)) 
    \rgf_selc1_rn_wb[0]_i_9 
       (.I0(ir1[6]),
        .I1(ir1[3]),
        .I2(\stat_reg[0]_55 ),
        .I3(ir1[0]),
        .I4(ir1[8]),
        .I5(ir1[7]),
        .O(\rgf_selc1_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \rgf_selc1_rn_wb[1]_i_1 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\rgf_selc1_rn_wb[1]_i_2_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .O(\stat_reg[2]_1 [1]));
  LUT6 #(
    .INIT(64'hFF0F0F0F8F8F0F0F)) 
    \rgf_selc1_rn_wb[1]_i_10 
       (.I0(\rgf_selc1_rn_wb[1]_i_19_n_0 ),
        .I1(\stat_reg[0]_55 ),
        .I2(ir1[11]),
        .I3(ir1[1]),
        .I4(ir1[7]),
        .I5(ir1[8]),
        .O(\rgf_selc1_rn_wb[1]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \rgf_selc1_rn_wb[1]_i_11 
       (.I0(ir1[4]),
        .I1(ir1[1]),
        .I2(ir1[7]),
        .O(\rgf_selc1_rn_wb[1]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_selc1_rn_wb[1]_i_12 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .O(\rgf_selc1_rn_wb[1]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_13 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .O(\rgf_selc1_rn_wb[1]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[1]_i_14 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .O(\rgf_selc1_rn_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8000AAAA80008000)) 
    \rgf_selc1_rn_wb[1]_i_15 
       (.I0(\badr[15]_INST_0_i_90_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_20_n_0 ),
        .I2(\badrx[15]_INST_0_i_5_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_21_n_0 ),
        .I5(ir1[4]),
        .O(\rgf_selc1_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_selc1_rn_wb[1]_i_16 
       (.I0(ir1[6]),
        .I1(\stat[2]_i_10__0_n_0 ),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_22_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_19 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .O(\rgf_selc1_rn_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABBBBAAAAAAAA)) 
    \rgf_selc1_rn_wb[1]_i_2 
       (.I0(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_7_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_8_n_0 ),
        .I3(ir1[1]),
        .I4(\rgf_selc1_rn_wb[1]_i_9_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_10_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00002000F0000100)) 
    \rgf_selc1_rn_wb[1]_i_20 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .I2(ir1[6]),
        .I3(ir1[1]),
        .I4(ir1[7]),
        .I5(ir1[5]),
        .O(\rgf_selc1_rn_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0FF7FFC00FFCF)) 
    \rgf_selc1_rn_wb[1]_i_21 
       (.I0(ir1[6]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[7]),
        .O(\rgf_selc1_rn_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF2200F2002200)) 
    \rgf_selc1_rn_wb[1]_i_3 
       (.I0(\rgf_selc1_rn_wb[1]_i_11_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_12_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I4(ir1[4]),
        .I5(rst_n_fl_reg_9),
        .O(\rgf_selc1_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h7707777777777777)) 
    \rgf_selc1_rn_wb[1]_i_4 
       (.I0(\rgf_selc1_rn_wb[1]_i_11_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_14_n_0 ),
        .I3(\stat[2]_i_11_n_0 ),
        .I4(\bdatw[14]_INST_0_i_29_n_0 ),
        .I5(\rgf_selc1_rn_wb_reg[2] ),
        .O(\rgf_selc1_rn_wb[1]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[1]_i_5 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\rgf_selc1_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAEAAAFFFFEAAA)) 
    \rgf_selc1_rn_wb[1]_i_6 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_2_0 ),
        .I3(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_2_1 ),
        .I5(\rgf_selc1_rn_wb[2]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFDDDFDFDFFFFFFFF)) 
    \rgf_selc1_rn_wb[1]_i_7 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[11]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(\rgf_selc1_wb[0]_i_6_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \rgf_selc1_rn_wb[1]_i_8 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\rgf_selc1_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5555555545555555)) 
    \rgf_selc1_rn_wb[1]_i_9 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(ir1[14]),
        .I5(ir1[15]),
        .O(\rgf_selc1_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5554555554545454)) 
    \rgf_selc1_rn_wb[2]_i_1 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_3_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_5_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .O(\stat_reg[2]_1 [2]));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_selc1_rn_wb[2]_i_10 
       (.I0(ir1[6]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .O(\rgf_selc1_rn_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF000000FB)) 
    \rgf_selc1_rn_wb[2]_i_11 
       (.I0(ir1[8]),
        .I1(ir1[2]),
        .I2(\rgf_selc1_wb[1]_i_12_n_0 ),
        .I3(ir1[11]),
        .I4(rst_n_fl_reg_9),
        .I5(\rgf_selc1_rn_wb[1]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_12 
       (.I0(ir1[2]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .I5(ir1[3]),
        .O(\rgf_selc1_rn_wb[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    \rgf_selc1_rn_wb[2]_i_13 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[2]),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .O(\rgf_selc1_rn_wb[2]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_selc1_rn_wb[2]_i_14 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \rgf_selc1_rn_wb[2]_i_15 
       (.I0(ir1[9]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \rgf_selc1_rn_wb[2]_i_16 
       (.I0(\stat_reg[0]_48 ),
        .I1(brdy),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[8]),
        .O(\rgf_selc1_rn_wb[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_17 
       (.I0(\rgf_selc1_wb[0]_i_20_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[2]),
        .I3(ir1[9]),
        .I4(ir1[11]),
        .I5(ir1[10]),
        .O(\rgf_selc1_rn_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEE00FF6EFFFF)) 
    \rgf_selc1_rn_wb[2]_i_18 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\rgf_selc1_rn_wb[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004F44)) 
    \rgf_selc1_rn_wb[2]_i_2 
       (.I0(\rgf_selc1_rn_wb[2]_i_7_n_0 ),
        .I1(ir1[10]),
        .I2(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_selc1_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF4F4F4F)) 
    \rgf_selc1_rn_wb[2]_i_3 
       (.I0(\stat[2]_i_11_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[11]),
        .I3(\rgf_selc1_rn_wb_reg[2] ),
        .I4(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF88F888888888)) 
    \rgf_selc1_rn_wb[2]_i_4 
       (.I0(ir1[5]),
        .I1(rst_n_fl_reg_9),
        .I2(\rgf_selc1_rn_wb_reg[2] ),
        .I3(\rgf_selc1_rn_wb[2]_i_12_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5555FF7F777FFF7F)) 
    \rgf_selc1_rn_wb[2]_i_5 
       (.I0(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .I2(ir1[2]),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .I5(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \rgf_selc1_rn_wb[2]_i_6 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_rn_wb[2]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hD5D57555)) 
    \rgf_selc1_rn_wb[2]_i_7 
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[14]),
        .O(\rgf_selc1_rn_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hA222A2AA0000A2AA)) 
    \rgf_selc1_rn_wb[2]_i_8 
       (.I0(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I2(ir1[8]),
        .I3(ir1[7]),
        .I4(ir1[5]),
        .I5(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc1_stat_i_1
       (.I0(\stat_reg[2]_2 [1]),
        .I1(\stat_reg[2]_2 [0]),
        .O(\stat_reg[2]_19 ));
  LUT6 #(
    .INIT(64'h5554555544444444)) 
    \rgf_selc1_wb[0]_i_1 
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(\rgf_selc1_wb[0]_i_2_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_6_n_0 ),
        .O(\stat_reg[2]_2 [0]));
  LUT5 #(
    .INIT(32'hCC3E003F)) 
    \rgf_selc1_wb[0]_i_10 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[8]),
        .O(\rgf_selc1_wb[0]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF0E0)) 
    \rgf_selc1_wb[0]_i_11 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .O(\rgf_selc1_wb[0]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \rgf_selc1_wb[0]_i_12 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_selc1_wb[0]_i_20_n_0 ),
        .O(\rgf_selc1_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hEFEAFFFFFFFFFFFF)) 
    \rgf_selc1_wb[0]_i_13 
       (.I0(\stat[0]_i_19__0_n_0 ),
        .I1(ir1[4]),
        .I2(ir1[6]),
        .I3(ir1[10]),
        .I4(ir1[8]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \rgf_selc1_wb[0]_i_15 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[10]),
        .I3(ir1[7]),
        .I4(ir1[9]),
        .O(\rgf_selc1_wb[0]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAABAA)) 
    \rgf_selc1_wb[0]_i_16 
       (.I0(\rgf_selc1_wb[0]_i_21_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_selc1_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00006545)) 
    \rgf_selc1_wb[0]_i_17 
       (.I0(ir1[8]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[9]),
        .O(\rgf_selc1_wb[0]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_selc1_wb[0]_i_18 
       (.I0(ir1[8]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .O(\rgf_selc1_wb[0]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_selc1_wb[0]_i_19 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .O(\rgf_selc1_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAEAAAAAAAA)) 
    \rgf_selc1_wb[0]_i_2 
       (.I0(\rgf_selc1_wb[0]_i_7_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_9_n_0 ),
        .I3(ir1[4]),
        .I4(ir1[9]),
        .I5(\stat[2]_i_13__0_n_0 ),
        .O(\rgf_selc1_wb[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFBFB7BE)) 
    \rgf_selc1_wb[0]_i_20 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .I2(ir1[7]),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .O(\rgf_selc1_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0404000000000004)) 
    \rgf_selc1_wb[0]_i_21 
       (.I0(\rgf_selc1_wb[1]_i_12_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(rst_n_fl_reg_9),
        .I4(ir1[11]),
        .I5(ir1[8]),
        .O(\rgf_selc1_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2E2EEE2)) 
    \rgf_selc1_wb[0]_i_3 
       (.I0(\rgf_selc1_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_12_n_0 ),
        .I3(\stat_reg[0]_55 ),
        .I4(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I5(\rgf_selc1_wb_reg[0] ),
        .O(\rgf_selc1_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00400000)) 
    \rgf_selc1_wb[0]_i_4 
       (.I0(\stat_reg[0]_48 ),
        .I1(brdy),
        .I2(ir1[11]),
        .I3(ir1[6]),
        .I4(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_16_n_0 ),
        .O(\rgf_selc1_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55551555)) 
    \rgf_selc1_wb[0]_i_5 
       (.I0(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\rgf_selc1_wb[0]_i_18_n_0 ),
        .I3(brdy),
        .I4(\stat_reg[0]_48 ),
        .I5(\rgf_selc1_wb[0]_i_19_n_0 ),
        .O(\rgf_selc1_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc1_wb[0]_i_6 
       (.I0(ir1[13]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(ir1[15]),
        .O(\rgf_selc1_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h228200008AAA0000)) 
    \rgf_selc1_wb[0]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_53_0 ),
        .I1(ir1[12]),
        .I2(ir1[11]),
        .I3(ir1[13]),
        .I4(ir1[15]),
        .I5(ir1[14]),
        .O(\rgf_selc1_wb[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0440)) 
    \rgf_selc1_wb[0]_i_8 
       (.I0(ir1[0]),
        .I1(ir1[2]),
        .I2(ir1[1]),
        .I3(ir1[3]),
        .O(\rgf_selc1_wb[0]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_wb[0]_i_9 
       (.I0(ir1[11]),
        .I1(ir1[10]),
        .O(\rgf_selc1_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFEEAE)) 
    \rgf_selc1_wb[1]_i_1 
       (.I0(\stat_reg[1]_6 ),
        .I1(\rgf_selc1_wb_reg[1]_0 ),
        .I2(\rgf_selc1_wb[1]_i_3_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_4_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_5_n_0 ),
        .I5(\rgf_selc1_wb_reg[1] [2]),
        .O(\stat_reg[2]_2 [1]));
  LUT5 #(
    .INIT(32'h0000FFDF)) 
    \rgf_selc1_wb[1]_i_10 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .I3(ir1[8]),
        .I4(rst_n_fl_reg_9),
        .O(\rgf_selc1_wb[1]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \rgf_selc1_wb[1]_i_11 
       (.I0(\stat_reg[0]_48 ),
        .I1(brdy),
        .I2(ir1[11]),
        .I3(ir1[6]),
        .O(\rgf_selc1_wb[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_selc1_wb[1]_i_12 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .I2(ir1[10]),
        .O(\rgf_selc1_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFFBFFF3FFFBFF)) 
    \rgf_selc1_wb[1]_i_13 
       (.I0(\sr_reg[15]_0 [6]),
        .I1(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I2(ir1[15]),
        .I3(ir1[13]),
        .I4(ir1[12]),
        .I5(ir1[14]),
        .O(\rgf_selc1_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEEEFEFE)) 
    \rgf_selc1_wb[1]_i_14 
       (.I0(\rgf_selc1_wb[1]_i_20_n_0 ),
        .I1(\rgf_selc1_wb_reg[1]_i_21_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_22_n_0 ),
        .I3(\stat_reg[0]_48 ),
        .I4(brdy),
        .I5(\rgf_selc1_wb[1]_i_23_n_0 ),
        .O(\rgf_selc1_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000303C0808)) 
    \rgf_selc1_wb[1]_i_15 
       (.I0(\stat_reg[0]_55 ),
        .I1(ir1[1]),
        .I2(ir1[3]),
        .I3(ir1[0]),
        .I4(ir1[2]),
        .I5(\rgf_selc1_wb[1]_i_24_n_0 ),
        .O(\rgf_selc1_wb[1]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h11110010)) 
    \rgf_selc1_wb[1]_i_16 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[13]),
        .I2(\rgf_selc1_wb[1]_i_5_0 ),
        .I3(\rgf_selc1_wb[1]_i_26_n_0 ),
        .I4(ir1[15]),
        .O(\rgf_selc1_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCC5D00C0CC5D0000)) 
    \rgf_selc1_wb[1]_i_17 
       (.I0(\rgf_selc1_wb[1]_i_5_1 ),
        .I1(\rgf_selc1_wb[1]_i_5_2 ),
        .I2(ir1[11]),
        .I3(ir1[14]),
        .I4(ir1[15]),
        .I5(\sr_reg[15]_0 [6]),
        .O(\rgf_selc1_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_selc1_wb[1]_i_18 
       (.I0(\bcmd[0]_INST_0_i_7_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I4(ir1[12]),
        .I5(ir1[14]),
        .O(\rgf_selc1_wb[1]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h10000111)) 
    \rgf_selc1_wb[1]_i_19 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[14]),
        .I2(\sr_reg[15]_0 [7]),
        .I3(ir1[12]),
        .I4(ir1[11]),
        .O(\rgf_selc1_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \rgf_selc1_wb[1]_i_2 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\rgf_selc1_wb[1]_i_6_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .O(\stat_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h55775577557755F7)) 
    \rgf_selc1_wb[1]_i_20 
       (.I0(ir1[8]),
        .I1(ir1[10]),
        .I2(ir1[11]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[1]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h80888888)) 
    \rgf_selc1_wb[1]_i_22 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[9]),
        .I2(ir1[5]),
        .I3(ir1[11]),
        .I4(ir1[10]),
        .O(\rgf_selc1_wb[1]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf_selc1_wb[1]_i_23 
       (.I0(\rgf_selc1_wb[1]_i_31_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_32_n_0 ),
        .I3(rst_n_fl_reg_9),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .O(\rgf_selc1_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    \rgf_selc1_wb[1]_i_24 
       (.I0(\stat[0]_i_11__0_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[13]),
        .I3(\bdatw[11]_INST_0_i_28_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_34_n_0 ),
        .O(\rgf_selc1_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0606060605000505)) 
    \rgf_selc1_wb[1]_i_26 
       (.I0(ir1[11]),
        .I1(\sr_reg[15]_0 [5]),
        .I2(ir1[12]),
        .I3(\badr[15]_INST_0_i_175_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I5(ir1[14]),
        .O(\rgf_selc1_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h77FF77FFFF0FFFFF)) 
    \rgf_selc1_wb[1]_i_29 
       (.I0(\rgf_selc1_wb[1]_i_35_n_0 ),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[11]),
        .I4(ir1[6]),
        .I5(ir1[9]),
        .O(\rgf_selc1_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFABFFABFFABAAAA)) 
    \rgf_selc1_wb[1]_i_3 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb[1]_i_7_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_8_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_9_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_10_n_0 ),
        .I5(\badrx[15]_INST_0_i_6_n_0 ),
        .O(\rgf_selc1_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEE00EE00F0FFFFFF)) 
    \rgf_selc1_wb[1]_i_30 
       (.I0(\stat[0]_i_19__0_n_0 ),
        .I1(\stat[0]_i_21__0_n_0 ),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(\rgf_selc1_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h000000041010001C)) 
    \rgf_selc1_wb[1]_i_31 
       (.I0(ir1[8]),
        .I1(ir1[11]),
        .I2(ir1[10]),
        .I3(ir1[7]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[9]),
        .O(\rgf_selc1_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000007F00000000)) 
    \rgf_selc1_wb[1]_i_32 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(ir1[10]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[11]),
        .O(\rgf_selc1_wb[1]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc1_wb[1]_i_33 
       (.I0(ir1[7]),
        .I1(ir1[5]),
        .I2(ir1[6]),
        .I3(ir1[4]),
        .O(\rgf_selc1_wb[1]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc1_wb[1]_i_34 
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .O(\rgf_selc1_wb[1]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h1E001F81)) 
    \rgf_selc1_wb[1]_i_35 
       (.I0(ir1[4]),
        .I1(ir1[6]),
        .I2(ir1[5]),
        .I3(ir1[7]),
        .I4(ir1[3]),
        .O(\rgf_selc1_wb[1]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000EA0000)) 
    \rgf_selc1_wb[1]_i_4 
       (.I0(\rgf_selc1_wb[1]_i_11_n_0 ),
        .I1(ir1[11]),
        .I2(ir1[8]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_12_n_0 ),
        .O(\rgf_selc1_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FFF1)) 
    \rgf_selc1_wb[1]_i_5 
       (.I0(\rgf_selc1_wb[1]_i_13_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_14_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_16_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(\rgf_selc1_wb[1]_i_17_n_0 ),
        .O(\rgf_selc1_wb[1]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_wb[1]_i_6 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .O(\rgf_selc1_wb[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h0020AAAA)) 
    \rgf_selc1_wb[1]_i_7 
       (.I0(ir1[0]),
        .I1(\stat_reg[0]_48 ),
        .I2(brdy),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[1]),
        .O(\rgf_selc1_wb[1]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    \rgf_selc1_wb[1]_i_8 
       (.I0(ir1[1]),
        .I1(ir1[3]),
        .I2(ir1[2]),
        .O(\rgf_selc1_wb[1]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFDFDFDDD)) 
    \rgf_selc1_wb[1]_i_9 
       (.I0(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I1(ir1[13]),
        .I2(ir1[0]),
        .I3(ir1[3]),
        .I4(ir1[2]),
        .O(\rgf_selc1_wb[1]_i_9_n_0 ));
  MUXF7 \rgf_selc1_wb_reg[1]_i_21 
       (.I0(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_30_n_0 ),
        .O(\rgf_selc1_wb_reg[1]_i_21_n_0 ),
        .S(\rgf_selc1_wb_reg[1] [0]));
  FDRE rst_n_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(rst_n_fl),
        .R(\<const0> ));
  LUT4 #(
    .INIT(16'hFD08)) 
    \sp[0]_i_2 
       (.I0(\stat_reg[0]_0 ),
        .I1(\sp_reg[0] ),
        .I2(\stat_reg[0]_1 ),
        .I3(\sp_reg[0]_0 ),
        .O(\sp[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFAFEFFBEFAFFFFBF)) 
    \sp[15]_i_10 
       (.I0(\sp[15]_i_21_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[3]),
        .I3(ir1[5]),
        .I4(ir1[6]),
        .I5(ir1[0]),
        .O(\sp[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF3EFF3EFF3EFFFF)) 
    \sp[15]_i_11 
       (.I0(ir1[2]),
        .I1(ir1[8]),
        .I2(ir1[9]),
        .I3(\sp[15]_i_22_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(ctl_fetch1_fl_i_20_n_0),
        .O(\sp[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF2FFFFFFFFFF2)) 
    \sp[15]_i_13 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .I2(ir0[8]),
        .I3(ir0[9]),
        .I4(\badr[15]_INST_0_i_195_n_0 ),
        .I5(ir0[7]),
        .O(\sp[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8FFF8FF88FFF8FFF)) 
    \sp[15]_i_14 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(\bcmd[0]_INST_0_i_23_n_0 ),
        .I2(ir0[6]),
        .I3(ir0[5]),
        .I4(ir0[3]),
        .I5(ir0[1]),
        .O(\sp[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0089008900890000)) 
    \sp[15]_i_15 
       (.I0(ir0[6]),
        .I1(ir0[7]),
        .I2(ir0[4]),
        .I3(\sp[15]_i_8_0 ),
        .I4(\bcmd[0]_INST_0_i_9_n_0 ),
        .I5(\ccmd[4]_INST_0_i_15_n_0 ),
        .O(\sp[15]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFEFFE)) 
    \sp[15]_i_16 
       (.I0(\sp[15]_i_23_n_0 ),
        .I1(\bcmd[0]_INST_0_i_16_n_0 ),
        .I2(ir1[7]),
        .I3(ir1[6]),
        .I4(ir1[4]),
        .I5(\sp[15]_i_24_n_0 ),
        .O(\sp[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    \sp[15]_i_17 
       (.I0(fch_irq_req),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[12]),
        .I3(ir0[11]),
        .I4(ir0[9]),
        .I5(ir0[6]),
        .O(\sp[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFEBFFFAEFEBFFFBF)) 
    \sp[15]_i_18 
       (.I0(\bcmd[1]_INST_0_i_9_n_0 ),
        .I1(ir0[5]),
        .I2(ir0[6]),
        .I3(ir0[3]),
        .I4(ir0[7]),
        .I5(ir0[0]),
        .O(\sp[15]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sp[15]_i_19 
       (.I0(ir0[11]),
        .I1(ir0[12]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\sp[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hBFBFBFBEFFFFBFBE)) 
    \sp[15]_i_20 
       (.I0(\sp[15]_i_8_0 ),
        .I1(ir0[7]),
        .I2(ir0[8]),
        .I3(ir0[1]),
        .I4(ir0[4]),
        .I5(ir0[6]),
        .O(\sp[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFBFFFFF00)) 
    \sp[15]_i_21 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[12]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(ir1[6]),
        .O(\sp[15]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3F3EFF3E)) 
    \sp[15]_i_22 
       (.I0(ir1[1]),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[4]),
        .I4(ir1[6]),
        .O(\sp[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFF7EFFFFFFFF7E7E)) 
    \sp[15]_i_23 
       (.I0(ir1[9]),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[12]),
        .I5(ir1[11]),
        .O(\sp[15]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFFFFFFEAFFFFFFF)) 
    \sp[15]_i_24 
       (.I0(\bcmd[1]_INST_0_i_17_n_0 ),
        .I1(ir1[2]),
        .I2(ir1[6]),
        .I3(ir1[5]),
        .I4(ir1[3]),
        .I5(ir1[1]),
        .O(\sp[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAFEAAAAAAAA)) 
    \sp[15]_i_5 
       (.I0(ctl_sp_dec0),
        .I1(\sp[15]_i_9_n_0 ),
        .I2(ir1[10]),
        .I3(\sp[15]_i_10_n_0 ),
        .I4(\sp[15]_i_11_n_0 ),
        .I5(\sp[15]_i_2 ),
        .O(\stat_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0100FFFF01000100)) 
    \sp[15]_i_6 
       (.I0(\sp[15]_i_13_n_0 ),
        .I1(\sp[15]_i_14_n_0 ),
        .I2(\bcmd[1]_INST_0_i_8_n_0 ),
        .I3(\sp[15]_i_15_n_0 ),
        .I4(\sp[15]_i_16_n_0 ),
        .I5(\sp[15]_i_2 ),
        .O(\stat_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0000000030220022)) 
    \sp[15]_i_8 
       (.I0(\sp[15]_i_17_n_0 ),
        .I1(\sp[15]_i_18_n_0 ),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(\sp[15]_i_19_n_0 ),
        .I5(\sp[15]_i_20_n_0 ),
        .O(ctl_sp_dec0));
  LUT4 #(
    .INIT(16'h1110)) 
    \sp[15]_i_9 
       (.I0(ir1[12]),
        .I1(ir1[11]),
        .I2(fch_irq_req),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .O(\sp[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF51BB0000)) 
    \sr[13]_i_11 
       (.I0(ir0[13]),
        .I1(ir0[14]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .I4(ir0[15]),
        .I5(\sr[13]_i_12_n_0 ),
        .O(\sr[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000003A0AFA0A)) 
    \sr[13]_i_12 
       (.I0(\sr[13]_i_13_n_0 ),
        .I1(\stat[0]_i_18_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_12_n_0 ),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(\sr[13]_i_14_n_0 ),
        .O(\sr[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AA040004)) 
    \sr[13]_i_13 
       (.I0(ir0[9]),
        .I1(ir0[6]),
        .I2(fctl_n_91),
        .I3(ir0[11]),
        .I4(ir0[10]),
        .I5(\sr[13]_i_15_n_0 ),
        .O(\sr[13]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \sr[13]_i_14 
       (.I0(ir0[15]),
        .I1(ir0[12]),
        .I2(ir0[13]),
        .O(\sr[13]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFBFF0FFC0FFC0FFC)) 
    \sr[13]_i_15 
       (.I0(ir0[3]),
        .I1(ir0[4]),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(ir0[9]),
        .I5(ir0[5]),
        .O(\sr[13]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00000200)) 
    \sr[13]_i_3 
       (.I0(\sr[13]_i_6_n_0 ),
        .I1(\sr[13]_i_7_n_0 ),
        .I2(ir0[3]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\sr[13]_i_8_n_0 ),
        .O(ctl_sr_ldie0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[13]_i_6 
       (.I0(\bcmd[1]_INST_0_i_13_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[10]),
        .I3(ir0[7]),
        .I4(ir0[9]),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\sr[13]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[13]_i_7 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(ir0[1]),
        .I2(ir0[2]),
        .O(\sr[13]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \sr[13]_i_8 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(ir0[11]),
        .I2(brdy),
        .I3(ir0[0]),
        .O(\sr[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    \sr[13]_i_9 
       (.I0(\sr[13]_i_11_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(\rgf_selc0_rn_wb_reg[0] [2]),
        .I4(ir0[14]),
        .I5(ir0[15]),
        .O(ctl_sr_upd0));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \sr[15]_i_5 
       (.I0(\sr[15]_i_2 ),
        .I1(ir1[11]),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(ir1[1]),
        .I4(\sr[15]_i_9_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .O(ctl_sr_ldie1));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \sr[15]_i_9 
       (.I0(ir1[2]),
        .I1(ir1[3]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .O(\sr[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFFEAFFFFFFEA)) 
    \sr[3]_i_7 
       (.I0(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(cbus_i[2]),
        .I3(\sr[3]_i_3 ),
        .I4(\rgf_c0bus_wb_reg[3] [3]),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\sr[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEFEFFFFEEFE)) 
    \sr[4]_i_10 
       (.I0(\sr[4]_i_29_n_0 ),
        .I1(\sr[4]_i_30_n_0 ),
        .I2(\sr[4]_i_31_n_0 ),
        .I3(\sr[4]_i_32_n_0 ),
        .I4(\sr[4]_i_33_n_0 ),
        .I5(\sr[4]_i_34_n_0 ),
        .O(\sr[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBABFBABAAAAAAAAA)) 
    \sr[4]_i_100 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\sr[4]_i_35_0 ),
        .I2(\rgf_c1bus_wb[15]_i_14_0 ),
        .I3(\sr[4]_i_170_n_0 ),
        .I4(\sr[4]_i_171_n_0 ),
        .I5(\tr_reg[4]_0 ),
        .O(\sr[4]_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h0A22FFFF0A220A22)) 
    \sr[4]_i_101 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_25_0 ),
        .I2(\sr[4]_i_36_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\stat_reg[2]_4 ),
        .I5(\rgf_c1bus_wb[15]_i_14_1 ),
        .O(\sr[4]_i_101_n_0 ));
  LUT6 #(
    .INIT(64'h00FD00FD000000FD)) 
    \sr[4]_i_102 
       (.I0(\rgf_c1bus_wb[15]_i_14_0 ),
        .I1(\sr[4]_i_172_n_0 ),
        .I2(\sr[4]_i_36_1 ),
        .I3(\sr[4]_i_174_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\sr[4]_i_36_2 ),
        .O(\sr[4]_i_102_n_0 ));
  LUT5 #(
    .INIT(32'h00088808)) 
    \sr[4]_i_103 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(\sr[4]_i_37_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb_reg[4]_1 ),
        .O(\sr[4]_i_103_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBBA)) 
    \sr[4]_i_104 
       (.I0(\stat_reg[2]_4 ),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(\sr[6]_i_6_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\sr[4]_i_104_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_106 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .O(\sr[4]_i_106_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[4]_i_107 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\rgf_c1bus_wb_reg[13]_6 ),
        .O(\sr[4]_i_107_n_0 ));
  LUT6 #(
    .INIT(64'h000F0B0B000F0000)) 
    \sr[4]_i_108 
       (.I0(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I1(\stat_reg[2]_8 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[13]_i_2_0 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .O(\sr[4]_i_108_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF2700)) 
    \sr[4]_i_109 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[11]_i_6_0 ),
        .I2(\rgf_c1bus_wb[15]_i_4_0 ),
        .I3(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_14_1 ),
        .I5(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .O(\sr[4]_i_109_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEEFFFFEFEE)) 
    \sr[4]_i_11 
       (.I0(\sr[4]_i_35_n_0 ),
        .I1(\sr[4]_i_36_n_0 ),
        .I2(\sr[4]_i_37_n_0 ),
        .I3(\sr[4]_i_38_n_0 ),
        .I4(\sr[4]_i_39_n_0 ),
        .I5(\sr[4]_i_40_n_0 ),
        .O(\sr[4]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \sr[4]_i_110 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_35_1 ),
        .O(\sr[4]_i_110_n_0 ));
  LUT6 #(
    .INIT(64'hFF005D0000005D00)) 
    \sr[4]_i_111 
       (.I0(\stat_reg[2]_8 ),
        .I1(\sr[4]_i_177_n_0 ),
        .I2(\sr[4]_i_178_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .I5(\sr[4]_i_41_0 ),
        .O(\sr[4]_i_111_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAABABF)) 
    \sr[4]_i_112 
       (.I0(\rgf_c1bus_wb[15]_i_14_1 ),
        .I1(\sr[4]_i_46_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_29_3 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\bdatw[9]_INST_0_i_16_0 ),
        .O(\sr[4]_i_112_n_0 ));
  LUT5 #(
    .INIT(32'h8A80FFFF)) 
    \sr[4]_i_113 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_43_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_43_1 ),
        .I4(\tr_reg[4]_0 ),
        .O(\sr[4]_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBEEFBBBFBAAFB)) 
    \sr[4]_i_114 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\sr[4]_i_43_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(\sr[4]_i_45_0 ),
        .I5(\sr[4]_i_34_0 ),
        .O(\sr[4]_i_114_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \sr[4]_i_116 
       (.I0(\stat_reg[2]_7 ),
        .I1(\rgf_c1bus_wb[15]_i_4_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_33_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .O(\sr[4]_i_116_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \sr[4]_i_117 
       (.I0(\stat_reg[2]_8 ),
        .I1(\rgf_c1bus_wb_reg[2]_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .O(\sr[4]_i_117_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAFBABFFFFFBAB)) 
    \sr[4]_i_118 
       (.I0(\stat_reg[2]_8 ),
        .I1(\sr[4]_i_43_2 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_43_1 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .I5(\sr[4]_i_46_1 ),
        .O(\sr[4]_i_118_n_0 ));
  LUT6 #(
    .INIT(64'h00002320FFFFFFFF)) 
    \sr[4]_i_119 
       (.I0(\sr[4]_i_46_1 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_46_2 ),
        .I4(\stat_reg[2]_4 ),
        .I5(\tr_reg[4]_0 ),
        .O(\sr[4]_i_119_n_0 ));
  LUT6 #(
    .INIT(64'h0000000054540054)) 
    \sr[4]_i_12 
       (.I0(\sr[4]_i_41_n_0 ),
        .I1(\sr[4]_i_42_n_0 ),
        .I2(\sr[4]_i_43_n_0 ),
        .I3(\sr[4]_i_44_n_0 ),
        .I4(\sr[4]_i_45_n_0 ),
        .I5(\sr[4]_i_46_n_0 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA00000000303F)) 
    \sr[4]_i_120 
       (.I0(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .I1(\sr[4]_i_29_3 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[9]_i_3_1 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\bdatw[9]_INST_0_i_16_0 ),
        .O(\sr[4]_i_120_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FDFFFDDD)) 
    \sr[4]_i_121 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\sr[4]_i_44_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\sr[4]_i_46_0 ),
        .I5(\rgf_c1bus_wb[15]_i_14_1 ),
        .O(\sr[4]_i_121_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFCFCFCFCFFF)) 
    \sr[4]_i_124 
       (.I0(tout__1_carry_i_14_n_0),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .O(\sr[4]_i_124_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \sr[4]_i_125 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(a0bus_0[6]),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\sr[4]_i_125_n_0 ));
  LUT6 #(
    .INIT(64'hE0E020E0FFFFFFFF)) 
    \sr[4]_i_126 
       (.I0(\sr[4]_i_54_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\tr_reg[4] ),
        .I3(\rgf_c0bus_wb[11]_i_3_0 ),
        .I4(\sr[4]_i_54_1 ),
        .I5(\rgf_c0bus_wb[15]_i_7_0 ),
        .O(\sr[4]_i_126_n_0 ));
  LUT6 #(
    .INIT(64'h1111303311113000)) 
    \sr[4]_i_127 
       (.I0(\sr[4]_i_185_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I2(\sr[4]_i_55_1 ),
        .I3(\bbus_o[2]_INST_0_i_1_0 ),
        .I4(\stat_reg[1]_1 ),
        .I5(\sr[4]_i_55_2 ),
        .O(\sr[4]_i_127_n_0 ));
  LUT6 #(
    .INIT(64'h8088AAAA80888888)) 
    \sr[4]_i_129 
       (.I0(\stat_reg[2]_10 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb_reg[11]_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr[4]_i_55_0 ),
        .O(\sr[4]_i_129_n_0 ));
  LUT6 #(
    .INIT(64'h2233332000000020)) 
    \sr[4]_i_13 
       (.I0(\sr_reg[15]_0 [4]),
        .I1(\sr[4]_i_3_0 ),
        .I2(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[2]_4 ),
        .I5(tout__1_carry_i_11_n_0),
        .O(\sr[4]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \sr[4]_i_132 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(a0bus_0[12]),
        .I2(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\rgf_c0bus_wb[13]_i_10_0 ));
  LUT6 #(
    .INIT(64'hA2A2A2808080A280)) 
    \sr[4]_i_134 
       (.I0(\stat_reg[2]_10 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\sr[4]_i_60_1 ),
        .I3(\sr[4]_i_65_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .I5(\sr[4]_i_60_0 ),
        .O(\sr[4]_i_134_n_0 ));
  LUT5 #(
    .INIT(32'hFFFBAAAA)) 
    \sr[4]_i_136 
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_3_1 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[4]_i_9_n_0 ),
        .O(\sr[4]_i_136_n_0 ));
  LUT5 #(
    .INIT(32'hAA22A2A2)) 
    \sr[4]_i_137 
       (.I0(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb_reg[8]_1 ),
        .I3(\rgf_c0bus_wb_reg[8]_2 ),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\sr[4]_i_137_n_0 ));
  LUT6 #(
    .INIT(64'hE4E4EE44FFFFFFFF)) 
    \sr[4]_i_139 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\sr[4]_i_63_0 ),
        .I2(\sr[4]_i_63_1 ),
        .I3(\rgf_c0bus_wb_reg[2]_0 ),
        .I4(\rgf_c0bus_wb[11]_i_3_0 ),
        .I5(\tr_reg[4] ),
        .O(\sr[4]_i_139_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \sr[4]_i_14 
       (.I0(\sr[4]_i_48_n_0 ),
        .I1(\sr[4]_i_49_n_0 ),
        .I2(\sr[4]_i_50_n_0 ),
        .I3(\sr[4]_i_51_n_0 ),
        .I4(\sr[4]_i_52_n_0 ),
        .I5(\sr[4]_i_53_n_0 ),
        .O(\sr[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \sr[4]_i_140 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_2 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_64_0 ),
        .I4(\bbus_o[2]_INST_0_i_1_0 ),
        .O(\sr[4]_i_140_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_141 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(a0bus_0[5]),
        .O(\sr[4]_i_141_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \sr[4]_i_143 
       (.I0(\sr[4]_i_201_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[1]_i_3_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\rgf_c0bus_wb[9]_i_3_0 ),
        .I5(\stat_reg[2]_10 ),
        .O(\sr[4]_i_143_n_0 ));
  LUT6 #(
    .INIT(64'h4F405F5F4F405050)) 
    \sr[4]_i_144 
       (.I0(\rgf_c0bus_wb[11]_i_3_0 ),
        .I1(\badr[1]_INST_0_i_2 ),
        .I2(\bbus_o[2]_INST_0_i_1_0 ),
        .I3(\sr[4]_i_66_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_0 ),
        .I5(\rgf_c0bus_wb[5]_i_2_0 ),
        .O(\sr[4]_i_144_n_0 ));
  LUT4 #(
    .INIT(16'hBAFE)) 
    \sr[4]_i_145 
       (.I0(\rgf_c0bus_wb[11]_i_11_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb[14]_i_5_0 ),
        .I3(\rgf_c0bus_wb[5]_i_2_1 ),
        .O(\sr[4]_i_145_n_0 ));
  LUT6 #(
    .INIT(64'hB080FFFFB080B080)) 
    \sr[4]_i_147 
       (.I0(\rgf_c0bus_wb[5]_i_3_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\stat_reg[2]_10 ),
        .I3(\sr[4]_i_67_0 ),
        .I4(\rgf_c0bus_wb[5]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\sr[4]_i_147_n_0 ));
  LUT5 #(
    .INIT(32'h14405400)) 
    \sr[4]_i_149 
       (.I0(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb_reg[5] ),
        .I2(a0bus_0[5]),
        .I3(\stat_reg[1]_1 ),
        .I4(\stat_reg[2]_10 ),
        .O(\sr[4]_i_149_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEFFFE)) 
    \sr[4]_i_15 
       (.I0(\sr[4]_i_54_n_0 ),
        .I1(\sr[4]_i_55_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I3(\tr_reg[4] ),
        .I4(\sr[4]_i_56_n_0 ),
        .I5(\sr[4]_i_6_0 ),
        .O(\sr[4]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF75770000)) 
    \sr[4]_i_150 
       (.I0(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .I2(\sr[4]_i_204_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .O(\sr[4]_i_150_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFFFEFCFFFCFCF)) 
    \sr[4]_i_151 
       (.I0(\ccmd[0]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[0]_3 ),
        .I2(\ccmd[4]_INST_0_i_2_n_0 ),
        .I3(\ccmd[2]_INST_0_i_1_n_0 ),
        .I4(\ccmd[1]_INST_0_i_1_n_0 ),
        .I5(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_151_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \sr[4]_i_153 
       (.I0(\stat_reg[1]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\sr[4]_i_153_n_0 ));
  LUT5 #(
    .INIT(32'hCCCC440C)) 
    \sr[4]_i_157 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(a1bus_0[8]),
        .I3(\stat_reg[1]_0 ),
        .I4(\stat_reg[2]_4 ),
        .O(\sr[4]_i_157_n_0 ));
  LUT5 #(
    .INIT(32'h33BF33B3)) 
    \sr[4]_i_158 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(\stat_reg[1]_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(a1bus_0[14]),
        .O(\sr[4]_i_158_n_0 ));
  LUT6 #(
    .INIT(64'h54FF000054540000)) 
    \sr[4]_i_16 
       (.I0(\sr[4]_i_58_n_0 ),
        .I1(\sr[4]_i_59_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_7_0 ),
        .I5(\sr[4]_i_60_n_0 ),
        .O(\sr[4]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFF47FFFF)) 
    \sr[4]_i_163 
       (.I0(a1bus_0[1]),
        .I1(\tr_reg[0] ),
        .I2(a1bus_0[0]),
        .I3(\bdatw[8]_INST_0_i_16_1 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .O(\sr[4]_i_163_n_0 ));
  LUT6 #(
    .INIT(64'hBBBFFFBFAAAEEEAE)) 
    \sr[4]_i_167 
       (.I0(\sr[4]_i_221_n_0 ),
        .I1(\bdatw[8]_INST_0_i_16_1 ),
        .I2(a1bus_0[13]),
        .I3(\tr_reg[0] ),
        .I4(a1bus_0[14]),
        .I5(\sr[4]_i_91 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'h1511155504000444)) 
    \sr[4]_i_168 
       (.I0(\sr[4]_i_222_n_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\sr[4]_i_98_0 ),
        .I3(\bdatw[8]_INST_0_i_16_1 ),
        .I4(\sr[4]_i_98_1 ),
        .I5(a1bus_0[15]),
        .O(\sr[4]_i_168_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFEFEFFFFFFFEF)) 
    \sr[4]_i_17 
       (.I0(\sr[4]_i_61_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr[4]_i_62_n_0 ),
        .O(\sr[4]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h08000888)) 
    \sr[4]_i_170 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\bdatw[8]_INST_0_i_16_0 ),
        .I2(\sr[4]_i_100_1 ),
        .I3(\bdatw[8]_INST_0_i_16_1 ),
        .I4(\sr[4]_i_100_2 ),
        .O(\sr[4]_i_170_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAFEE)) 
    \sr[4]_i_171 
       (.I0(\stat_reg[2]_4 ),
        .I1(\sr[4]_i_91 ),
        .I2(\sr[4]_i_100_0 ),
        .I3(\bdatw[8]_INST_0_i_16_1 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\bdatw[8]_INST_0_i_16_0 ),
        .O(\sr[4]_i_171_n_0 ));
  LUT6 #(
    .INIT(64'h080808A8A8A808A8)) 
    \sr[4]_i_172 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_102_0 ),
        .I2(\bdatw[8]_INST_0_i_16_1 ),
        .I3(a1bus_0[14]),
        .I4(\tr_reg[0] ),
        .I5(a1bus_0[15]),
        .O(\sr[4]_i_172_n_0 ));
  LUT5 #(
    .INIT(32'h0004FFFF)) 
    \sr[4]_i_174 
       (.I0(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\stat_reg[2]_8 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\tr_reg[4]_0 ),
        .O(\sr[4]_i_174_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \sr[4]_i_176 
       (.I0(\stat_reg[1]_0 ),
        .I1(a1bus_0[15]),
        .I2(\stat_reg[2]_4 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .O(\stat_reg[2]_9 ));
  LUT6 #(
    .INIT(64'hABFBAAAAABFBFFFF)) 
    \sr[4]_i_177 
       (.I0(\bdatw[8]_INST_0_i_16_0 ),
        .I1(a1bus_0[9]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[10]),
        .I4(\bdatw[8]_INST_0_i_16_1 ),
        .I5(\sr[4]_i_111_0 ),
        .O(\sr[4]_i_177_n_0 ));
  LUT6 #(
    .INIT(64'hA808FD5D00000000)) 
    \sr[4]_i_178 
       (.I0(\bdatw[8]_INST_0_i_16_1 ),
        .I1(a1bus_0[13]),
        .I2(\tr_reg[0] ),
        .I3(a1bus_0[14]),
        .I4(\sr[4]_i_91 ),
        .I5(\bdatw[8]_INST_0_i_16_0 ),
        .O(\sr[4]_i_178_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002022)) 
    \sr[4]_i_18 
       (.I0(\sr[4]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I2(\sr[4]_i_64_n_0 ),
        .I3(\sr[4]_i_65_n_0 ),
        .I4(\sr[4]_i_66_n_0 ),
        .I5(\sr[4]_i_67_n_0 ),
        .O(\sr[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8D888DDDCCCCCCCC)) 
    \sr[4]_i_185 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(a0bus_0[15]),
        .I2(\sr[4]_i_127_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_0 ),
        .I4(\sr[4]_i_127_1 ),
        .I5(\bbus_o[1]_INST_0_i_1_0 ),
        .O(\sr[4]_i_185_n_0 ));
  LUT5 #(
    .INIT(32'h000000C5)) 
    \sr[4]_i_188 
       (.I0(\sr[4]_i_128 ),
        .I1(\sr[4]_i_128_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_0 ),
        .I4(\stat_reg[1]_1 ),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hF5FF000055440000)) 
    \sr[4]_i_19 
       (.I0(\rgf_c0bus_wb[12]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_7_n_0 ),
        .I3(\tr_reg[4] ),
        .I4(\rgf_c0bus_wb[15]_i_7_0 ),
        .I5(\sr[4]_i_68_n_0 ),
        .O(\sr[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h010001000100FFFF)) 
    \sr[4]_i_20 
       (.I0(\sr[4]_i_69_n_0 ),
        .I1(\sr[4]_i_70_n_0 ),
        .I2(\sr[4]_i_71_n_0 ),
        .I3(\sr[4]_i_72_n_0 ),
        .I4(\sr[4]_i_73_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\sr[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00007F007F007F00)) 
    \sr[4]_i_201 
       (.I0(\ccmd[0]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[15]),
        .I2(\stat_reg[1]_1 ),
        .I3(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I4(a0bus_0[8]),
        .I5(\rgf_c0bus_wb[11]_i_3_0 ),
        .O(\sr[4]_i_201_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \sr[4]_i_204 
       (.I0(a0bus_0[12]),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .I2(\stat_reg[1]_1 ),
        .O(\sr[4]_i_204_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \sr[4]_i_21 
       (.I0(ir1[9]),
        .I1(ir1[10]),
        .I2(ir1[8]),
        .O(\sr[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1100000111004001)) 
    \sr[4]_i_22 
       (.I0(\sr[4]_i_74_n_0 ),
        .I1(\sr[4]_i_75_n_0 ),
        .I2(ir1[4]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(ir1[3]),
        .O(\sr[4]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hAAFBFFAE)) 
    \sr[4]_i_221 
       (.I0(\stat_reg[1]_0 ),
        .I1(\tr_reg[0] ),
        .I2(\bdatw[9]_INST_0_i_16_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\bdatw[10]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_221_n_0 ));
  LUT6 #(
    .INIT(64'hFF0400FBFFFFFFFF)) 
    \sr[4]_i_222 
       (.I0(\bdatw[9]_INST_0_i_16_n_0 ),
        .I1(\tr_reg[0] ),
        .I2(\bdatw[10]_INST_0_i_16_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\sr[4]_i_222_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAFFEAAFFFF)) 
    \sr[4]_i_23 
       (.I0(\sr[4]_i_76_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[9]),
        .I3(ir1[10]),
        .I4(ir1[11]),
        .I5(ir1[8]),
        .O(\sr[4]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0A02A2A2)) 
    \sr[4]_i_24 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[11]),
        .I4(ir1[12]),
        .O(\sr[4]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFFFEAAAAAAAA)) 
    \sr[4]_i_25 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I2(\sr[4]_i_77_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb_reg[12]_0 ),
        .I5(\rgf_c1bus_wb[12]_i_10_n_0 ),
        .O(\sr[4]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \sr[4]_i_258 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [11]),
        .O(\sr_reg[1]_2 ));
  LUT6 #(
    .INIT(64'h4444040044444444)) 
    \sr[4]_i_26 
       (.I0(\rgf_c1bus_wb[12]_i_9_n_0 ),
        .I1(\sr[4]_i_78_n_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb_reg[12]_1 ),
        .I4(\sr[4]_i_79_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_6_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \sr[4]_i_260 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [9]),
        .O(\sr_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \sr[4]_i_262 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\i_/rgf_c1bus_wb[4]_i_86 [0]),
        .O(\sr_reg[0]_35 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \sr[4]_i_264 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [0]),
        .O(\sr_reg[1]_13 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \sr[4]_i_266 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [4]),
        .O(\sr_reg[1]_9 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \sr[4]_i_268 
       (.I0(\stat_reg[2]_14 ),
        .I1(\stat_reg[2]_15 ),
        .I2(\stat_reg[2]_16 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\i_/rgf_c1bus_wb[4]_i_96 [6]),
        .O(\sr_reg[1]_7 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \sr[4]_i_27 
       (.I0(\sr[4]_i_9_0 ),
        .I1(\sr[4]_i_81_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\sr[4]_i_82_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h3022332230223022)) 
    \sr[4]_i_28 
       (.I0(\sr[4]_i_83_n_0 ),
        .I1(\sr[4]_i_84_n_0 ),
        .I2(\sr[4]_i_85_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\rgf_c1bus_wb_reg[6]_2 ),
        .I5(\bdatw[9]_INST_0_i_16_0 ),
        .O(\sr[4]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AAFE)) 
    \sr[4]_i_29 
       (.I0(\sr[4]_i_86_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I3(\sr[4]_i_87_n_0 ),
        .I4(\sr[4]_i_88_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0100)) 
    \sr[4]_i_3 
       (.I0(\sr[4]_i_9_n_0 ),
        .I1(\sr[4]_i_10_n_0 ),
        .I2(\sr[4]_i_11_n_0 ),
        .I3(\sr[4]_i_12_n_0 ),
        .I4(\sr[4]_i_13_n_0 ),
        .I5(\sr[4]_i_14_n_0 ),
        .O(alu_sr_flag1));
  LUT6 #(
    .INIT(64'h00FF000E0000000E)) 
    \sr[4]_i_30 
       (.I0(\sr[4]_i_10_1 ),
        .I1(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I3(\sr[4]_i_90_n_0 ),
        .I4(\tr_reg[4]_0 ),
        .I5(\sr[4]_i_10_2 ),
        .O(\sr[4]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEFAAAF)) 
    \sr[4]_i_31 
       (.I0(\tr_reg[4]_0 ),
        .I1(\sr[4]_i_92_n_0 ),
        .I2(\sr[4]_i_93_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_8_n_0 ),
        .I4(\stat_reg[2]_7 ),
        .I5(\sr[4]_i_10_0 ),
        .O(\sr[4]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFFFBAAAAAAAA)) 
    \sr[4]_i_32 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\sr[4]_i_95_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .I3(\sr[4]_i_96_n_0 ),
        .I4(\rgf_c1bus_wb_reg[13]_2 ),
        .I5(\tr_reg[4]_0 ),
        .O(\sr[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAAFAAEFAAEF)) 
    \sr[4]_i_33 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_8_n_0 ),
        .O(\sr[4]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFBBBAAAAAAAA)) 
    \sr[4]_i_34 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\sr[4]_i_97_n_0 ),
        .I2(\rgf_c1bus_wb_reg[6]_2 ),
        .I3(\rgf_c1bus_wb[15]_i_14_0 ),
        .I4(\rgf_c1bus_wb[6]_i_7_n_0 ),
        .I5(\tr_reg[4]_0 ),
        .O(\sr[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF08AA)) 
    \sr[4]_i_35 
       (.I0(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .I2(\sr[4]_i_98_n_0 ),
        .I3(\sr[4]_i_99_n_0 ),
        .I4(\tr_reg[4]_0 ),
        .I5(\sr[4]_i_100_n_0 ),
        .O(\sr[4]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF8A)) 
    \sr[4]_i_36 
       (.I0(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .I1(\sr[4]_i_101_n_0 ),
        .I2(\rgf_c1bus_wb_reg[8]_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\sr[4]_i_102_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFBBBAAAAAAAA)) 
    \sr[4]_i_37 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb_reg[13]_1 ),
        .I3(\rgf_c1bus_wb[15]_i_14_0 ),
        .I4(\sr[4]_i_103_n_0 ),
        .I5(\tr_reg[4]_0 ),
        .O(\sr[4]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBAAFBAAFBAAFB)) 
    \sr[4]_i_38 
       (.I0(\tr_reg[4]_0 ),
        .I1(\sr[4]_i_104_n_0 ),
        .I2(\sr[4]_i_11_0 ),
        .I3(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I4(\stat_reg[2]_8 ),
        .I5(a1bus_0[3]),
        .O(\sr[4]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBABABBBA)) 
    \sr[4]_i_39 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_11_n_0 ),
        .I3(\sr[4]_i_106_n_0 ),
        .I4(\rgf_c1bus_wb_reg[13]_0 ),
        .I5(\sr[4]_i_107_n_0 ),
        .O(\sr[4]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAAA)) 
    \sr[4]_i_40 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[13]_1 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_108_n_0 ),
        .I4(\tr_reg[4]_0 ),
        .O(\sr[4]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF0E)) 
    \sr[4]_i_41 
       (.I0(\sr[4]_i_109_n_0 ),
        .I1(\sr[4]_i_110_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_9_n_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\sr[4]_i_111_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455555455)) 
    \sr[4]_i_42 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .I5(\sr[4]_i_112_n_0 ),
        .O(\sr[4]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_43 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\sr[4]_i_113_n_0 ),
        .I2(\sr[4]_i_114_n_0 ),
        .O(\sr[4]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAAAA)) 
    \sr[4]_i_44 
       (.I0(\tr_reg[4]_0 ),
        .I1(\rgf_c1bus_wb[2]_i_12_n_0 ),
        .I2(\sr[4]_i_12_0 ),
        .I3(\stat_reg[2]_4 ),
        .I4(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .I5(\sr[4]_i_116_n_0 ),
        .O(\sr[4]_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFEFAAAA)) 
    \sr[4]_i_45 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_7_n_0 ),
        .I3(\sr[4]_i_117_n_0 ),
        .I4(\tr_reg[4]_0 ),
        .O(\sr[4]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0404040455045555)) 
    \sr[4]_i_46 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\sr[4]_i_118_n_0 ),
        .I2(\sr[4]_i_119_n_0 ),
        .I3(\sr[4]_i_120_n_0 ),
        .I4(\sr[4]_i_121_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_4_n_0 ),
        .O(\sr[4]_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_48 
       (.I0(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .O(\sr[4]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_49 
       (.I0(\rgf_c1bus_wb[0]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I2(\sr[4]_i_124_n_0 ),
        .O(\sr[4]_i_49_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_50 
       (.I0(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_15_n_0 ),
        .O(\sr[4]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[4]_i_51 
       (.I0(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\sr[4]_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_52 
       (.I0(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[9]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb_reg[12]_i_15_n_0 ),
        .O(\sr[4]_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_53 
       (.I0(\rgf_c1bus_wb[6]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .O(\sr[4]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00AB)) 
    \sr[4]_i_54 
       (.I0(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_0 ),
        .I2(\rgf_c0bus_wb_reg[7]_1 ),
        .I3(\sr[4]_i_125_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr[4]_i_126_n_0 ),
        .O(\sr[4]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0220000)) 
    \sr[4]_i_55 
       (.I0(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I1(\sr[4]_i_127_n_0 ),
        .I2(\sr[4]_i_15_0 ),
        .I3(\tr_reg[4] ),
        .I4(\rgf_c0bus_wb[15]_i_7_0 ),
        .I5(\sr[4]_i_129_n_0 ),
        .O(\sr[4]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFF040000FFFFFFFF)) 
    \sr[4]_i_56 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\rgf_c0bus_wb[11]_i_3_0 ),
        .I2(\rgf_c0bus_wb_reg[9]_0 ),
        .I3(\rgf_c0bus_wb[1]_i_5_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c0bus_wb[15]_i_7_0 ),
        .O(\sr[4]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h0455555504040404)) 
    \sr[4]_i_58 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I3(a0bus_0[13]),
        .I4(\rgf_c0bus_wb[11]_i_3_0 ),
        .I5(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\sr[4]_i_58_n_0 ));
  LUT5 #(
    .INIT(32'h888B3333)) 
    \sr[4]_i_59 
       (.I0(\sr[4]_i_16_0 ),
        .I1(\tr_reg[4] ),
        .I2(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_0 ),
        .I4(\stat_reg[2]_10 ),
        .O(\sr[4]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000100)) 
    \sr[4]_i_6 
       (.I0(\sr[4]_i_15_n_0 ),
        .I1(\sr[4]_i_16_n_0 ),
        .I2(\sr[4]_i_17_n_0 ),
        .I3(\sr[4]_i_18_n_0 ),
        .I4(\sr[4]_i_19_n_0 ),
        .I5(\sr[4]_i_20_n_0 ),
        .O(alu_sr_flag0[0]));
  LUT6 #(
    .INIT(64'hABABABABABABABAA)) 
    \sr[4]_i_60 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[2]_i_12_n_0 ),
        .I2(\sr[4]_i_134_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_11_n_0 ),
        .O(\sr[4]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFF008A0000008A00)) 
    \sr[4]_i_61 
       (.I0(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .I1(\sr[4]_i_17_1 ),
        .I2(\sr[4]_i_136_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_7_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c0bus_wb[4]_i_2_n_0 ),
        .O(\sr[4]_i_61_n_0 ));
  LUT5 #(
    .INIT(32'hD0D000D0)) 
    \sr[4]_i_62 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\sr[4]_i_137_n_0 ),
        .I2(\tr_reg[4] ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\sr[4]_i_17_0 ),
        .O(\sr[4]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hFF5D0000FFFFFFFF)) 
    \sr[4]_i_63 
       (.I0(\sr[4]_i_18_3 ),
        .I1(\rgf_c0bus_wb_reg[10]_1 ),
        .I2(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .I4(\sr[4]_i_139_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_7_0 ),
        .O(\sr[4]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFF5D0000FFFFFFFF)) 
    \sr[4]_i_64 
       (.I0(\sr[4]_i_140_n_0 ),
        .I1(\rgf_c0bus_wb_reg[6]_1 ),
        .I2(\rgf_c0bus_wb[11]_i_11_0 ),
        .I3(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .I4(\tr_reg[4] ),
        .I5(\rgf_c0bus_wb[15]_i_7_0 ),
        .O(\sr[4]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBAAAA)) 
    \sr[4]_i_65 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\sr[4]_i_141_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_8_n_0 ),
        .O(\sr[4]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h0020F02000200020)) 
    \sr[4]_i_66 
       (.I0(\sr[4]_i_18_2 ),
        .I1(\sr[4]_i_143_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_0 ),
        .I3(\tr_reg[4] ),
        .I4(\sr[4]_i_144_n_0 ),
        .I5(\sr[4]_i_145_n_0 ),
        .O(\sr[4]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFF000E0000000E00)) 
    \sr[4]_i_67 
       (.I0(\sr[4]_i_18_0 ),
        .I1(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I2(\sr[4]_i_147_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_7_0 ),
        .I4(\tr_reg[4] ),
        .I5(\sr[4]_i_18_1 ),
        .O(\sr[4]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFBBBBAAAAAAAA)) 
    \sr[4]_i_68 
       (.I0(\tr_reg[4] ),
        .I1(\rgf_c0bus_wb[3]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_5_n_0 ),
        .O(\sr[4]_i_68_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEA)) 
    \sr[4]_i_69 
       (.I0(\rgf_c0bus_wb[9]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb_reg[7]_i_11_n_0 ),
        .O(\sr[4]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_70 
       (.I0(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .I3(\sr[4]_i_149_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_15_n_0 ),
        .I5(\sr[4]_i_150_n_0 ),
        .O(\sr[4]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_71 
       (.I0(\rgf_c0bus_wb[2]_i_13_n_0 ),
        .I1(\sr[4]_i_151_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb_reg[15]_i_3_n_0 ),
        .O(\sr[4]_i_71_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \sr[4]_i_72 
       (.I0(\rgf_c0bus_wb[13]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_19_n_0 ),
        .O(\sr[4]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEFEAEAEA)) 
    \sr[4]_i_73 
       (.I0(\sr[4]_i_20_0 ),
        .I1(\sr[4]_i_153_n_0 ),
        .I2(\stat_reg[2]_10 ),
        .I3(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\sr_reg[15]_0 [4]),
        .O(\sr[4]_i_73_n_0 ));
  LUT4 #(
    .INIT(16'h3DFD)) 
    \sr[4]_i_74 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .I2(ir1[11]),
        .I3(ir1[10]),
        .O(\sr[4]_i_74_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_75 
       (.I0(ir1[5]),
        .I1(ir1[9]),
        .O(\sr[4]_i_75_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \sr[4]_i_76 
       (.I0(ir1[12]),
        .I1(ir1[15]),
        .I2(ir1[13]),
        .O(\sr[4]_i_76_n_0 ));
  LUT5 #(
    .INIT(32'h2020202A)) 
    \sr[4]_i_77 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_25_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[6]_i_6_0 ),
        .I4(\stat_reg[1]_0 ),
        .O(\sr[4]_i_77_n_0 ));
  LUT5 #(
    .INIT(32'hFDFFCCCC)) 
    \sr[4]_i_78 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\sr[4]_i_25_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\stat_reg[2]_4 ),
        .O(\sr[4]_i_78_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_79 
       (.I0(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I1(\bdatw[9]_INST_0_i_16_0 ),
        .I2(\stat_reg[2]_8 ),
        .O(\sr[4]_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF0D0000)) 
    \sr[4]_i_8 
       (.I0(\sr[4]_i_21_n_0 ),
        .I1(\sr[4]_i_22_n_0 ),
        .I2(\sr[4]_i_23_n_0 ),
        .I3(\sr[4]_i_24_n_0 ),
        .I4(\stat[0]_i_2__1_0 ),
        .I5(\stat[2]_i_5__1_n_0 ),
        .O(ctl_sr_upd1));
  LUT6 #(
    .INIT(64'hFFFBBBFBAAAAAAAA)) 
    \sr[4]_i_81 
       (.I0(\sr[4]_i_157_n_0 ),
        .I1(\bdatw[9]_INST_0_i_16_0 ),
        .I2(\sr[4]_i_29_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[9]_i_3_1 ),
        .I5(\stat_reg[2]_4 ),
        .O(\sr[4]_i_81_n_0 ));
  LUT4 #(
    .INIT(16'h08A8)) 
    \sr[4]_i_82 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_2_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_27_0 ),
        .O(\sr[4]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA0A02AAAA0002)) 
    \sr[4]_i_83 
       (.I0(\sr[4]_i_158_n_0 ),
        .I1(\sr[4]_i_28_0 ),
        .I2(\stat_reg[1]_0 ),
        .I3(\bdatw[9]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .I5(\sr[4]_i_28_1 ),
        .O(\sr[4]_i_83_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_84 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[15]_1 ),
        .I2(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .O(\sr[4]_i_84_n_0 ));
  LUT4 #(
    .INIT(16'h5101)) 
    \sr[4]_i_85 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb_reg[7]_3 ),
        .O(\sr[4]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hCCCECCCCCCCECECE)) 
    \sr[4]_i_86 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\tr_reg[4]_0 ),
        .I2(\rgf_c1bus_wb[1]_i_12_n_0 ),
        .I3(\sr[4]_i_46_0 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\sr[4]_i_29_3 ),
        .O(\sr[4]_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFECCCCCCCC)) 
    \sr[4]_i_87 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[1]_i_12_n_0 ),
        .I2(\sr[4]_i_29_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[9]_i_3_1 ),
        .I5(\stat_reg[2]_4 ),
        .O(\sr[4]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h80AA8AAA800A8A0A)) 
    \sr[4]_i_88 
       (.I0(\tr_reg[4]_0 ),
        .I1(\sr[4]_i_29_1 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\stat_reg[2]_8 ),
        .I4(\sr[4]_i_29_2 ),
        .I5(\sr[4]_i_163_n_0 ),
        .O(\sr[4]_i_88_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEFE)) 
    \sr[4]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_4_n_0 ),
        .I2(\sr[4]_i_25_n_0 ),
        .I3(\sr[4]_i_26_n_0 ),
        .I4(\sr[4]_i_27_n_0 ),
        .I5(\sr[4]_i_28_n_0 ),
        .O(\sr[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAEFFAAAAAEAFAAAA)) 
    \sr[4]_i_90 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\sr[4]_i_30_0 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\stat_reg[2]_4 ),
        .I5(\sr[4]_i_30_1 ),
        .O(\sr[4]_i_90_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \sr[4]_i_92 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I2(\stat_reg[2]_4 ),
        .O(\sr[4]_i_92_n_0 ));
  LUT4 #(
    .INIT(16'hFD5D)) 
    \sr[4]_i_93 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\rgf_c1bus_wb[9]_i_3_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_29_3 ),
        .O(\sr[4]_i_93_n_0 ));
  LUT5 #(
    .INIT(32'hEAEFAAAA)) 
    \sr[4]_i_95 
       (.I0(\stat_reg[2]_8 ),
        .I1(\rgf_c1bus_wb[13]_i_2_0 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .O(\sr[4]_i_95_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_96 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[2]_8 ),
        .O(\sr[4]_i_96_n_0 ));
  LUT5 #(
    .INIT(32'hEAEFAAAA)) 
    \sr[4]_i_97 
       (.I0(\stat_reg[2]_8 ),
        .I1(\sr[4]_i_43_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[4]_i_43_2 ),
        .I4(\bdatw[9]_INST_0_i_16_0 ),
        .O(\sr[4]_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h1011100011111111)) 
    \sr[4]_i_98 
       (.I0(\sr[4]_i_168_n_0 ),
        .I1(\stat_reg[2]_7 ),
        .I2(\rgf_c1bus_wb_reg[11]_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb[11]_i_6_0 ),
        .I5(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .O(\sr[4]_i_98_n_0 ));
  LUT4 #(
    .INIT(16'hFD5D)) 
    \sr[4]_i_99 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[4]_i_35_1 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\sr[6]_i_6_2 ),
        .O(\sr[4]_i_99_n_0 ));
  LUT6 #(
    .INIT(64'h0000001E00E10000)) 
    \sr[5]_i_10 
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[15] ),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb_reg[15] [3]),
        .I5(a0bus_0[15]),
        .O(\sr[5]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[5]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I1(\tr_reg[4]_0 ),
        .O(\sr[5]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00090600)) 
    \sr[5]_i_8 
       (.I0(\stat_reg[2]_3 ),
        .I1(fch_leir_nir_reg),
        .I2(tout__1_carry_i_11_0),
        .I3(\rgf_c1bus_wb_reg[15] [1]),
        .I4(a1bus_0[15]),
        .O(\sr[5]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[5]_i_9 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\sr[5]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[6]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\bdatw[9]_INST_0_i_16_0 ),
        .I2(\rgf_c1bus_wb_reg[7]_2 ),
        .O(\sr[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hDF555555DF55FFFF)) 
    \sr[6]_i_11 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\stat_reg[1]_0 ),
        .I2(\sr[6]_i_6_0 ),
        .I3(\sr[6]_i_6_3 ),
        .I4(\bdatw[8]_INST_0_i_16_0 ),
        .I5(\sr[6]_i_6_2 ),
        .O(\sr[6]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFEFFAEA)) 
    \sr[6]_i_14 
       (.I0(\bbus_o[2]_INST_0_i_1_0 ),
        .I1(\sr[6]_i_18_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\sr[6]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb_reg[7]_2 ),
        .O(\sr[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h220A220A000AAA0A)) 
    \sr[6]_i_15 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[6]_i_9_1 ),
        .I2(\sr[6]_i_9_0 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\rgf_c1bus_wb_reg[3]_0 ),
        .I5(\stat_reg[1]_0 ),
        .O(\sr[6]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \sr[6]_i_18 
       (.I0(\bbus_o[0]_INST_0_i_1_0 ),
        .I1(a0bus_0[13]),
        .I2(\tr_reg[0]_0 ),
        .I3(a0bus_0[14]),
        .O(\sr[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h000000008C0FBF0F)) 
    \sr[6]_i_19 
       (.I0(\stat_reg[2]_10 ),
        .I1(\stat_reg[1]_1 ),
        .I2(a0bus_0[15]),
        .I3(\tr_reg[0]_0 ),
        .I4(\sr_reg[15]_0 [6]),
        .I5(\bbus_o[0]_INST_0_i_1_0 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h04FF)) 
    \sr[6]_i_21 
       (.I0(\bdatw[8]_INST_0_i_16_2 ),
        .I1(a1bus_0[15]),
        .I2(\stat_reg[2]_4 ),
        .I3(\stat_reg[1]_0 ),
        .O(\stat_reg[2]_13 ));
  LUT6 #(
    .INIT(64'h00000000ACAFACAC)) 
    \sr[6]_i_6 
       (.I0(\sr[6]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb_reg[15]_1 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\sr[6]_i_10_n_0 ),
        .I4(\sr[6]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h020202A2A2A2A2A2)) 
    \sr[6]_i_7 
       (.I0(\rgf_c0bus_wb[15]_i_7_0 ),
        .I1(\sr[6]_i_5 ),
        .I2(\tr_reg[4] ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\sr[4]_i_17_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\sr[6]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h00E1)) 
    \sr[6]_i_8 
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\sr[6]_i_5_0 ),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\sr[6]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h0000EEFA)) 
    \sr[6]_i_9 
       (.I0(\bdatw[9]_INST_0_i_16_0 ),
        .I1(\sr[6]_i_6_1 ),
        .I2(\rgf_c1bus_wb_reg[4]_1 ),
        .I3(\bdatw[8]_INST_0_i_16_0 ),
        .I4(\sr[6]_i_15_n_0 ),
        .O(\sr[6]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \sr[7]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[15] [3]),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(alu_sr_flag0[3]));
  LUT6 #(
    .INIT(64'h00000000F3005555)) 
    \stat[0]_i_1 
       (.I0(\stat_reg[0]_49 ),
        .I1(\stat[0]_i_3__0_n_0 ),
        .I2(\stat[0]_i_4__1_n_0 ),
        .I3(\stat_reg[0]_50 ),
        .I4(ir0[14]),
        .I5(ir0[15]),
        .O(\stat_reg[0]_4 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00D0F0F0)) 
    \stat[0]_i_10 
       (.I0(ir0[7]),
        .I1(ir0[6]),
        .I2(\ccmd[3]_INST_0_i_14_n_0 ),
        .I3(ir0[8]),
        .I4(ir0[9]),
        .I5(ir0[11]),
        .O(\stat[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0440044400000000)) 
    \stat[0]_i_10__0 
       (.I0(ir0[8]),
        .I1(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[0]),
        .I4(ir0[1]),
        .I5(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .O(\stat[0]_i_10__0_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \stat[0]_i_10__1 
       (.I0(\sr_reg[15]_0 [10]),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .O(\stat[0]_i_10__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000077F70000)) 
    \stat[0]_i_11 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .I2(\stat[0]_i_19_n_0 ),
        .I3(\stat[0]_i_20_n_0 ),
        .I4(ir0[11]),
        .I5(\stat[0]_i_21_n_0 ),
        .O(\stat[0]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_11__0 
       (.I0(ir1[10]),
        .I1(ir1[11]),
        .I2(ir1[9]),
        .I3(ir1[8]),
        .O(\stat[0]_i_11__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_11__1 
       (.I0(ir0[4]),
        .I1(ir0[6]),
        .O(\stat[0]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'hC0CCC040CCCCCC44)) 
    \stat[0]_i_12 
       (.I0(ir0[11]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(\stat[0]_i_22_n_0 ),
        .I3(brdy),
        .I4(ir0[8]),
        .I5(\stat[0]_i_23__0_n_0 ),
        .O(\stat[0]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF12F)) 
    \stat[0]_i_12__1 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(ir1[0]),
        .I3(ir1[2]),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .O(\stat[0]_i_12__1_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAAAEA)) 
    \stat[0]_i_13 
       (.I0(\stat[0]_i_24_n_0 ),
        .I1(\stat[0]_i_25_n_0 ),
        .I2(\stat[0]_i_26_n_0 ),
        .I3(ir0[11]),
        .I4(\stat[0]_i_27_n_0 ),
        .O(\stat[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \stat[0]_i_13__0 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .I2(ir1[7]),
        .I3(ir1[3]),
        .I4(ir1[1]),
        .I5(ir1[6]),
        .O(\stat[0]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFFFFFFF)) 
    \stat[0]_i_14 
       (.I0(ir1[3]),
        .I1(ir1[1]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[4]),
        .I4(ir1[6]),
        .I5(\fadr[15]_INST_0_i_16_n_0 ),
        .O(\stat[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFEFEFEEEEEEEE)) 
    \stat[0]_i_14__0 
       (.I0(\stat[0]_i_28__0_n_0 ),
        .I1(ir0[2]),
        .I2(ir0[0]),
        .I3(ir0[1]),
        .I4(\iv_reg[15]_0 [0]),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\stat[0]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000100)) 
    \stat[0]_i_15 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(ir0[11]),
        .I2(\stat[0]_i_8_0 ),
        .I3(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I4(\bdatw[10]_INST_0_i_18_n_0 ),
        .I5(\stat[0]_i_30_n_0 ),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0020202000200000)) 
    \stat[0]_i_15__0 
       (.I0(\stat[0]_i_18__0_n_0 ),
        .I1(\stat[0]_i_19__0_n_0 ),
        .I2(\stat[0]_i_20__0_n_0 ),
        .I3(\stat[0]_i_21__0_n_0 ),
        .I4(ir1[11]),
        .I5(\stat[0]_i_22__0_n_0 ),
        .O(\stat[0]_i_15__0_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \stat[0]_i_16 
       (.I0(ir0[8]),
        .I1(crdy),
        .I2(ir0[9]),
        .O(\stat[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00AE00AE000000AE)) 
    \stat[0]_i_16__0 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(\badrx[15]_INST_0_i_5_n_0 ),
        .I2(\stat[0]_i_24__0_n_0 ),
        .I3(\stat[0]_i_25__0_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\stat[0]_i_26__0_n_0 ),
        .O(\stat[0]_i_16__0_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \stat[0]_i_17 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[6]),
        .I3(brdy),
        .O(\stat[0]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_17__0 
       (.I0(ir1[11]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .O(\stat[0]_i_17__0_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_18 
       (.I0(ir0[9]),
        .I1(ir0[7]),
        .O(\stat[0]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \stat[0]_i_18__0 
       (.I0(ir1[8]),
        .I1(\stat_reg[0]_48 ),
        .I2(brdy),
        .O(\stat[0]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'hF2FF3333FFFFFFFF)) 
    \stat[0]_i_19 
       (.I0(ir0[3]),
        .I1(brdy),
        .I2(ir0[4]),
        .I3(ir0[7]),
        .I4(ir0[10]),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\stat[0]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h2AAAAAAA)) 
    \stat[0]_i_19__0 
       (.I0(ir1[6]),
        .I1(ir1[5]),
        .I2(ir1[7]),
        .I3(ir1[10]),
        .I4(ir1[3]),
        .O(\stat[0]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45454544)) 
    \stat[0]_i_1__2 
       (.I0(\stat[0]_i_2__1_n_0 ),
        .I1(\stat_reg[0]_53 ),
        .I2(\stat[0]_i_3__1_n_0 ),
        .I3(\stat[0]_i_4__0_n_0 ),
        .I4(\stat[0]_i_5__0_n_0 ),
        .I5(\stat[0]_i_6_n_0 ),
        .O(\stat_reg[2]_12 [0]));
  LUT6 #(
    .INIT(64'h8000000000880088)) 
    \stat[0]_i_20 
       (.I0(ir0[5]),
        .I1(brdy),
        .I2(ir0[7]),
        .I3(ir0[6]),
        .I4(ir0[3]),
        .I5(ir0[10]),
        .O(\stat[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_20__0 
       (.I0(ir1[9]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .O(\stat[0]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'h4044404440000000)) 
    \stat[0]_i_21 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .I2(crdy),
        .I3(ir0[8]),
        .I4(\sr_reg[15]_0 [11]),
        .I5(ir0[7]),
        .O(\stat[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h4444444444044444)) 
    \stat[0]_i_21__0 
       (.I0(ir1[6]),
        .I1(ir1[10]),
        .I2(ir1[7]),
        .I3(ir1[4]),
        .I4(ir1[3]),
        .I5(ir1[5]),
        .O(\stat[0]_i_21__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_22 
       (.I0(ir0[5]),
        .I1(ir0[3]),
        .O(\stat[0]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_22__0 
       (.I0(ir1[10]),
        .I1(ir1[6]),
        .O(\stat[0]_i_22__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000EA00FFFFFFFF)) 
    \stat[0]_i_23 
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(\sr_reg[15]_0 [11]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(ir1[11]),
        .O(\stat[0]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \stat[0]_i_23__0 
       (.I0(ir0[9]),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .O(\stat[0]_i_23__0_n_0 ));
  LUT6 #(
    .INIT(64'h00AA00AA00EB00AA)) 
    \stat[0]_i_24 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(ir0[8]),
        .I2(ir0[11]),
        .I3(crdy),
        .I4(ir0[7]),
        .I5(\ccmd[4]_INST_0_i_20_n_0 ),
        .O(\stat[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h000000007CFCFFFF)) 
    \stat[0]_i_24__0 
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(ir1[10]),
        .I3(ir1[3]),
        .I4(\rgf_selc1_rn_wb_reg[2] ),
        .I5(\stat[0]_i_27__0_n_0 ),
        .O(\stat[0]_i_24__0_n_0 ));
  LUT5 #(
    .INIT(32'h8000FFFF)) 
    \stat[0]_i_25 
       (.I0(ir0[10]),
        .I1(ir0[7]),
        .I2(ir0[5]),
        .I3(ir0[3]),
        .I4(ir0[6]),
        .O(\stat[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00A000AF00A000BF)) 
    \stat[0]_i_25__0 
       (.I0(\stat[0]_i_28_n_0 ),
        .I1(\bdatw[15]_INST_0_i_197_n_0 ),
        .I2(ir1[10]),
        .I3(ir1[11]),
        .I4(\stat[0]_i_29_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .O(\stat[0]_i_25__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000DC0000000000)) 
    \stat[0]_i_26 
       (.I0(ir0[6]),
        .I1(ir0[11]),
        .I2(ir0[10]),
        .I3(ir0[8]),
        .I4(brdy),
        .I5(ir0[9]),
        .O(\stat[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00004000F0F040F0)) 
    \stat[0]_i_26__0 
       (.I0(\stat[0]_i_30__0_n_0 ),
        .I1(\stat[0]_i_31__0_n_0 ),
        .I2(ir1[11]),
        .I3(brdy),
        .I4(\stat_reg[0]_48 ),
        .I5(ir1[8]),
        .O(\stat[0]_i_26__0_n_0 ));
  LUT6 #(
    .INIT(64'hDDDFDDDDDDDDDDDD)) 
    \stat[0]_i_27 
       (.I0(ir0[10]),
        .I1(ir0[6]),
        .I2(ir0[5]),
        .I3(ir0[4]),
        .I4(ir0[7]),
        .I5(ir0[3]),
        .O(\stat[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h5D000C0C00000000)) 
    \stat[0]_i_27__0 
       (.I0(ir1[3]),
        .I1(brdy),
        .I2(\stat_reg[0]_48 ),
        .I3(\stat[0]_i_32__0_n_0 ),
        .I4(ir1[10]),
        .I5(\stat[0]_i_33__0_n_0 ),
        .O(\stat[0]_i_27__0_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \stat[0]_i_28 
       (.I0(\sr_reg[15]_0 [11]),
        .I1(ir1[9]),
        .I2(ir1[7]),
        .O(\stat[0]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_28__0 
       (.I0(ir0[11]),
        .I1(\rgf_selc0_rn_wb_reg[0] [2]),
        .O(\stat[0]_i_28__0_n_0 ));
  LUT5 #(
    .INIT(32'h40CC44CC)) 
    \stat[0]_i_29 
       (.I0(ir1[8]),
        .I1(rst_n_fl_reg_9),
        .I2(ir1[6]),
        .I3(ir1[9]),
        .I4(ir1[7]),
        .O(\stat[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h1100110000000001)) 
    \stat[0]_i_2__0 
       (.I0(ir0[8]),
        .I1(ir0[9]),
        .I2(ir0[5]),
        .I3(ir0[11]),
        .I4(ir0[3]),
        .I5(ir0[7]),
        .O(\stat[0]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h008A0000000000FF)) 
    \stat[0]_i_2__1 
       (.I0(ir1[0]),
        .I1(ir1[1]),
        .I2(\iv_reg[15]_0 [0]),
        .I3(\stat[0]_i_7__0_n_0 ),
        .I4(\stat_reg[0]_55 ),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(\stat[0]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000FB)) 
    \stat[0]_i_30 
       (.I0(ir0[2]),
        .I1(\rgf_selc0_rn_wb_reg[0]_0 ),
        .I2(fch_irq_req),
        .I3(\stat[0]_i_31_n_0 ),
        .I4(\stat[0]_i_15_0 ),
        .I5(\stat[0]_i_33_n_0 ),
        .O(\stat[0]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[0]_i_30__0 
       (.I0(ir1[10]),
        .I1(ir1[9]),
        .O(\stat[0]_i_30__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF21FF)) 
    \stat[0]_i_31 
       (.I0(ir0[3]),
        .I1(ir0[1]),
        .I2(ir0[0]),
        .I3(\stat[0]_i_34_n_0 ),
        .I4(\bcmd[0]_INST_0_i_22_n_0 ),
        .I5(\stat[0]_i_30_0 ),
        .O(\stat[0]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_31__0 
       (.I0(ir1[3]),
        .I1(ir1[5]),
        .O(\stat[0]_i_31__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_32__0 
       (.I0(ir1[7]),
        .I1(ir1[4]),
        .O(\stat[0]_i_32__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \stat[0]_i_33 
       (.I0(\rgf_selc0_rn_wb_reg[0] [0]),
        .I1(ir0[2]),
        .I2(ir0[10]),
        .I3(ir0[9]),
        .I4(ir0[6]),
        .I5(\bdatw[10]_INST_0_i_18_n_0 ),
        .O(\stat[0]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_33__0 
       (.I0(ir1[5]),
        .I1(ir1[6]),
        .O(\stat[0]_i_33__0_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_34 
       (.I0(ir0[8]),
        .I1(ir0[7]),
        .O(\stat[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8778)) 
    \stat[0]_i_3__0 
       (.I0(ir0[12]),
        .I1(\sr_reg[15]_0 [7]),
        .I2(\sr_reg[15]_0 [5]),
        .I3(ir0[11]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(ir0[13]),
        .O(\stat[0]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFDDCCFC)) 
    \stat[0]_i_3__1 
       (.I0(\stat[0]_i_8__1_n_0 ),
        .I1(\stat[0]_i_9__0_n_0 ),
        .I2(\stat[0]_i_10__1_n_0 ),
        .I3(ir1[1]),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(\stat[0]_i_11__0_n_0 ),
        .O(\stat[0]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h67FF0000FFFFFFFF)) 
    \stat[0]_i_3__2 
       (.I0(ir0[5]),
        .I1(ir0[6]),
        .I2(ir0[3]),
        .I3(ir0[7]),
        .I4(\stat[0]_i_7_n_0 ),
        .I5(\stat[2]_i_12_n_0 ),
        .O(\stat[0]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEFEE)) 
    \stat[0]_i_4 
       (.I0(\stat[0]_i_8__0_n_0 ),
        .I1(\stat_reg[0]_52 ),
        .I2(ir0[7]),
        .I3(ir0[2]),
        .I4(ir0[8]),
        .I5(\stat[0]_i_10__0_n_0 ),
        .O(\stat[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000033332)) 
    \stat[0]_i_4__0 
       (.I0(fch_irq_req),
        .I1(\stat[0]_i_12__1_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[2]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\stat[0]_i_13__0_n_0 ),
        .O(\stat[0]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h5555005400000054)) 
    \stat[0]_i_4__1 
       (.I0(\bcmd[2]_INST_0_i_9_n_0 ),
        .I1(\stat[0]_i_9_n_0 ),
        .I2(\stat[0]_i_10_n_0 ),
        .I3(\stat[0]_i_11_n_0 ),
        .I4(\stat[0]_i_12_n_0 ),
        .I5(\stat[0]_i_13_n_0 ),
        .O(\stat[0]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'hB5BFB5BFF7FFF7AA)) 
    \stat[0]_i_5 
       (.I0(ir0[9]),
        .I1(ir0[11]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[12]),
        .I4(ir0[6]),
        .I5(ir0[10]),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000000E3E0E1E)) 
    \stat[0]_i_5__0 
       (.I0(ir1[1]),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(ir1[2]),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(\sr_reg[15]_0 [10]),
        .I5(\stat[0]_i_14_n_0 ),
        .O(\stat[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFE00000000000)) 
    \stat[0]_i_6 
       (.I0(\stat[0]_i_15__0_n_0 ),
        .I1(\stat[0]_i_16__0_n_0 ),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(\stat_reg[0]_16 ),
        .I5(\stat_reg[0]_54 ),
        .O(\stat[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hBBABAAAAAAAABBAB)) 
    \stat[0]_i_6__1 
       (.I0(\sr_reg[4]_0 ),
        .I1(\stat[0]_i_14__0_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(ir0[1]),
        .I4(brdy),
        .I5(\rgf_selc0_rn_wb_reg[0] [0]),
        .O(\stat_reg[1]_7 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_7 
       (.I0(ir0[11]),
        .I1(ir0[10]),
        .O(\stat[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFDCFFDCFFFFFFDC)) 
    \stat[0]_i_7__0 
       (.I0(ir1[1]),
        .I1(ir1[2]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\stat[0]_i_17__0_n_0 ),
        .I4(\stat[0]_i_2__1_0 ),
        .I5(\stat[2]_i_2__1 ),
        .O(\stat[0]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h20222A2222222A22)) 
    \stat[0]_i_8 
       (.I0(\stat[0]_i_15_n_0 ),
        .I1(\rgf_selc0_rn_wb_reg[0] [2]),
        .I2(ir0[1]),
        .I3(ir0[0]),
        .I4(ir0[3]),
        .I5(\sr_reg[15]_0 [10]),
        .O(\stat_reg[2]_11 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4040FF40)) 
    \stat[0]_i_8__0 
       (.I0(\bcmd[2]_INST_0_i_11_n_0 ),
        .I1(\ccmd[4]_INST_0_i_20_n_0 ),
        .I2(\stat[0]_i_11__1_n_0 ),
        .I3(\bcmd[2]_INST_0_i_9_n_0 ),
        .I4(\stat[1]_i_9__0_n_0 ),
        .I5(\sp[15]_i_8_0 ),
        .O(\stat[0]_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_8__1 
       (.I0(ir1[0]),
        .I1(ir1[3]),
        .O(\stat[0]_i_8__1_n_0 ));
  LUT6 #(
    .INIT(64'h5700570000005700)) 
    \stat[0]_i_9 
       (.I0(\stat[0]_i_16_n_0 ),
        .I1(fctl_n_91),
        .I2(\stat[0]_i_17_n_0 ),
        .I3(ir0[10]),
        .I4(\sr_reg[15]_0 [11]),
        .I5(\stat[0]_i_18_n_0 ),
        .O(\stat[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFEFEFEFE)) 
    \stat[0]_i_9__0 
       (.I0(ir1[14]),
        .I1(ir1[13]),
        .I2(ir1[15]),
        .I3(\sr_reg[15]_0 [4]),
        .I4(ir1[11]),
        .I5(ir1[12]),
        .O(\stat[0]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAEA0000)) 
    \stat[1]_i_10 
       (.I0(\stat[1]_i_12__0_n_0 ),
        .I1(\sr_reg[15]_0 [10]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(\ccmd[4]_INST_0_i_17_n_0 ),
        .I4(ir0[8]),
        .I5(\rgf_selc0_rn_wb_reg[0] [1]),
        .O(\stat[1]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEFCCEECC)) 
    \stat[1]_i_10__0 
       (.I0(ir1[0]),
        .I1(ir1[9]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[3]),
        .I4(\sr_reg[15]_0 [10]),
        .O(\stat[1]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF000400)) 
    \stat[1]_i_11 
       (.I0(ir0[6]),
        .I1(ir0[9]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[7]),
        .I4(ir0[10]),
        .I5(\stat[1]_i_13_n_0 ),
        .O(\stat[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[1]_i_11__0 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(ir1[12]),
        .O(\stat[1]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8FFF)) 
    \stat[1]_i_12 
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\stat[1]_i_17_n_0 ),
        .I2(\fadr[15]_INST_0_i_16_n_0 ),
        .I3(\stat[2]_i_5__1_n_0 ),
        .I4(ir1[4]),
        .I5(ir1[6]),
        .O(\stat[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000090)) 
    \stat[1]_i_12__0 
       (.I0(ir0[3]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(ir0[9]),
        .I3(ir0[6]),
        .I4(ir0[5]),
        .I5(ir0[4]),
        .O(\stat[1]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFDFFFDFFFD)) 
    \stat[1]_i_13 
       (.I0(\stat[1]_i_14_n_0 ),
        .I1(\bdatw[15]_INST_0_i_223_n_0 ),
        .I2(ir0[11]),
        .I3(\bcmd[2]_INST_0_i_9_n_0 ),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\sr_reg[15]_0 [10]),
        .O(\stat[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0100001001000100)) 
    \stat[1]_i_13__0 
       (.I0(ir1[9]),
        .I1(\stat[1]_i_18_n_0 ),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(\stat_reg[0]_48 ),
        .I5(brdy),
        .O(\stat[1]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[1]_i_14 
       (.I0(ir0[9]),
        .I1(ir0[10]),
        .O(\stat[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hDDD1FFFFDDDDFFF3)) 
    \stat[1]_i_14__0 
       (.I0(\sr_reg[15]_0 [10]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(\stat[2]_i_10__0_n_0 ),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(ir1[3]),
        .O(\stat[1]_i_14__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[1]_i_15 
       (.I0(ir1[10]),
        .I1(ir1[7]),
        .O(\stat[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDFFFDFFFDF)) 
    \stat[1]_i_16 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(ir1[8]),
        .I2(ir1[7]),
        .I3(ir1[11]),
        .I4(\rgf_selc1_wb_reg[1] [0]),
        .I5(\sr_reg[15]_0 [10]),
        .O(\stat[1]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[1]_i_17 
       (.I0(ir1[1]),
        .I1(ir1[0]),
        .I2(ir1[3]),
        .O(\stat[1]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[1]_i_18 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .O(\stat[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h000F00DD000000DD)) 
    \stat[1]_i_1__0 
       (.I0(\stat_reg[1]_8 ),
        .I1(\stat[1]_i_2__0_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [2]),
        .I3(ir0[15]),
        .I4(ir0[14]),
        .I5(\stat[1]_i_3_n_0 ),
        .O(\stat_reg[0]_4 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFF0101FF01)) 
    \stat[1]_i_1__1 
       (.I0(\stat[1]_i_2__1_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [2]),
        .I2(\bcmd[2]_INST_0_i_7_n_0 ),
        .I3(\stat[1]_i_3__0_n_0 ),
        .I4(\stat[1]_i_4__0_n_0 ),
        .I5(\stat_reg[0]_53 ),
        .O(\stat_reg[2]_12 [1]));
  LUT6 #(
    .INIT(64'h0426000000000000)) 
    \stat[1]_i_2__0 
       (.I0(\rgf_selc0_rn_wb_reg[0] [1]),
        .I1(\rgf_selc0_rn_wb_reg[0] [0]),
        .I2(\stat[1]_i_4__1_n_0 ),
        .I3(\stat[1]_i_5__0_n_0 ),
        .I4(\stat[1]_i_6_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_6_n_0 ),
        .O(\stat[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000AAA82220AAA8)) 
    \stat[1]_i_2__1 
       (.I0(\stat[1]_i_5_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\stat[1]_i_6__0_n_0 ),
        .I4(\stat[1]_i_7__0_n_0 ),
        .I5(rst_n_fl_reg_9),
        .O(\stat[1]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF20000000)) 
    \stat[1]_i_3 
       (.I0(ir0[11]),
        .I1(\bcmd[2]_INST_0_i_9_n_0 ),
        .I2(ir0[7]),
        .I3(ir0[10]),
        .I4(\stat[1]_i_7_n_0 ),
        .I5(\stat[1]_i_8_n_0 ),
        .O(\stat[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0044034403440044)) 
    \stat[1]_i_3__0 
       (.I0(\stat[1]_i_9_n_0 ),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\rgf_selc1_wb_reg[1] [2]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ir1[0]),
        .I5(ir1[2]),
        .O(\stat[1]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \stat[1]_i_4__0 
       (.I0(\stat[1]_i_10__0_n_0 ),
        .I1(\stat[1]_i_11__0_n_0 ),
        .I2(\bdatw[14]_INST_0_i_29_n_0 ),
        .I3(ir1[8]),
        .I4(ir1[10]),
        .I5(\stat[1]_i_12_n_0 ),
        .O(\stat[1]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFCCCC55FFFF0C77)) 
    \stat[1]_i_4__1 
       (.I0(brdy),
        .I1(ir0[1]),
        .I2(\sr_reg[15]_0 [10]),
        .I3(ir0[2]),
        .I4(\rgf_selc0_rn_wb_reg[0] [2]),
        .I5(ir0[0]),
        .O(\stat[1]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h5551FFFFFFFFFFFF)) 
    \stat[1]_i_5 
       (.I0(\stat[1]_i_13__0_n_0 ),
        .I1(ir1[8]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\stat[1]_i_14__0_n_0 ),
        .I4(\stat[2]_i_9__0_n_0 ),
        .I5(\stat[1]_i_15_n_0 ),
        .O(\stat[1]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hEB)) 
    \stat[1]_i_5__0 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(ir0[0]),
        .I2(ir0[2]),
        .O(\stat[1]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h222822222228222A)) 
    \stat[1]_i_6 
       (.I0(\stat[1]_i_9__0_n_0 ),
        .I1(ir0[3]),
        .I2(ir0[0]),
        .I3(ir0[1]),
        .I4(\rgf_selc0_rn_wb_reg[0] [1]),
        .I5(\sr_reg[15]_0 [10]),
        .O(\stat[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEABFBFEA)) 
    \stat[1]_i_6__0 
       (.I0(ir1[13]),
        .I1(\sr_reg[15]_0 [7]),
        .I2(ir1[12]),
        .I3(\sr_reg[15]_0 [5]),
        .I4(ir1[11]),
        .O(\stat[1]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00400400)) 
    \stat[1]_i_7 
       (.I0(ir0[6]),
        .I1(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I2(brdy),
        .I3(\rgf_selc0_rn_wb_reg[0] [1]),
        .I4(\rgf_selc0_rn_wb_reg[0] [0]),
        .I5(\stat[1]_i_10_n_0 ),
        .O(\stat[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000F00010000)) 
    \stat[1]_i_7__0 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[6]),
        .I2(\stat[1]_i_16_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ir1[9]),
        .I5(ir1[10]),
        .O(\stat[1]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h0D0D0D050DFD0D05)) 
    \stat[1]_i_8 
       (.I0(\stat[0]_i_3__0_n_0 ),
        .I1(\stat[1]_i_11_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [1]),
        .I3(\rgf_selc0_rn_wb_reg[0] [0]),
        .I4(\ccmd[4]_INST_0_i_12_n_0 ),
        .I5(crdy),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \stat[1]_i_8__0 
       (.I0(ir1[15]),
        .I1(ir1[14]),
        .I2(ir1[12]),
        .I3(ir1[13]),
        .I4(ir1[10]),
        .I5(ir1[11]),
        .O(rst_n_fl_reg_9));
  LUT6 #(
    .INIT(64'hFFCFC403FFCFF733)) 
    \stat[1]_i_9 
       (.I0(\sr_reg[15]_0 [10]),
        .I1(ir1[2]),
        .I2(ir1[0]),
        .I3(ir1[1]),
        .I4(\rgf_selc1_wb_reg[1] [2]),
        .I5(\stat_reg[0]_55 ),
        .O(\stat[1]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[1]_i_9__0 
       (.I0(ir0[12]),
        .I1(ir0[11]),
        .I2(ir0[13]),
        .O(\stat[1]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000007)) 
    \stat[2]_i_10 
       (.I0(\rgf_selc0_rn_wb_reg[0] [2]),
        .I1(\rgf_selc0_rn_wb_reg[0] [1]),
        .I2(ir0[9]),
        .I3(ir0[10]),
        .I4(ir0[4]),
        .I5(ir0[2]),
        .O(\stat[2]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[2]_i_10__0 
       (.I0(ir1[5]),
        .I1(ir1[4]),
        .O(\stat[2]_i_10__0_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[2]_i_11 
       (.I0(ir1[8]),
        .I1(ir1[7]),
        .O(\stat[2]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[2]_i_12 
       (.I0(ir0[9]),
        .I1(ir0[8]),
        .O(\stat[2]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \stat[2]_i_12__0 
       (.I0(ir1[6]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .O(\stat[2]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \stat[2]_i_13 
       (.I0(\bcmd[0]_INST_0_i_22_n_0 ),
        .I1(ir0[7]),
        .I2(ir0[13]),
        .I3(ir0[11]),
        .I4(ir0[6]),
        .I5(ir0[10]),
        .O(\stat[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \stat[2]_i_13__0 
       (.I0(ir1[8]),
        .I1(ir1[6]),
        .I2(\fadr[15]_INST_0_i_16_n_0 ),
        .I3(\stat[2]_i_5__1_n_0 ),
        .I4(ir1[12]),
        .I5(ir1[13]),
        .O(\stat[2]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_14 
       (.I0(ir1[4]),
        .I1(ir1[3]),
        .O(\stat[2]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[2]_i_15 
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[10]),
        .O(\stat[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000000000F00DDDD)) 
    \stat[2]_i_2__0 
       (.I0(\stat_reg[1]_8 ),
        .I1(\stat[2]_i_4__0_n_0 ),
        .I2(\stat[2]_i_5_n_0 ),
        .I3(\stat_reg[0]_50 ),
        .I4(ir0[14]),
        .I5(ir0[15]),
        .O(\stat_reg[0]_4 [2]));
  LUT6 #(
    .INIT(64'h0000000000440040)) 
    \stat[2]_i_4__0 
       (.I0(\stat[2]_i_9_n_0 ),
        .I1(\stat[2]_i_10_n_0 ),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[3]),
        .I4(ir0[0]),
        .I5(\stat_reg[2]_21 ),
        .O(\stat[2]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h0111100010000111)) 
    \stat[2]_i_4__1 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[13]),
        .I2(\sr_reg[15]_0 [7]),
        .I3(ir1[12]),
        .I4(\sr_reg[15]_0 [5]),
        .I5(ir1[11]),
        .O(\stat_reg[0]_16 ));
  LUT6 #(
    .INIT(64'h28AAAAAAAAAAAAAA)) 
    \stat[2]_i_5 
       (.I0(\stat[0]_i_3__0_n_0 ),
        .I1(ir0[3]),
        .I2(\rgf_selc0_rn_wb_reg[0] [0]),
        .I3(ir0[12]),
        .I4(\stat[2]_i_12_n_0 ),
        .I5(\stat[2]_i_13_n_0 ),
        .O(\stat[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF6FFFFFFFFF)) 
    \stat[2]_i_5__0 
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(ir1[3]),
        .I2(\stat[2]_i_9__0_n_0 ),
        .I3(\stat[2]_i_10__0_n_0 ),
        .I4(\stat[2]_i_11_n_0 ),
        .I5(\stat[2]_i_12__0_n_0 ),
        .O(\stat_reg[0]_17 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_5__1 
       (.I0(ir1[14]),
        .I1(ir1[15]),
        .O(\stat[2]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hDDDFFFFFFFFFFFFF)) 
    \stat[2]_i_6__0 
       (.I0(\stat[2]_i_13__0_n_0 ),
        .I1(ir1[2]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[0]),
        .I4(\stat[2]_i_14_n_0 ),
        .I5(\stat[2]_i_15_n_0 ),
        .O(\stat_reg[0]_18 ));
  LUT5 #(
    .INIT(32'hBBBBBBB0)) 
    \stat[2]_i_8 
       (.I0(\stat[0]_i_9__0_n_0 ),
        .I1(ir1[11]),
        .I2(\stat[2]_i_2__1 ),
        .I3(ir1[14]),
        .I4(ir1[15]),
        .O(\sr_reg[4] ));
  LUT4 #(
    .INIT(16'hDFCC)) 
    \stat[2]_i_8__0 
       (.I0(\sr_reg[15]_0 [4]),
        .I1(ir0[13]),
        .I2(ir0[11]),
        .I3(ir0[12]),
        .O(\sr_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[2]_i_9 
       (.I0(ir0[6]),
        .I1(ir0[5]),
        .I2(ir0[8]),
        .I3(ir0[7]),
        .I4(\ccmd[1]_INST_0_i_9_n_0 ),
        .I5(ir0[12]),
        .O(\stat[2]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \stat[2]_i_9__0 
       (.I0(ir1[13]),
        .I1(ir1[11]),
        .I2(ir1[12]),
        .O(\stat[2]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__0_i_1
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bbus_o_6_sn_1),
        .I3(a0bus_0[6]),
        .O(\badr[6]_INST_0_i_2 [3]));
  LUT4 #(
    .INIT(16'hE100)) 
    tout__1_carry__0_i_2
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\rgf_c0bus_wb_reg[5] ),
        .I3(a0bus_0[5]),
        .O(\badr[6]_INST_0_i_2 [2]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__0_i_3
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\tr_reg[4] ),
        .I3(a0bus_0[4]),
        .O(\badr[6]_INST_0_i_2 [1]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_3__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\tr_reg[4]_0 ),
        .I2(a1bus_0[4]),
        .O(\badr[4]_INST_0_i_1 [1]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__0_i_4
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[3]),
        .O(\badr[6]_INST_0_i_2 [0]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_4__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[3]),
        .O(\badr[4]_INST_0_i_1 [0]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__0_i_5
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bbus_o_7_sn_1),
        .I3(a0bus_0[7]),
        .I4(\badr[6]_INST_0_i_2 [3]),
        .O(tout__1_carry__0_i_1_0[3]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__0_i_6
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bbus_o_6_sn_1),
        .I3(a0bus_0[6]),
        .I4(\badr[6]_INST_0_i_2 [2]),
        .O(tout__1_carry__0_i_1_0[2]));
  LUT5 #(
    .INIT(32'hE11E1EE1)) 
    tout__1_carry__0_i_7
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\rgf_c0bus_wb_reg[5] ),
        .I3(a0bus_0[5]),
        .I4(\badr[6]_INST_0_i_2 [1]),
        .O(tout__1_carry__0_i_1_0[1]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_7__0
       (.I0(\stat_reg[2]_3 ),
        .I1(tout__1_carry__0),
        .I2(a1bus_0[5]),
        .I3(\badr[4]_INST_0_i_1 [1]),
        .O(tout__1_carry__0_i_3__0_0[1]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__0_i_8
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\tr_reg[4] ),
        .I3(a0bus_0[4]),
        .I4(\badr[6]_INST_0_i_2 [0]),
        .O(tout__1_carry__0_i_1_0[0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_8__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\tr_reg[4]_0 ),
        .I2(a1bus_0[4]),
        .I3(\badr[4]_INST_0_i_1 [0]),
        .O(tout__1_carry__0_i_3__0_0[0]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__1_i_1
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[10]_0 ),
        .I3(a0bus_0[10]),
        .O(\badr[10]_INST_0_i_2 [3]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__1_i_2
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bdatw_9_sn_1),
        .I3(a0bus_0[9]),
        .O(\badr[10]_INST_0_i_2 [2]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__1_i_3
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[8]_0 ),
        .I3(a0bus_0[8]),
        .O(\badr[10]_INST_0_i_2 [1]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__1_i_4
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bbus_o_7_sn_1),
        .I3(a0bus_0[7]),
        .O(\badr[10]_INST_0_i_2 [0]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__1_i_5
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bdatw_11_sn_1),
        .I3(a0bus_0[11]),
        .I4(\badr[10]_INST_0_i_2 [3]),
        .O(tout__1_carry__1_i_1_0[3]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__1_i_6
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[10]_0 ),
        .I3(a0bus_0[10]),
        .I4(\badr[10]_INST_0_i_2 [2]),
        .O(tout__1_carry__1_i_1_0[2]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__1_i_7
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bdatw_9_sn_1),
        .I3(a0bus_0[9]),
        .I4(\badr[10]_INST_0_i_2 [1]),
        .O(tout__1_carry__1_i_1_0[1]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__1_i_8
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[8]_0 ),
        .I3(a0bus_0[8]),
        .I4(\badr[10]_INST_0_i_2 [0]),
        .O(tout__1_carry__1_i_1_0[0]));
  LUT3 #(
    .INIT(8'h69)) 
    tout__1_carry__2_i_1
       (.I0(\stat_reg[2]_3 ),
        .I1(fch_leir_nir_reg),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1_1 ));
  LUT4 #(
    .INIT(16'hE11E)) 
    tout__1_carry__2_i_1__0
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[15] ),
        .I3(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_2_0 [3]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__2_i_2
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bbus_o_13_sn_1),
        .I3(a0bus_0[13]),
        .O(\badr[15]_INST_0_i_2_0 [2]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__2_i_3
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bdatw_12_sn_1),
        .I3(a0bus_0[12]),
        .O(\badr[15]_INST_0_i_2_0 [1]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry__2_i_4
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bdatw_11_sn_1),
        .I3(a0bus_0[11]),
        .O(\badr[15]_INST_0_i_2_0 [0]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__2_i_6__0
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bbus_o_14_sn_1),
        .I3(\badr[15]_INST_0_i_2_0 [2]),
        .I4(a0bus_0[14]),
        .O(\badr[14]_INST_0_i_2 [2]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__2_i_7
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bbus_o_13_sn_1),
        .I3(a0bus_0[13]),
        .I4(\badr[15]_INST_0_i_2_0 [1]),
        .O(\badr[14]_INST_0_i_2 [1]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry__2_i_8
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(bdatw_12_sn_1),
        .I3(a0bus_0[12]),
        .I4(\badr[15]_INST_0_i_2_0 [0]),
        .O(\badr[14]_INST_0_i_2 [0]));
  LUT3 #(
    .INIT(8'h9F)) 
    tout__1_carry__3_i_1
       (.I0(\stat_reg[2]_3 ),
        .I1(fch_leir_nir_reg),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1_0 ));
  LUT4 #(
    .INIT(16'h1EFF)) 
    tout__1_carry__3_i_1__0
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[15] ),
        .I3(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_2_1 ));
  LUT3 #(
    .INIT(8'h96)) 
    tout__1_carry__3_i_2
       (.I0(\stat_reg[2]_3 ),
        .I1(fch_leir_nir_reg),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1 [1]));
  LUT4 #(
    .INIT(16'h1EE1)) 
    tout__1_carry__3_i_2__0
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[15] ),
        .I3(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_2_2 [1]));
  LUT3 #(
    .INIT(8'hF9)) 
    tout__1_carry__3_i_3
       (.I0(\stat_reg[2]_3 ),
        .I1(fch_leir_nir_reg),
        .I2(a1bus_0[15]),
        .O(\badr[15]_INST_0_i_1 [0]));
  LUT4 #(
    .INIT(16'hFF1E)) 
    tout__1_carry__3_i_3__0
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bdatw[15] ),
        .I3(a0bus_0[15]),
        .O(\badr[15]_INST_0_i_2_2 [0]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry_i_1
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[2]),
        .O(\badr[2]_INST_0_i_2 [2]));
  LUT3 #(
    .INIT(8'h01)) 
    tout__1_carry_i_10
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(tout__1_carry_i_13_n_0),
        .I2(tout__1_carry_i_14_n_0),
        .O(\stat_reg[2]_4 ));
  LUT4 #(
    .INIT(16'h000E)) 
    tout__1_carry_i_11
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .O(tout__1_carry_i_11_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    tout__1_carry_i_12
       (.I0(\stat_reg[2]_3 ),
        .I1(\tr_reg[0] ),
        .O(tout__1_carry_i_12_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF4F44)) 
    tout__1_carry_i_13
       (.I0(tout__1_carry_i_15_n_0),
        .I1(tout__1_carry_i_16_n_0),
        .I2(tout__1_carry_i_17_n_0),
        .I3(tout__1_carry_i_18_n_0),
        .I4(ir1[11]),
        .I5(tout__1_carry_i_19_n_0),
        .O(tout__1_carry_i_13_n_0));
  MUXF7 tout__1_carry_i_14
       (.I0(tout__1_carry_i_21_n_0),
        .I1(tout__1_carry_i_22_n_0),
        .O(tout__1_carry_i_14_n_0),
        .S(tout__1_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    tout__1_carry_i_15
       (.I0(ir1[7]),
        .I1(ir1[8]),
        .I2(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I3(\stat[2]_i_10__0_n_0 ),
        .I4(ir1[6]),
        .I5(ir1[2]),
        .O(tout__1_carry_i_15_n_0));
  LUT6 #(
    .INIT(64'h00003F003F007700)) 
    tout__1_carry_i_16
       (.I0(\rgf_selc1_wb_reg[1] [0]),
        .I1(\rgf_selc1_wb_reg[1] [1]),
        .I2(ir1[0]),
        .I3(ctl_fetch1_fl_i_20_n_0),
        .I4(ir1[3]),
        .I5(ir1[1]),
        .O(tout__1_carry_i_16_n_0));
  LUT6 #(
    .INIT(64'h99989888FFFFFFFF)) 
    tout__1_carry_i_17
       (.I0(\rgf_selc1_wb_reg[1] [1]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(ir1[8]),
        .I3(ir1[10]),
        .I4(ir1[9]),
        .I5(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .O(tout__1_carry_i_17_n_0));
  LUT6 #(
    .INIT(64'hAAAEAAAFAAAAAAAA)) 
    tout__1_carry_i_18
       (.I0(rst_n_fl_reg_9),
        .I1(ir1[7]),
        .I2(ir1[8]),
        .I3(ir1[9]),
        .I4(\rgf_selc1_wb_reg[1] [1]),
        .I5(ir1[10]),
        .O(tout__1_carry_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFEEFEEEEEEEEE)) 
    tout__1_carry_i_19
       (.I0(\rgf_selc1_wb_reg[1] [2]),
        .I1(ir1[15]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(tout__1_carry_i_23_n_0),
        .I4(tout__1_carry_i_24_n_0),
        .I5(ir1[11]),
        .O(tout__1_carry_i_19_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_1__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[10]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[2]),
        .O(DI[2]));
  LUT4 #(
    .INIT(16'h1E00)) 
    tout__1_carry_i_2
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[1]),
        .O(\badr[2]_INST_0_i_2 [1]));
  LUT6 #(
    .INIT(64'hFF00FF00EF00FF00)) 
    tout__1_carry_i_20
       (.I0(ir1[12]),
        .I1(ir1[14]),
        .I2(\sr_reg[15]_0 [6]),
        .I3(ir1[13]),
        .I4(\rgf_c1bus_wb[14]_i_53_0 ),
        .I5(ir1[15]),
        .O(tout__1_carry_i_20_n_0));
  LUT6 #(
    .INIT(64'h14FF14FFFFFF0000)) 
    tout__1_carry_i_21
       (.I0(ir1[15]),
        .I1(\badr[15]_INST_0_i_25_0 ),
        .I2(ir1[11]),
        .I3(\rgf_c1bus_wb[14]_i_53_0 ),
        .I4(tout__1_carry_i_25_n_0),
        .I5(ir1[12]),
        .O(tout__1_carry_i_21_n_0));
  LUT6 #(
    .INIT(64'hBFFFBFBFAAAAAAAA)) 
    tout__1_carry_i_22
       (.I0(ir1[15]),
        .I1(ir1[12]),
        .I2(ir1[14]),
        .I3(tout__1_carry_i_26_n_0),
        .I4(tout__1_carry_i_27_n_0),
        .I5(tout__1_carry_i_28_n_0),
        .O(tout__1_carry_i_22_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    tout__1_carry_i_23
       (.I0(ir1[7]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .O(tout__1_carry_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF7FFFFFFF)) 
    tout__1_carry_i_24
       (.I0(ir1[8]),
        .I1(ir1[14]),
        .I2(ir1[13]),
        .I3(ir1[12]),
        .I4(ir1[10]),
        .I5(ir1[9]),
        .O(tout__1_carry_i_24_n_0));
  LUT6 #(
    .INIT(64'h00000000F55F75DF)) 
    tout__1_carry_i_25
       (.I0(\rgf_c1bus_wb[14]_i_53_0 ),
        .I1(\sr_reg[15]_0 [5]),
        .I2(ir1[14]),
        .I3(ir1[11]),
        .I4(ir1[15]),
        .I5(tout__1_carry_i_29_n_0),
        .O(tout__1_carry_i_25_n_0));
  LUT6 #(
    .INIT(64'hAAAAFFEFAAAAFAEA)) 
    tout__1_carry_i_26
       (.I0(\rgf_selc1_wb[0]_i_21_n_0 ),
        .I1(ir1[7]),
        .I2(ir1[11]),
        .I3(\stat[1]_i_18_n_0 ),
        .I4(tout__1_carry_i_30_n_0),
        .I5(tout__1_carry_i_31_n_0),
        .O(tout__1_carry_i_26_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBAAAAABAA)) 
    tout__1_carry_i_27
       (.I0(tout__1_carry_i_22_0),
        .I1(tout__1_carry_i_32_n_0),
        .I2(\rgf_selc1_rn_wb[1]_i_9_n_0 ),
        .I3(\rgf_selc1_wb_reg[1] [0]),
        .I4(ir1[8]),
        .I5(tout__1_carry_i_33_n_0),
        .O(tout__1_carry_i_27_n_0));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFEFC)) 
    tout__1_carry_i_28
       (.I0(ir1[12]),
        .I1(\rgf_selc1_wb_reg[1] [0]),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(\sr_reg[15]_0 [7]),
        .I4(ir1[14]),
        .I5(ir1[11]),
        .O(tout__1_carry_i_28_n_0));
  LUT6 #(
    .INIT(64'h0001001101411101)) 
    tout__1_carry_i_29
       (.I0(tout__1_carry_i_34_n_0),
        .I1(tout__1_carry_i_25_0),
        .I2(\rgf_selc1_wb_reg[1] [1]),
        .I3(ir1[3]),
        .I4(ir1[0]),
        .I5(ir1[1]),
        .O(tout__1_carry_i_29_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_2__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[9]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[1]),
        .O(DI[1]));
  LUT6 #(
    .INIT(64'hFFFF8B338B330000)) 
    tout__1_carry_i_3
       (.I0(\stat_reg[1]_0 ),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\stat_reg[2]_4 ),
        .I3(tout__1_carry_i_11_n_0),
        .I4(tout__1_carry_i_12_n_0),
        .I5(a1bus_0[0]),
        .O(DI[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD8)) 
    tout__1_carry_i_30
       (.I0(ir1[11]),
        .I1(ir1[9]),
        .I2(ir1[6]),
        .I3(\rgf_selc1_wb_reg[1] [1]),
        .I4(ir1[10]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(tout__1_carry_i_30_n_0));
  LUT3 #(
    .INIT(8'h2A)) 
    tout__1_carry_i_31
       (.I0(rst_n_fl_reg_9),
        .I1(ir1[9]),
        .I2(ir1[8]),
        .O(tout__1_carry_i_31_n_0));
  LUT5 #(
    .INIT(32'h80000000)) 
    tout__1_carry_i_32
       (.I0(tout__1_carry_i_36_n_0),
        .I1(ir1[9]),
        .I2(ir1[11]),
        .I3(ir1[8]),
        .I4(tout__1_carry_i_37_n_0),
        .O(tout__1_carry_i_32_n_0));
  LUT6 #(
    .INIT(64'hFFFF06FFFFFF0406)) 
    tout__1_carry_i_33
       (.I0(ir1[7]),
        .I1(ir1[6]),
        .I2(\rgf_selc1_wb_reg[1] [0]),
        .I3(ir1[11]),
        .I4(ir1[9]),
        .I5(ir1[8]),
        .O(tout__1_carry_i_33_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    tout__1_carry_i_34
       (.I0(ctl_fetch1_fl_i_36_n_0),
        .I1(ir1[14]),
        .I2(ir1[15]),
        .I3(ir1[11]),
        .I4(ir1[6]),
        .O(tout__1_carry_i_34_n_0));
  LUT6 #(
    .INIT(64'h5555F7F55D55F5F5)) 
    tout__1_carry_i_36
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[7]),
        .I4(ir1[6]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(tout__1_carry_i_36_n_0));
  LUT6 #(
    .INIT(64'hAA0AAA0AAA3BEA0A)) 
    tout__1_carry_i_37
       (.I0(ir1[3]),
        .I1(ir1[4]),
        .I2(ir1[5]),
        .I3(ir1[6]),
        .I4(ir1[7]),
        .I5(\rgf_selc1_wb_reg[1] [0]),
        .O(tout__1_carry_i_37_n_0));
  LUT5 #(
    .INIT(32'h1EFF001E)) 
    tout__1_carry_i_3__0
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\tr_reg[0]_0 ),
        .I3(tout__1_carry_i_9_n_0),
        .I4(a0bus_0[0]),
        .O(\badr[2]_INST_0_i_2 [0]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry_i_4
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[3]),
        .I4(\badr[2]_INST_0_i_2 [2]),
        .O(tout__1_carry_i_1_0[3]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_4__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[3]),
        .I3(DI[2]),
        .O(tout__1_carry_i_1__0_0[3]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry_i_5
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[2]),
        .I4(\badr[2]_INST_0_i_2 [1]),
        .O(tout__1_carry_i_1_0[2]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_5__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[10]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[2]),
        .I3(DI[1]),
        .O(tout__1_carry_i_1__0_0[2]));
  LUT5 #(
    .INIT(32'h1EE1E11E)) 
    tout__1_carry_i_6
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[1]),
        .I4(\badr[2]_INST_0_i_2 [0]),
        .O(tout__1_carry_i_1_0[1]));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_6__0
       (.I0(\stat_reg[2]_3 ),
        .I1(\bdatw[9]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[1]),
        .I3(DI[0]),
        .O(tout__1_carry_i_1__0_0[1]));
  LUT6 #(
    .INIT(64'h8B3374CC74CC8B33)) 
    tout__1_carry_i_7
       (.I0(\stat_reg[1]_0 ),
        .I1(\sr_reg[15]_0 [6]),
        .I2(\stat_reg[2]_4 ),
        .I3(tout__1_carry_i_11_n_0),
        .I4(a1bus_0[0]),
        .I5(tout__1_carry_i_12_n_0),
        .O(tout__1_carry_i_1__0_0[0]));
  LUT5 #(
    .INIT(32'hE11E1EE1)) 
    tout__1_carry_i_7__0
       (.I0(\stat_reg[2]_10 ),
        .I1(\rgf_c0bus_wb[15]_i_8_0 ),
        .I2(\tr_reg[0]_0 ),
        .I3(tout__1_carry_i_9_n_0),
        .I4(a0bus_0[0]),
        .O(tout__1_carry_i_1_0[0]));
  LUT6 #(
    .INIT(64'hFD00FDFDFDFDFDFD)) 
    tout__1_carry_i_8
       (.I0(\stat_reg[1]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I3(\stat_reg[2]_10 ),
        .I4(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_8_0 ));
  LUT6 #(
    .INIT(64'h00000000000E0001)) 
    tout__1_carry_i_8__0
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\stat_reg[2]_4 ),
        .O(\stat_reg[2]_3 ));
  LUT6 #(
    .INIT(64'hF0F0F0F0BFB0B0B0)) 
    tout__1_carry_i_9
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\stat_reg[1]_1 ),
        .I2(\sr_reg[15]_0 [6]),
        .I3(\stat_reg[2]_10 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\stat_reg[0]_2 ),
        .O(tout__1_carry_i_9_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    tout__1_carry_i_9__0
       (.I0(tout__1_carry_i_13_n_0),
        .I1(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .O(\stat_reg[1]_0 ));
endmodule

module mcss_fch_fsm
   (fch_wrbufn1,
    p_2_in,
    rst_n_fl_reg,
    \sr_reg[15] ,
    rst_n_0,
    rgf_selc1_stat_reg,
    D,
    \stat_reg[1]_0 ,
    \sp_reg[15] ,
    fch_issu1_ir,
    \stat_reg[2]_0 ,
    E,
    brdy_0,
    fadr,
    \stat_reg[0]_0 ,
    \stat_reg[1]_1 ,
    S,
    rst_n_fl_reg_0,
    ctl_fetch0,
    crdy_0,
    ctl_fetch1,
    \stat_reg[0]_1 ,
    \stat_reg[1]_2 ,
    rst_n_fl_reg_1,
    rst_n_fl_reg_2,
    rst_n_fl_reg_3,
    fch_memacc1,
    in0,
    ir1,
    fch_issu1,
    rst_n_fl_reg_4,
    eir,
    \pc_reg[7] ,
    \pc_reg[11] ,
    \pc_reg[12] ,
    fch_irq_req_fl_reg,
    \sr_reg[1] ,
    \sr_reg[0] ,
    \sr_reg[0]_0 ,
    \sr_reg[0]_1 ,
    \sr_reg[1]_0 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[1]_1 ,
    \sr_reg[0]_5 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[1]_2 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[1]_3 ,
    \sr_reg[0]_11 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[1]_4 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[0]_17 ,
    \sr_reg[1]_5 ,
    \sr_reg[0]_18 ,
    \sr_reg[0]_19 ,
    \iv_reg[15] ,
    \tr_reg[15] ,
    rgf_selc1_stat_reg_0,
    rgf_selc1_stat_reg_1,
    rgf_selc1_stat_reg_2,
    rgf_selc1_stat_reg_3,
    rgf_selc1_stat_reg_4,
    rgf_selc1_stat_reg_5,
    rgf_selc1_stat_reg_6,
    rgf_selc1_stat_reg_7,
    rgf_selc1_stat_reg_8,
    rgf_selc1_stat_reg_9,
    rgf_selc1_stat_reg_10,
    rgf_selc1_stat_reg_11,
    rgf_selc1_stat_reg_12,
    rgf_selc1_stat_reg_13,
    rgf_selc1_stat_reg_14,
    rgf_selc1_stat_reg_15,
    rgf_selc1_stat_reg_16,
    rgf_selc1_stat_reg_17,
    rgf_selc1_stat_reg_18,
    rgf_selc1_stat_reg_19,
    rgf_selc1_stat_reg_20,
    rgf_selc1_stat_reg_21,
    rgf_selc1_stat_reg_22,
    rgf_selc1_stat_reg_23,
    rgf_selc1_stat_reg_24,
    rgf_selc1_stat_reg_25,
    rgf_selc1_stat_reg_26,
    rgf_selc1_stat_reg_27,
    rgf_selc1_stat_reg_28,
    rgf_selc1_stat_reg_29,
    rgf_selc1_stat_reg_30,
    rgf_selc1_stat_reg_31,
    \sr_reg[0]_20 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[1]_6 ,
    clk,
    \grn_reg[15] ,
    \pc_reg[15] ,
    rgf_selc1_stat,
    Q,
    \pc_reg[15]_0 ,
    rgf_selc0_stat,
    \pc_reg[15]_1 ,
    \pc_reg[14] ,
    \pc_reg[14]_0 ,
    \sr_reg[3] ,
    \sr_reg[3]_0 ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \grn[15]_i_3__5_0 ,
    \grn[15]_i_3__5_1 ,
    \sr[13]_i_5_0 ,
    \sr[13]_i_5_1 ,
    \sr[13]_i_5_2 ,
    \sr[13]_i_5_3 ,
    alu_sr_flag1,
    \sr_reg[4] ,
    alu_sr_flag0,
    \sr_reg[5] ,
    \sr_reg[5]_0 ,
    \sr_reg[5]_1 ,
    \sr_reg[5]_2 ,
    \sr_reg[5]_3 ,
    \sr_reg[5]_4 ,
    \sr_reg[15]_0 ,
    \sr_reg[6] ,
    \sr_reg[6]_0 ,
    \sr_reg[7] ,
    \sr_reg[5]_5 ,
    \sr_reg[5]_6 ,
    \sr_reg[5]_7 ,
    \sr_reg[5]_8 ,
    \sr_reg[5]_9 ,
    \sr_reg[6]_1 ,
    ctl_sr_ldie1,
    ctl_sr_upd0,
    fch_irq_lev,
    rst_n,
    ctl_sr_upd1,
    \pc_reg[15]_2 ,
    \pc_reg[14]_1 ,
    \pc_reg[13] ,
    \pc_reg[0] ,
    \pc0_reg[12] ,
    \pc0_reg[3] ,
    fch_irq_req,
    p_2_in_0,
    \sp_reg[15]_0 ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[1] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[0] ,
    \sp_reg[2] ,
    O,
    \fadr[8] ,
    \fadr[12] ,
    fch_leir_nir_reg_0,
    ctl_fetch1_fl_i_21_0,
    fch_leir_nir_reg_1,
    \stat_reg[0]_2 ,
    \stat[2]_i_4_0 ,
    ctl_fetch0_fl_reg,
    ctl_fetch0_fl_reg_0,
    \stat[2]_i_4_1 ,
    \stat[2]_i_4_2 ,
    ctl_fetch0_fl_reg_1,
    ctl_fetch0_fl_reg_2,
    ctl_fetch0_fl_reg_3,
    ctl_fetch0_fl_reg_4,
    ctl_fetch0_fl_i_15_0,
    \sr[13]_i_13 ,
    crdy,
    brdy,
    \stat_reg[0]_3 ,
    ctl_fetch1_fl_reg,
    ctl_fetch1_fl_reg_i_6_0,
    ctl_fetch1_fl_reg_i_6_1,
    ctl_fetch1_fl_reg_i_6_2,
    ctl_fetch1_fl_i_2_0,
    ctl_fetch1_fl_i_16_0,
    \stat_reg[0]_4 ,
    \stat_reg[0]_5 ,
    \stat_reg[0]_6 ,
    \stat_reg[0]_7 ,
    ctl_fetch0_fl_reg_5,
    ctl_fetch0_fl_i_2_0,
    ctl_fetch0_fl_i_8_0,
    ctl_fetch0_fl_i_4_0,
    ctl_fetch0_fl_i_4_1,
    ctl_fetch0_fl_i_16_0,
    ctl_fetch0_fl_i_16_1,
    ctl_fetch1_fl_i_25_0,
    ctl_fetch1_fl_i_25_1,
    ctl_fetch1_fl_i_27_0,
    ctl_fetch1_fl_i_27_1,
    ctl_fetch1_fl_i_2_1,
    ctl_fetch1_fl_i_2_2,
    ctl_fetch1_fl_i_2_3,
    ctl_fetch1_fl_reg_0,
    ctl_fetch1_fl_reg_1,
    ctl_fetch1_fl_i_2_4,
    ctl_fetch1_fl_i_27_2,
    \fch_irq_lev[1]_i_2 ,
    \fch_irq_lev[1]_i_2_0 ,
    ctl_fetch1_fl_i_34_0,
    ctl_fetch1_fl_i_2_5,
    \ir0_fl_reg[0] ,
    \stat_reg[0]_8 ,
    rst_n_fl,
    \ir1_id_fl_reg[21] ,
    fch_term_fl,
    out,
    ctl_fetch0_fl,
    \ir0_fl_reg[15] ,
    \ir0_id_fl_reg[21] ,
    \ir1_id_fl_reg[20] ,
    \ir0_id_fl_reg[20] ,
    fch_issu1_inferred_i_11_0,
    \ir1_id_fl_reg[21]_0 ,
    fadr_1_fl,
    \ir1_id_fl_reg[21]_1 ,
    \ir1_fl_reg[0] ,
    ctl_fetch1_fl,
    \ir1_fl_reg[15] ,
    fdat,
    fdatx,
    fch_issu1_inferred_i_8_0,
    fch_issu1_inferred_i_8_1,
    fch_issu1_inferred_i_8_2,
    fch_issu1_inferred_i_20_0,
    fch_issu1_inferred_i_20_1,
    fch_issu1_inferred_i_20_2,
    fch_issu1_inferred_i_2_0,
    fch_issu1_inferred_i_8_3,
    fch_issu1_inferred_i_8_4,
    fch_issu1_inferred_i_8_5,
    fch_issu1_inferred_i_7_0,
    fch_issu1_inferred_i_6_0,
    fch_issu1_inferred_i_8_6,
    fch_issu1_inferred_i_8_7,
    fch_issu1_inferred_i_8_8,
    fch_issu1_inferred_i_8_9,
    fch_issu1_inferred_i_8_10,
    fch_issu1_inferred_i_33_0,
    fch_issu1_inferred_i_33_1,
    fch_issu1_inferred_i_33_2,
    fch_issu1_inferred_i_33_3,
    fch_issu1_inferred_i_7_1,
    fch_issu1_inferred_i_7_2,
    fch_issu1_inferred_i_7_3,
    fch_issu1_inferred_i_7_4,
    fch_issu1_inferred_i_41_0,
    fch_issu1_inferred_i_41_1,
    fch_issu1_inferred_i_7_5,
    fch_issu1_inferred_i_6_1,
    fch_issu1_inferred_i_7_6,
    fch_issu1_inferred_i_2_1,
    fch_issu1_inferred_i_2_2,
    fch_issu1_inferred_i_1_0,
    fch_issu1_inferred_i_1_1,
    fch_issu1_inferred_i_1_2,
    fch_issu1_inferred_i_6_2,
    fch_issu1_inferred_i_6_3,
    fch_issu1_inferred_i_6_4,
    fch_issu1_inferred_i_41_2,
    fch_issu1_inferred_i_41_3,
    fch_issu1_inferred_i_11_1,
    fch_issu1_inferred_i_11_2,
    fch_issu1_inferred_i_1_3,
    fch_issu1_inferred_i_1_4,
    fch_issu1_inferred_i_5_0,
    fch_issu1_inferred_i_5_1,
    fch_issu1_inferred_i_1_5,
    fch_issu1_inferred_i_1_6,
    fch_issu1_inferred_i_11_3,
    fch_issu1_inferred_i_11_4,
    fch_issu1_inferred_i_11_5,
    fch_issu1_inferred_i_28_0,
    fch_issu1_inferred_i_28_1,
    fch_issu1_inferred_i_28_2,
    fch_issu1_inferred_i_28_3,
    \eir_fl_reg[15] ,
    fch_issu1_inferred_i_32_0,
    fch_issu1_inferred_i_32_1,
    fch_issu1_inferred_i_32_2,
    fch_issu1_inferred_i_31_0,
    ctl_fetch0_fl_i_27_0,
    fch_issu1_fl,
    ctl_fetch_ext_fl,
    \eir_fl_reg[15]_0 ,
    fch_leir_lir_reg_0,
    fch_leir_lir_reg_1,
    ctl_fetch1_fl_i_2_6,
    ctl_sr_ldie0,
    cpuid,
    \sr_reg[7]_0 ,
    \sr_reg[7]_1 ,
    \iv_reg[15]_0 ,
    \tr_reg[15]_0 );
  output fch_wrbufn1;
  output p_2_in;
  output rst_n_fl_reg;
  output [15:0]\sr_reg[15] ;
  output rst_n_0;
  output [15:0]rgf_selc1_stat_reg;
  output [12:0]D;
  output \stat_reg[1]_0 ;
  output [15:0]\sp_reg[15] ;
  output fch_issu1_ir;
  output \stat_reg[2]_0 ;
  output [0:0]E;
  output [0:0]brdy_0;
  output [12:0]fadr;
  output \stat_reg[0]_0 ;
  output \stat_reg[1]_1 ;
  output [3:0]S;
  output rst_n_fl_reg_0;
  output ctl_fetch0;
  output crdy_0;
  output ctl_fetch1;
  output [0:0]\stat_reg[0]_1 ;
  output \stat_reg[1]_2 ;
  output rst_n_fl_reg_1;
  output rst_n_fl_reg_2;
  output [1:0]rst_n_fl_reg_3;
  output fch_memacc1;
  output [15:0]in0;
  output [15:0]ir1;
  output fch_issu1;
  output rst_n_fl_reg_4;
  output [15:0]eir;
  output [3:0]\pc_reg[7] ;
  output [3:0]\pc_reg[11] ;
  output [0:0]\pc_reg[12] ;
  output fch_irq_req_fl_reg;
  output [0:0]\sr_reg[1] ;
  output [0:0]\sr_reg[0] ;
  output [0:0]\sr_reg[0]_0 ;
  output [0:0]\sr_reg[0]_1 ;
  output [0:0]\sr_reg[1]_0 ;
  output [0:0]\sr_reg[0]_2 ;
  output [0:0]\sr_reg[0]_3 ;
  output [0:0]\sr_reg[0]_4 ;
  output [0:0]\sr_reg[1]_1 ;
  output [0:0]\sr_reg[0]_5 ;
  output [0:0]\sr_reg[0]_6 ;
  output [0:0]\sr_reg[0]_7 ;
  output [0:0]\sr_reg[1]_2 ;
  output [0:0]\sr_reg[0]_8 ;
  output [0:0]\sr_reg[0]_9 ;
  output [0:0]\sr_reg[0]_10 ;
  output [0:0]\sr_reg[1]_3 ;
  output [0:0]\sr_reg[0]_11 ;
  output [0:0]\sr_reg[0]_12 ;
  output [0:0]\sr_reg[0]_13 ;
  output [0:0]\sr_reg[1]_4 ;
  output [0:0]\sr_reg[0]_14 ;
  output [0:0]\sr_reg[0]_15 ;
  output [0:0]\sr_reg[0]_16 ;
  output [0:0]\sr_reg[0]_17 ;
  output [0:0]\sr_reg[1]_5 ;
  output [0:0]\sr_reg[0]_18 ;
  output [0:0]\sr_reg[0]_19 ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15] ;
  output [15:0]rgf_selc1_stat_reg_0;
  output [15:0]rgf_selc1_stat_reg_1;
  output [15:0]rgf_selc1_stat_reg_2;
  output [15:0]rgf_selc1_stat_reg_3;
  output [15:0]rgf_selc1_stat_reg_4;
  output [15:0]rgf_selc1_stat_reg_5;
  output [15:0]rgf_selc1_stat_reg_6;
  output [15:0]rgf_selc1_stat_reg_7;
  output [15:0]rgf_selc1_stat_reg_8;
  output [15:0]rgf_selc1_stat_reg_9;
  output [15:0]rgf_selc1_stat_reg_10;
  output [15:0]rgf_selc1_stat_reg_11;
  output [15:0]rgf_selc1_stat_reg_12;
  output [15:0]rgf_selc1_stat_reg_13;
  output [15:0]rgf_selc1_stat_reg_14;
  output [15:0]rgf_selc1_stat_reg_15;
  output [15:0]rgf_selc1_stat_reg_16;
  output [15:0]rgf_selc1_stat_reg_17;
  output [15:0]rgf_selc1_stat_reg_18;
  output [15:0]rgf_selc1_stat_reg_19;
  output [15:0]rgf_selc1_stat_reg_20;
  output [15:0]rgf_selc1_stat_reg_21;
  output [15:0]rgf_selc1_stat_reg_22;
  output [15:0]rgf_selc1_stat_reg_23;
  output [15:0]rgf_selc1_stat_reg_24;
  output [15:0]rgf_selc1_stat_reg_25;
  output [15:0]rgf_selc1_stat_reg_26;
  output [15:0]rgf_selc1_stat_reg_27;
  output [15:0]rgf_selc1_stat_reg_28;
  output [15:0]rgf_selc1_stat_reg_29;
  output [15:0]rgf_selc1_stat_reg_30;
  output [15:0]rgf_selc1_stat_reg_31;
  output [0:0]\sr_reg[0]_20 ;
  output [0:0]\sr_reg[0]_21 ;
  output [0:0]\sr_reg[0]_22 ;
  output [0:0]\sr_reg[1]_6 ;
  input clk;
  input \grn_reg[15] ;
  input [15:0]\pc_reg[15] ;
  input rgf_selc1_stat;
  input [15:0]Q;
  input [13:0]\pc_reg[15]_0 ;
  input rgf_selc0_stat;
  input [15:0]\pc_reg[15]_1 ;
  input \pc_reg[14] ;
  input \pc_reg[14]_0 ;
  input \sr_reg[3] ;
  input \sr_reg[3]_0 ;
  input [2:0]\grn_reg[15]_0 ;
  input [2:0]\grn_reg[15]_1 ;
  input [1:0]\grn[15]_i_3__5_0 ;
  input [1:0]\grn[15]_i_3__5_1 ;
  input [2:0]\sr[13]_i_5_0 ;
  input [2:0]\sr[13]_i_5_1 ;
  input [1:0]\sr[13]_i_5_2 ;
  input [1:0]\sr[13]_i_5_3 ;
  input [0:0]alu_sr_flag1;
  input \sr_reg[4] ;
  input [1:0]alu_sr_flag0;
  input \sr_reg[5] ;
  input \sr_reg[5]_0 ;
  input \sr_reg[5]_1 ;
  input \sr_reg[5]_2 ;
  input \sr_reg[5]_3 ;
  input \sr_reg[5]_4 ;
  input [15:0]\sr_reg[15]_0 ;
  input \sr_reg[6] ;
  input [0:0]\sr_reg[6]_0 ;
  input \sr_reg[7] ;
  input \sr_reg[5]_5 ;
  input \sr_reg[5]_6 ;
  input \sr_reg[5]_7 ;
  input \sr_reg[5]_8 ;
  input \sr_reg[5]_9 ;
  input \sr_reg[6]_1 ;
  input ctl_sr_ldie1;
  input ctl_sr_upd0;
  input [1:0]fch_irq_lev;
  input rst_n;
  input ctl_sr_upd1;
  input \pc_reg[15]_2 ;
  input \pc_reg[14]_1 ;
  input \pc_reg[13] ;
  input \pc_reg[0] ;
  input [12:0]\pc0_reg[12] ;
  input \pc0_reg[3] ;
  input fch_irq_req;
  input [12:0]p_2_in_0;
  input \sp_reg[15]_0 ;
  input \sp_reg[14] ;
  input \sp_reg[13] ;
  input \sp_reg[12] ;
  input \sp_reg[11] ;
  input \sp_reg[10] ;
  input \sp_reg[9] ;
  input \sp_reg[8] ;
  input \sp_reg[7] ;
  input \sp_reg[6] ;
  input \sp_reg[5] ;
  input \sp_reg[1] ;
  input \sp_reg[3] ;
  input \sp_reg[4] ;
  input \sp_reg[0] ;
  input \sp_reg[2] ;
  input [3:0]O;
  input [3:0]\fadr[8] ;
  input [3:0]\fadr[12] ;
  input fch_leir_nir_reg_0;
  input [15:0]ctl_fetch1_fl_i_21_0;
  input fch_leir_nir_reg_1;
  input \stat_reg[0]_2 ;
  input \stat[2]_i_4_0 ;
  input [15:0]ctl_fetch0_fl_reg;
  input [2:0]ctl_fetch0_fl_reg_0;
  input \stat[2]_i_4_1 ;
  input \stat[2]_i_4_2 ;
  input ctl_fetch0_fl_reg_1;
  input ctl_fetch0_fl_reg_2;
  input ctl_fetch0_fl_reg_3;
  input ctl_fetch0_fl_reg_4;
  input ctl_fetch0_fl_i_15_0;
  input \sr[13]_i_13 ;
  input crdy;
  input brdy;
  input \stat_reg[0]_3 ;
  input [2:0]ctl_fetch1_fl_reg;
  input ctl_fetch1_fl_reg_i_6_0;
  input ctl_fetch1_fl_reg_i_6_1;
  input ctl_fetch1_fl_reg_i_6_2;
  input ctl_fetch1_fl_i_2_0;
  input ctl_fetch1_fl_i_16_0;
  input \stat_reg[0]_4 ;
  input \stat_reg[0]_5 ;
  input \stat_reg[0]_6 ;
  input \stat_reg[0]_7 ;
  input ctl_fetch0_fl_reg_5;
  input ctl_fetch0_fl_i_2_0;
  input ctl_fetch0_fl_i_8_0;
  input ctl_fetch0_fl_i_4_0;
  input ctl_fetch0_fl_i_4_1;
  input ctl_fetch0_fl_i_16_0;
  input ctl_fetch0_fl_i_16_1;
  input ctl_fetch1_fl_i_25_0;
  input ctl_fetch1_fl_i_25_1;
  input ctl_fetch1_fl_i_27_0;
  input ctl_fetch1_fl_i_27_1;
  input ctl_fetch1_fl_i_2_1;
  input ctl_fetch1_fl_i_2_2;
  input ctl_fetch1_fl_i_2_3;
  input ctl_fetch1_fl_reg_0;
  input ctl_fetch1_fl_reg_1;
  input ctl_fetch1_fl_i_2_4;
  input ctl_fetch1_fl_i_27_2;
  input \fch_irq_lev[1]_i_2 ;
  input \fch_irq_lev[1]_i_2_0 ;
  input ctl_fetch1_fl_i_34_0;
  input ctl_fetch1_fl_i_2_5;
  input \ir0_fl_reg[0] ;
  input [1:0]\stat_reg[0]_8 ;
  input rst_n_fl;
  input [1:0]\ir1_id_fl_reg[21] ;
  input fch_term_fl;
  input out;
  input ctl_fetch0_fl;
  input [15:0]\ir0_fl_reg[15] ;
  input [1:0]\ir0_id_fl_reg[21] ;
  input \ir1_id_fl_reg[20] ;
  input \ir0_id_fl_reg[20] ;
  input [10:0]fch_issu1_inferred_i_11_0;
  input [5:0]\ir1_id_fl_reg[21]_0 ;
  input fadr_1_fl;
  input \ir1_id_fl_reg[21]_1 ;
  input \ir1_fl_reg[0] ;
  input ctl_fetch1_fl;
  input [15:0]\ir1_fl_reg[15] ;
  input [15:0]fdat;
  input [15:0]fdatx;
  input fch_issu1_inferred_i_8_0;
  input fch_issu1_inferred_i_8_1;
  input fch_issu1_inferred_i_8_2;
  input fch_issu1_inferred_i_20_0;
  input fch_issu1_inferred_i_20_1;
  input fch_issu1_inferred_i_20_2;
  input fch_issu1_inferred_i_2_0;
  input fch_issu1_inferred_i_8_3;
  input fch_issu1_inferred_i_8_4;
  input fch_issu1_inferred_i_8_5;
  input fch_issu1_inferred_i_7_0;
  input fch_issu1_inferred_i_6_0;
  input fch_issu1_inferred_i_8_6;
  input fch_issu1_inferred_i_8_7;
  input fch_issu1_inferred_i_8_8;
  input fch_issu1_inferred_i_8_9;
  input fch_issu1_inferred_i_8_10;
  input fch_issu1_inferred_i_33_0;
  input fch_issu1_inferred_i_33_1;
  input fch_issu1_inferred_i_33_2;
  input fch_issu1_inferred_i_33_3;
  input fch_issu1_inferred_i_7_1;
  input fch_issu1_inferred_i_7_2;
  input fch_issu1_inferred_i_7_3;
  input fch_issu1_inferred_i_7_4;
  input fch_issu1_inferred_i_41_0;
  input fch_issu1_inferred_i_41_1;
  input fch_issu1_inferred_i_7_5;
  input fch_issu1_inferred_i_6_1;
  input fch_issu1_inferred_i_7_6;
  input fch_issu1_inferred_i_2_1;
  input fch_issu1_inferred_i_2_2;
  input fch_issu1_inferred_i_1_0;
  input fch_issu1_inferred_i_1_1;
  input fch_issu1_inferred_i_1_2;
  input fch_issu1_inferred_i_6_2;
  input fch_issu1_inferred_i_6_3;
  input fch_issu1_inferred_i_6_4;
  input fch_issu1_inferred_i_41_2;
  input fch_issu1_inferred_i_41_3;
  input fch_issu1_inferred_i_11_1;
  input fch_issu1_inferred_i_11_2;
  input fch_issu1_inferred_i_1_3;
  input fch_issu1_inferred_i_1_4;
  input fch_issu1_inferred_i_5_0;
  input fch_issu1_inferred_i_5_1;
  input fch_issu1_inferred_i_1_5;
  input fch_issu1_inferred_i_1_6;
  input fch_issu1_inferred_i_11_3;
  input fch_issu1_inferred_i_11_4;
  input fch_issu1_inferred_i_11_5;
  input fch_issu1_inferred_i_28_0;
  input fch_issu1_inferred_i_28_1;
  input fch_issu1_inferred_i_28_2;
  input fch_issu1_inferred_i_28_3;
  input [15:0]\eir_fl_reg[15] ;
  input fch_issu1_inferred_i_32_0;
  input fch_issu1_inferred_i_32_1;
  input fch_issu1_inferred_i_32_2;
  input fch_issu1_inferred_i_31_0;
  input ctl_fetch0_fl_i_27_0;
  input fch_issu1_fl;
  input ctl_fetch_ext_fl;
  input [15:0]\eir_fl_reg[15]_0 ;
  input fch_leir_lir_reg_0;
  input fch_leir_lir_reg_1;
  input ctl_fetch1_fl_i_2_6;
  input ctl_sr_ldie0;
  input [1:0]cpuid;
  input \sr_reg[7]_0 ;
  input [0:0]\sr_reg[7]_1 ;
  input [15:0]\iv_reg[15]_0 ;
  input [15:0]\tr_reg[15]_0 ;

  wire \<const1> ;
  wire [12:0]D;
  wire [0:0]E;
  wire [3:0]O;
  wire [15:0]Q;
  wire [3:0]S;
  wire [1:0]alu_sr_flag0;
  wire [0:0]alu_sr_flag1;
  wire brdy;
  wire [0:0]brdy_0;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire crdy_0;
  wire ctl_fetch0;
  wire ctl_fetch0_fl;
  wire ctl_fetch0_fl_i_11_n_0;
  wire ctl_fetch0_fl_i_12_n_0;
  wire ctl_fetch0_fl_i_13_n_0;
  wire ctl_fetch0_fl_i_14_n_0;
  wire ctl_fetch0_fl_i_15_0;
  wire ctl_fetch0_fl_i_15_n_0;
  wire ctl_fetch0_fl_i_16_0;
  wire ctl_fetch0_fl_i_16_1;
  wire ctl_fetch0_fl_i_16_n_0;
  wire ctl_fetch0_fl_i_17_n_0;
  wire ctl_fetch0_fl_i_19_n_0;
  wire ctl_fetch0_fl_i_20_n_0;
  wire ctl_fetch0_fl_i_21_n_0;
  wire ctl_fetch0_fl_i_22_n_0;
  wire ctl_fetch0_fl_i_23_n_0;
  wire ctl_fetch0_fl_i_24_n_0;
  wire ctl_fetch0_fl_i_25_n_0;
  wire ctl_fetch0_fl_i_26_n_0;
  wire ctl_fetch0_fl_i_27_0;
  wire ctl_fetch0_fl_i_27_n_0;
  wire ctl_fetch0_fl_i_28_n_0;
  wire ctl_fetch0_fl_i_29_n_0;
  wire ctl_fetch0_fl_i_2_0;
  wire ctl_fetch0_fl_i_2_n_0;
  wire ctl_fetch0_fl_i_30_n_0;
  wire ctl_fetch0_fl_i_31_n_0;
  wire ctl_fetch0_fl_i_32_n_0;
  wire ctl_fetch0_fl_i_33_n_0;
  wire ctl_fetch0_fl_i_34_n_0;
  wire ctl_fetch0_fl_i_36_n_0;
  wire ctl_fetch0_fl_i_37_n_0;
  wire ctl_fetch0_fl_i_38_n_0;
  wire ctl_fetch0_fl_i_39_n_0;
  wire ctl_fetch0_fl_i_3_n_0;
  wire ctl_fetch0_fl_i_40_n_0;
  wire ctl_fetch0_fl_i_41_n_0;
  wire ctl_fetch0_fl_i_43_n_0;
  wire ctl_fetch0_fl_i_45_n_0;
  wire ctl_fetch0_fl_i_4_0;
  wire ctl_fetch0_fl_i_4_1;
  wire ctl_fetch0_fl_i_4_n_0;
  wire ctl_fetch0_fl_i_5_n_0;
  wire ctl_fetch0_fl_i_6_n_0;
  wire ctl_fetch0_fl_i_8_0;
  wire ctl_fetch0_fl_i_8_n_0;
  wire ctl_fetch0_fl_i_9_n_0;
  wire [15:0]ctl_fetch0_fl_reg;
  wire [2:0]ctl_fetch0_fl_reg_0;
  wire ctl_fetch0_fl_reg_1;
  wire ctl_fetch0_fl_reg_2;
  wire ctl_fetch0_fl_reg_3;
  wire ctl_fetch0_fl_reg_4;
  wire ctl_fetch0_fl_reg_5;
  wire ctl_fetch1;
  wire ctl_fetch1_fl;
  wire ctl_fetch1_fl_i_10_n_0;
  wire ctl_fetch1_fl_i_12_n_0;
  wire ctl_fetch1_fl_i_13_n_0;
  wire ctl_fetch1_fl_i_14_n_0;
  wire ctl_fetch1_fl_i_15_n_0;
  wire ctl_fetch1_fl_i_16_0;
  wire ctl_fetch1_fl_i_16_n_0;
  wire ctl_fetch1_fl_i_17_n_0;
  wire ctl_fetch1_fl_i_18_n_0;
  wire ctl_fetch1_fl_i_19_n_0;
  wire [15:0]ctl_fetch1_fl_i_21_0;
  wire ctl_fetch1_fl_i_21_n_0;
  wire ctl_fetch1_fl_i_22_n_0;
  wire ctl_fetch1_fl_i_24_n_0;
  wire ctl_fetch1_fl_i_25_0;
  wire ctl_fetch1_fl_i_25_1;
  wire ctl_fetch1_fl_i_25_n_0;
  wire ctl_fetch1_fl_i_27_0;
  wire ctl_fetch1_fl_i_27_1;
  wire ctl_fetch1_fl_i_27_2;
  wire ctl_fetch1_fl_i_27_n_0;
  wire ctl_fetch1_fl_i_28_n_0;
  wire ctl_fetch1_fl_i_29_n_0;
  wire ctl_fetch1_fl_i_2_0;
  wire ctl_fetch1_fl_i_2_1;
  wire ctl_fetch1_fl_i_2_2;
  wire ctl_fetch1_fl_i_2_3;
  wire ctl_fetch1_fl_i_2_4;
  wire ctl_fetch1_fl_i_2_5;
  wire ctl_fetch1_fl_i_2_6;
  wire ctl_fetch1_fl_i_2_n_0;
  wire ctl_fetch1_fl_i_30_n_0;
  wire ctl_fetch1_fl_i_31_n_0;
  wire ctl_fetch1_fl_i_32_n_0;
  wire ctl_fetch1_fl_i_34_0;
  wire ctl_fetch1_fl_i_34_n_0;
  wire ctl_fetch1_fl_i_35_n_0;
  wire ctl_fetch1_fl_i_37_n_0;
  wire ctl_fetch1_fl_i_39_n_0;
  wire ctl_fetch1_fl_i_3_n_0;
  wire ctl_fetch1_fl_i_4_n_0;
  wire ctl_fetch1_fl_i_5_n_0;
  wire ctl_fetch1_fl_i_7_n_0;
  wire ctl_fetch1_fl_i_8_n_0;
  wire ctl_fetch1_fl_i_9_n_0;
  wire [2:0]ctl_fetch1_fl_reg;
  wire ctl_fetch1_fl_reg_0;
  wire ctl_fetch1_fl_reg_1;
  wire ctl_fetch1_fl_reg_i_6_0;
  wire ctl_fetch1_fl_reg_i_6_1;
  wire ctl_fetch1_fl_reg_i_6_2;
  wire ctl_fetch1_fl_reg_i_6_n_0;
  wire ctl_fetch_ext0;
  wire ctl_fetch_ext_fl;
  wire ctl_sr_ldie0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  wire [15:0]eir;
  wire [15:0]\eir_fl_reg[15] ;
  wire [15:0]\eir_fl_reg[15]_0 ;
  wire eir_inferred_i_17_n_0;
  wire eir_inferred_i_18_n_0;
  wire eir_inferred_i_19_n_0;
  wire eir_inferred_i_20_n_0;
  wire eir_inferred_i_21_n_0;
  wire eir_inferred_i_22_n_0;
  wire eir_inferred_i_23_n_0;
  wire eir_inferred_i_24_n_0;
  wire eir_inferred_i_25_n_0;
  wire eir_inferred_i_26_n_0;
  wire eir_inferred_i_27_n_0;
  wire eir_inferred_i_28_n_0;
  wire eir_inferred_i_29_n_0;
  wire eir_inferred_i_30_n_0;
  wire eir_inferred_i_31_n_0;
  wire eir_inferred_i_32_n_0;
  wire [12:0]fadr;
  wire [3:0]\fadr[12] ;
  wire \fadr[15]_INST_0_i_12_n_0 ;
  wire \fadr[15]_INST_0_i_15_n_0 ;
  wire \fadr[15]_INST_0_i_4_n_0 ;
  wire \fadr[15]_INST_0_i_5_n_0 ;
  wire \fadr[15]_INST_0_i_6_n_0 ;
  wire \fadr[15]_INST_0_i_9_n_0 ;
  wire [3:0]\fadr[8] ;
  wire fadr_1_fl;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[1]_i_2 ;
  wire \fch_irq_lev[1]_i_2_0 ;
  wire fch_irq_req;
  wire fch_irq_req_fl_reg;
  wire fch_issu1;
  wire fch_issu1_fl;
  wire fch_issu1_inferred_i_10_n_0;
  wire fch_issu1_inferred_i_112_n_0;
  wire [10:0]fch_issu1_inferred_i_11_0;
  wire fch_issu1_inferred_i_11_1;
  wire fch_issu1_inferred_i_11_2;
  wire fch_issu1_inferred_i_11_3;
  wire fch_issu1_inferred_i_11_4;
  wire fch_issu1_inferred_i_11_5;
  wire fch_issu1_inferred_i_11_n_0;
  wire fch_issu1_inferred_i_12_n_0;
  wire fch_issu1_inferred_i_13_n_0;
  wire fch_issu1_inferred_i_144_n_0;
  wire fch_issu1_inferred_i_18_n_0;
  wire fch_issu1_inferred_i_19_n_0;
  wire fch_issu1_inferred_i_1_0;
  wire fch_issu1_inferred_i_1_1;
  wire fch_issu1_inferred_i_1_2;
  wire fch_issu1_inferred_i_1_3;
  wire fch_issu1_inferred_i_1_4;
  wire fch_issu1_inferred_i_1_5;
  wire fch_issu1_inferred_i_1_6;
  wire fch_issu1_inferred_i_20_0;
  wire fch_issu1_inferred_i_20_1;
  wire fch_issu1_inferred_i_20_2;
  wire fch_issu1_inferred_i_20_n_0;
  wire fch_issu1_inferred_i_21_n_0;
  wire fch_issu1_inferred_i_22_n_0;
  wire fch_issu1_inferred_i_23_n_0;
  wire fch_issu1_inferred_i_24_n_0;
  wire fch_issu1_inferred_i_28_0;
  wire fch_issu1_inferred_i_28_1;
  wire fch_issu1_inferred_i_28_2;
  wire fch_issu1_inferred_i_28_3;
  wire fch_issu1_inferred_i_28_n_0;
  wire fch_issu1_inferred_i_29_n_0;
  wire fch_issu1_inferred_i_2_0;
  wire fch_issu1_inferred_i_2_1;
  wire fch_issu1_inferred_i_2_2;
  wire fch_issu1_inferred_i_2_n_0;
  wire fch_issu1_inferred_i_30_n_0;
  wire fch_issu1_inferred_i_31_0;
  wire fch_issu1_inferred_i_31_n_0;
  wire fch_issu1_inferred_i_32_0;
  wire fch_issu1_inferred_i_32_1;
  wire fch_issu1_inferred_i_32_2;
  wire fch_issu1_inferred_i_32_n_0;
  wire fch_issu1_inferred_i_33_0;
  wire fch_issu1_inferred_i_33_1;
  wire fch_issu1_inferred_i_33_2;
  wire fch_issu1_inferred_i_33_3;
  wire fch_issu1_inferred_i_33_n_0;
  wire fch_issu1_inferred_i_34_n_0;
  wire fch_issu1_inferred_i_35_n_0;
  wire fch_issu1_inferred_i_38_n_0;
  wire fch_issu1_inferred_i_3_n_0;
  wire fch_issu1_inferred_i_40_n_0;
  wire fch_issu1_inferred_i_41_0;
  wire fch_issu1_inferred_i_41_1;
  wire fch_issu1_inferred_i_41_2;
  wire fch_issu1_inferred_i_41_3;
  wire fch_issu1_inferred_i_41_n_0;
  wire fch_issu1_inferred_i_42_n_0;
  wire fch_issu1_inferred_i_48_n_0;
  wire fch_issu1_inferred_i_4_n_0;
  wire fch_issu1_inferred_i_50_n_0;
  wire fch_issu1_inferred_i_59_n_0;
  wire fch_issu1_inferred_i_5_0;
  wire fch_issu1_inferred_i_5_1;
  wire fch_issu1_inferred_i_5_n_0;
  wire fch_issu1_inferred_i_60_n_0;
  wire fch_issu1_inferred_i_61_n_0;
  wire fch_issu1_inferred_i_6_0;
  wire fch_issu1_inferred_i_6_1;
  wire fch_issu1_inferred_i_6_2;
  wire fch_issu1_inferred_i_6_3;
  wire fch_issu1_inferred_i_6_4;
  wire fch_issu1_inferred_i_6_n_0;
  wire fch_issu1_inferred_i_70_n_0;
  wire fch_issu1_inferred_i_74_n_0;
  wire fch_issu1_inferred_i_75_n_0;
  wire fch_issu1_inferred_i_79_n_0;
  wire fch_issu1_inferred_i_7_0;
  wire fch_issu1_inferred_i_7_1;
  wire fch_issu1_inferred_i_7_2;
  wire fch_issu1_inferred_i_7_3;
  wire fch_issu1_inferred_i_7_4;
  wire fch_issu1_inferred_i_7_5;
  wire fch_issu1_inferred_i_7_6;
  wire fch_issu1_inferred_i_7_n_0;
  wire fch_issu1_inferred_i_80_n_0;
  wire fch_issu1_inferred_i_8_0;
  wire fch_issu1_inferred_i_8_1;
  wire fch_issu1_inferred_i_8_10;
  wire fch_issu1_inferred_i_8_2;
  wire fch_issu1_inferred_i_8_3;
  wire fch_issu1_inferred_i_8_4;
  wire fch_issu1_inferred_i_8_5;
  wire fch_issu1_inferred_i_8_6;
  wire fch_issu1_inferred_i_8_7;
  wire fch_issu1_inferred_i_8_8;
  wire fch_issu1_inferred_i_8_9;
  wire fch_issu1_inferred_i_8_n_0;
  wire fch_issu1_inferred_i_98_n_0;
  wire fch_issu1_inferred_i_9_n_0;
  wire fch_issu1_ir;
  wire fch_leir_hir;
  wire fch_leir_hir_i_2_n_0;
  wire fch_leir_hir_t;
  wire fch_leir_lir;
  wire fch_leir_lir_i_1_n_0;
  wire fch_leir_lir_reg_0;
  wire fch_leir_lir_reg_1;
  wire fch_leir_nir;
  wire fch_leir_nir_reg_0;
  wire fch_leir_nir_reg_1;
  wire fch_leir_nir_t;
  wire fch_memacc1;
  wire fch_term_fl;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire [15:0]fdat;
  wire [15:0]fdatx;
  wire \grn[15]_i_3__1_n_0 ;
  wire [1:0]\grn[15]_i_3__5_0 ;
  wire [1:0]\grn[15]_i_3__5_1 ;
  wire \grn[15]_i_3__5_n_0 ;
  wire \grn[15]_i_3_n_0 ;
  wire \grn[15]_i_5__0_n_0 ;
  wire \grn[15]_i_7_n_0 ;
  wire \grn_reg[15] ;
  wire [2:0]\grn_reg[15]_0 ;
  wire [2:0]\grn_reg[15]_1 ;
  wire [15:0]in0;
  wire \ir0_fl_reg[0] ;
  wire [15:0]\ir0_fl_reg[15] ;
  wire \ir0_id_fl[20]_i_2_n_0 ;
  wire \ir0_id_fl[21]_i_2_n_0 ;
  wire \ir0_id_fl_reg[20] ;
  wire [1:0]\ir0_id_fl_reg[21] ;
  wire ir0_inferred_i_17_n_0;
  wire ir0_inferred_i_18_n_0;
  wire ir0_inferred_i_19_n_0;
  wire ir0_inferred_i_20_n_0;
  wire ir0_inferred_i_21_n_0;
  wire ir0_inferred_i_22_n_0;
  wire ir0_inferred_i_23_n_0;
  wire ir0_inferred_i_24_n_0;
  wire ir0_inferred_i_25_n_0;
  wire ir0_inferred_i_26_n_0;
  wire ir0_inferred_i_27_n_0;
  wire ir0_inferred_i_28_n_0;
  wire ir0_inferred_i_29_n_0;
  wire ir0_inferred_i_30_n_0;
  wire ir0_inferred_i_31_n_0;
  wire ir0_inferred_i_32_n_0;
  wire [15:0]ir1;
  wire \ir1_fl_reg[0] ;
  wire [15:0]\ir1_fl_reg[15] ;
  wire \ir1_id_fl[20]_i_2_n_0 ;
  wire \ir1_id_fl[21]_i_2_n_0 ;
  wire \ir1_id_fl_reg[20] ;
  wire [1:0]\ir1_id_fl_reg[21] ;
  wire [5:0]\ir1_id_fl_reg[21]_0 ;
  wire \ir1_id_fl_reg[21]_1 ;
  wire ir1_inferred_i_18_n_0;
  wire ir1_inferred_i_19_n_0;
  wire ir1_inferred_i_20_n_0;
  wire ir1_inferred_i_21_n_0;
  wire ir1_inferred_i_22_n_0;
  wire ir1_inferred_i_23_n_0;
  wire ir1_inferred_i_24_n_0;
  wire ir1_inferred_i_25_n_0;
  wire ir1_inferred_i_26_n_0;
  wire ir1_inferred_i_27_n_0;
  wire ir1_inferred_i_28_n_0;
  wire ir1_inferred_i_29_n_0;
  wire ir1_inferred_i_30_n_0;
  wire ir1_inferred_i_31_n_0;
  wire ir1_inferred_i_32_n_0;
  wire ir1_inferred_i_33_n_0;
  wire [15:0]\iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire \nir_id[24]_i_3_n_0 ;
  wire \nir_id[24]_i_4_n_0 ;
  wire out;
  wire p_2_in;
  wire [12:0]p_2_in_0;
  wire [12:0]\pc0_reg[12] ;
  wire \pc0_reg[3] ;
  wire \pc[0]_i_2_n_0 ;
  wire \pc[10]_i_2_n_0 ;
  wire \pc[11]_i_2_n_0 ;
  wire \pc[12]_i_4_n_0 ;
  wire \pc[1]_i_2_n_0 ;
  wire \pc[2]_i_2_n_0 ;
  wire \pc[3]_i_2_n_0 ;
  wire \pc[4]_i_4_n_0 ;
  wire \pc[5]_i_3_n_0 ;
  wire \pc[6]_i_2_n_0 ;
  wire \pc[7]_i_2_n_0 ;
  wire \pc[8]_i_4_n_0 ;
  wire \pc[9]_i_2_n_0 ;
  wire \pc_reg[0] ;
  wire [3:0]\pc_reg[11] ;
  wire [0:0]\pc_reg[12] ;
  wire \pc_reg[13] ;
  wire \pc_reg[14] ;
  wire \pc_reg[14]_0 ;
  wire \pc_reg[14]_1 ;
  wire [15:0]\pc_reg[15] ;
  wire [13:0]\pc_reg[15]_0 ;
  wire [15:0]\pc_reg[15]_1 ;
  wire \pc_reg[15]_2 ;
  wire [3:0]\pc_reg[7] ;
  wire \rgf/bank02/grn00/grn1 ;
  wire \rgf/bank02/grn01/grn1 ;
  wire \rgf/bank02/grn02/grn1 ;
  wire \rgf/bank02/grn03/grn1 ;
  wire \rgf/bank02/grn04/grn1 ;
  wire \rgf/bank02/grn05/grn1 ;
  wire \rgf/bank02/grn06/grn1 ;
  wire \rgf/bank02/grn07/grn1 ;
  wire \rgf/bank02/grn20/grn1 ;
  wire \rgf/bank02/grn21/grn1 ;
  wire \rgf/bank02/grn22/grn1 ;
  wire \rgf/bank02/grn23/grn1 ;
  wire \rgf/bank02/grn24/grn1 ;
  wire \rgf/bank02/grn25/grn1 ;
  wire \rgf/bank02/grn26/grn1 ;
  wire \rgf/bank02/grn27/grn1 ;
  wire \rgf/bank13/grn00/grn1 ;
  wire \rgf/bank13/grn01/grn1 ;
  wire \rgf/bank13/grn02/grn1 ;
  wire \rgf/bank13/grn03/grn1 ;
  wire \rgf/bank13/grn04/grn1 ;
  wire \rgf/bank13/grn05/grn1 ;
  wire \rgf/bank13/grn06/grn1 ;
  wire \rgf/bank13/grn07/grn1 ;
  wire \rgf/bank13/grn20/grn1 ;
  wire \rgf/bank13/grn21/grn1 ;
  wire \rgf/bank13/grn22/grn1 ;
  wire \rgf/bank13/grn23/grn1 ;
  wire \rgf/bank13/grn24/grn1 ;
  wire \rgf/bank13/grn25/grn1 ;
  wire \rgf/bank13/grn26/grn1 ;
  wire \rgf/bank13/grn27/grn1 ;
  wire [5:5]\rgf/c0bus_sel_0 ;
  wire [4:1]\rgf/c0bus_sel_cr ;
  wire [4:1]\rgf/c1bus_sel_cr ;
  wire [4:0]\rgf/rctl/p_0_in ;
  wire [0:0]\rgf/rctl/rgf_selc1 ;
  wire [2:0]\rgf/rctl/rgf_selc1_rn ;
  wire [15:0]\rgf/rgf_c0bus_0 ;
  wire [15:0]\rgf/rgf_c1bus_0 ;
  wire rgf_selc0_stat;
  wire rgf_selc1_stat;
  wire [15:0]rgf_selc1_stat_reg;
  wire [15:0]rgf_selc1_stat_reg_0;
  wire [15:0]rgf_selc1_stat_reg_1;
  wire [15:0]rgf_selc1_stat_reg_10;
  wire [15:0]rgf_selc1_stat_reg_11;
  wire [15:0]rgf_selc1_stat_reg_12;
  wire [15:0]rgf_selc1_stat_reg_13;
  wire [15:0]rgf_selc1_stat_reg_14;
  wire [15:0]rgf_selc1_stat_reg_15;
  wire [15:0]rgf_selc1_stat_reg_16;
  wire [15:0]rgf_selc1_stat_reg_17;
  wire [15:0]rgf_selc1_stat_reg_18;
  wire [15:0]rgf_selc1_stat_reg_19;
  wire [15:0]rgf_selc1_stat_reg_2;
  wire [15:0]rgf_selc1_stat_reg_20;
  wire [15:0]rgf_selc1_stat_reg_21;
  wire [15:0]rgf_selc1_stat_reg_22;
  wire [15:0]rgf_selc1_stat_reg_23;
  wire [15:0]rgf_selc1_stat_reg_24;
  wire [15:0]rgf_selc1_stat_reg_25;
  wire [15:0]rgf_selc1_stat_reg_26;
  wire [15:0]rgf_selc1_stat_reg_27;
  wire [15:0]rgf_selc1_stat_reg_28;
  wire [15:0]rgf_selc1_stat_reg_29;
  wire [15:0]rgf_selc1_stat_reg_3;
  wire [15:0]rgf_selc1_stat_reg_30;
  wire [15:0]rgf_selc1_stat_reg_31;
  wire [15:0]rgf_selc1_stat_reg_4;
  wire [15:0]rgf_selc1_stat_reg_5;
  wire [15:0]rgf_selc1_stat_reg_6;
  wire [15:0]rgf_selc1_stat_reg_7;
  wire [15:0]rgf_selc1_stat_reg_8;
  wire [15:0]rgf_selc1_stat_reg_9;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_fl;
  wire rst_n_fl_reg;
  wire rst_n_fl_reg_0;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_2;
  wire [1:0]rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire [15:0]\sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[11]_i_2_n_0 ;
  wire \sr[11]_i_5_n_0 ;
  wire \sr[11]_i_9_n_0 ;
  wire \sr[13]_i_10_n_0 ;
  wire \sr[13]_i_13 ;
  wire \sr[13]_i_2_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire [2:0]\sr[13]_i_5_0 ;
  wire [2:0]\sr[13]_i_5_1 ;
  wire [1:0]\sr[13]_i_5_2 ;
  wire [1:0]\sr[13]_i_5_3 ;
  wire \sr[13]_i_5_n_0 ;
  wire \sr[15]_i_2_n_0 ;
  wire \sr[15]_i_3_n_0 ;
  wire \sr[15]_i_4_n_0 ;
  wire \sr[15]_i_6_n_0 ;
  wire \sr[15]_i_7_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[3]_i_5_n_0 ;
  wire \sr[3]_i_6_n_0 ;
  wire \sr[3]_i_8_n_0 ;
  wire \sr[4]_i_2_n_0 ;
  wire \sr[4]_i_4_n_0 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[5]_i_2_n_0 ;
  wire \sr[5]_i_3_n_0 ;
  wire \sr[5]_i_6_n_0 ;
  wire \sr[6]_i_2_n_0 ;
  wire \sr[6]_i_5_n_0 ;
  wire \sr[7]_i_2_n_0 ;
  wire \sr[7]_i_4_n_0 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_7_n_0 ;
  wire [0:0]\sr_reg[0] ;
  wire [0:0]\sr_reg[0]_0 ;
  wire [0:0]\sr_reg[0]_1 ;
  wire [0:0]\sr_reg[0]_10 ;
  wire [0:0]\sr_reg[0]_11 ;
  wire [0:0]\sr_reg[0]_12 ;
  wire [0:0]\sr_reg[0]_13 ;
  wire [0:0]\sr_reg[0]_14 ;
  wire [0:0]\sr_reg[0]_15 ;
  wire [0:0]\sr_reg[0]_16 ;
  wire [0:0]\sr_reg[0]_17 ;
  wire [0:0]\sr_reg[0]_18 ;
  wire [0:0]\sr_reg[0]_19 ;
  wire [0:0]\sr_reg[0]_2 ;
  wire [0:0]\sr_reg[0]_20 ;
  wire [0:0]\sr_reg[0]_21 ;
  wire [0:0]\sr_reg[0]_22 ;
  wire [0:0]\sr_reg[0]_3 ;
  wire [0:0]\sr_reg[0]_4 ;
  wire [0:0]\sr_reg[0]_5 ;
  wire [0:0]\sr_reg[0]_6 ;
  wire [0:0]\sr_reg[0]_7 ;
  wire [0:0]\sr_reg[0]_8 ;
  wire [0:0]\sr_reg[0]_9 ;
  wire [15:0]\sr_reg[15] ;
  wire [15:0]\sr_reg[15]_0 ;
  wire [0:0]\sr_reg[1] ;
  wire [0:0]\sr_reg[1]_0 ;
  wire [0:0]\sr_reg[1]_1 ;
  wire [0:0]\sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_3 ;
  wire [0:0]\sr_reg[1]_4 ;
  wire [0:0]\sr_reg[1]_5 ;
  wire [0:0]\sr_reg[1]_6 ;
  wire \sr_reg[3] ;
  wire \sr_reg[3]_0 ;
  wire \sr_reg[4] ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[5]_3 ;
  wire \sr_reg[5]_4 ;
  wire \sr_reg[5]_5 ;
  wire \sr_reg[5]_6 ;
  wire \sr_reg[5]_7 ;
  wire \sr_reg[5]_8 ;
  wire \sr_reg[5]_9 ;
  wire \sr_reg[6] ;
  wire [0:0]\sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire [0:0]\sr_reg[7]_1 ;
  wire [2:0]stat;
  wire \stat[0]_i_2__2_n_0 ;
  wire \stat[0]_i_3_n_0 ;
  wire \stat[0]_i_6__0_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3__1_n_0 ;
  wire \stat[1]_i_4_n_0 ;
  wire \stat[2]_i_1__1_n_0 ;
  wire \stat[2]_i_3_n_0 ;
  wire \stat[2]_i_4_0 ;
  wire \stat[2]_i_4_1 ;
  wire \stat[2]_i_4_2 ;
  wire \stat[2]_i_6__1_n_0 ;
  wire [2:0]stat_nx;
  wire \stat_reg[0]_0 ;
  wire [0:0]\stat_reg[0]_1 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire [1:0]\stat_reg[0]_8 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[2]_0 ;
  wire [15:0]\tr_reg[15] ;
  wire [15:0]\tr_reg[15]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_0[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_1[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_2[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_3[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_4[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_5[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_6[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_7[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_8[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_9[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_10[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_11[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_12[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_13[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_14[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_15[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(rgf_selc1_stat_reg_16[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(rgf_selc1_stat_reg_17[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(rgf_selc1_stat_reg_18[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(rgf_selc1_stat_reg_19[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(rgf_selc1_stat_reg_20[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(rgf_selc1_stat_reg_21[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(rgf_selc1_stat_reg_22[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(rgf_selc1_stat_reg_23[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(rgf_selc1_stat_reg_24[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(rgf_selc1_stat_reg_25[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(rgf_selc1_stat_reg_26[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(rgf_selc1_stat_reg_27[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(rgf_selc1_stat_reg_28[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(rgf_selc1_stat_reg_29[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(rgf_selc1_stat_reg_30[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(rgf_selc1_stat_reg_31[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_20 
       (.I0(ctl_fetch0_fl_reg[2]),
        .I1(ctl_fetch0_fl_reg[1]),
        .O(rst_n_fl_reg_4));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[9]_INST_0_i_28 
       (.I0(ctl_fetch1_fl_i_21_0[1]),
        .I1(ctl_fetch1_fl_i_21_0[2]),
        .O(rst_n_fl_reg_1));
  LUT5 #(
    .INIT(32'h00008000)) 
    \ccmd[0]_INST_0_i_20 
       (.I0(ctl_fetch0_fl_reg[9]),
        .I1(ctl_fetch0_fl_reg[8]),
        .I2(ctl_fetch0_fl_reg[11]),
        .I3(ctl_fetch0_fl_reg[10]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .O(\stat_reg[1]_2 ));
  LUT6 #(
    .INIT(64'h00000000EFEEEFEF)) 
    ctl_fetch0_fl_i_1
       (.I0(ctl_fetch0_fl_i_2_n_0),
        .I1(ctl_fetch0_fl_i_3_n_0),
        .I2(ctl_fetch0_fl_reg[11]),
        .I3(ctl_fetch0_fl_i_4_n_0),
        .I4(ctl_fetch0_fl_i_5_n_0),
        .I5(ctl_fetch0_fl_i_6_n_0),
        .O(ctl_fetch0));
  LUT6 #(
    .INIT(64'h00000047FF000047)) 
    ctl_fetch0_fl_i_11
       (.I0(ctl_fetch0_fl_reg[3]),
        .I1(\sr_reg[15]_0 [10]),
        .I2(rst_n_fl_reg_4),
        .I3(ctl_fetch0_fl_reg[14]),
        .I4(ctl_fetch0_fl_reg[12]),
        .I5(ctl_fetch0_fl_reg_0[1]),
        .O(ctl_fetch0_fl_i_11_n_0));
  LUT6 #(
    .INIT(64'hFF04FF04FFFFFF04)) 
    ctl_fetch0_fl_i_12
       (.I0(crdy_0),
        .I1(ctl_fetch0_fl_reg[12]),
        .I2(ctl_fetch0_fl_reg[7]),
        .I3(ctl_fetch0_fl_i_24_n_0),
        .I4(ctl_fetch0_fl_i_25_n_0),
        .I5(\sr_reg[15]_0 [10]),
        .O(ctl_fetch0_fl_i_12_n_0));
  LUT6 #(
    .INIT(64'h000000001111BAAA)) 
    ctl_fetch0_fl_i_13
       (.I0(ctl_fetch0_fl_reg[9]),
        .I1(ctl_fetch0_fl_reg[7]),
        .I2(\sr_reg[15]_0 [11]),
        .I3(crdy),
        .I4(ctl_fetch0_fl_reg[8]),
        .I5(ctl_fetch0_fl_i_26_n_0),
        .O(ctl_fetch0_fl_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000C80000008B00)) 
    ctl_fetch0_fl_i_14
       (.I0(ctl_fetch0_fl_reg[3]),
        .I1(ctl_fetch0_fl_reg[0]),
        .I2(ctl_fetch0_fl_reg[1]),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ctl_fetch0_fl_reg[12]),
        .I5(ctl_fetch0_fl_reg[2]),
        .O(ctl_fetch0_fl_i_14_n_0));
  LUT6 #(
    .INIT(64'hA8AAA8A8AAAAAAAA)) 
    ctl_fetch0_fl_i_15
       (.I0(ctl_fetch0_fl_i_27_n_0),
        .I1(ctl_fetch0_fl_reg_0[2]),
        .I2(ctl_fetch0_fl_reg[15]),
        .I3(crdy_0),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .I5(ctl_fetch0_fl_i_28_n_0),
        .O(ctl_fetch0_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'h0008080808080808)) 
    ctl_fetch0_fl_i_16
       (.I0(ctl_fetch0_fl_i_29_n_0),
        .I1(ctl_fetch0_fl_i_4_0),
        .I2(ctl_fetch0_fl_i_4_1),
        .I3(crdy),
        .I4(ctl_fetch0_fl_reg[0]),
        .I5(ctl_fetch0_fl_i_30_n_0),
        .O(ctl_fetch0_fl_i_16_n_0));
  LUT5 #(
    .INIT(32'h03000055)) 
    ctl_fetch0_fl_i_17
       (.I0(ctl_fetch0_fl_i_31_n_0),
        .I1(ctl_fetch0_fl_reg[6]),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_reg[9]),
        .I4(ctl_fetch0_fl_reg[10]),
        .O(ctl_fetch0_fl_i_17_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_18
       (.I0(\sr[13]_i_13 ),
        .I1(crdy),
        .O(crdy_0));
  LUT6 #(
    .INIT(64'hAEBFAEBAAEEFAEEA)) 
    ctl_fetch0_fl_i_19
       (.I0(ctl_fetch0_fl_i_31_n_0),
        .I1(\sr_reg[15]_0 [7]),
        .I2(ctl_fetch0_fl_reg[14]),
        .I3(ctl_fetch0_fl_reg[13]),
        .I4(\sr_reg[15]_0 [4]),
        .I5(\sr_reg[15]_0 [5]),
        .O(ctl_fetch0_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'h0000FE00FF00FE00)) 
    ctl_fetch0_fl_i_2
       (.I0(ctl_fetch0_fl_reg_1),
        .I1(ctl_fetch0_fl_i_8_n_0),
        .I2(ctl_fetch0_fl_i_9_n_0),
        .I3(ctl_fetch0_fl_reg[11]),
        .I4(ctl_fetch0_fl_reg_2),
        .I5(ctl_fetch0_fl_reg_3),
        .O(ctl_fetch0_fl_i_2_n_0));
  LUT6 #(
    .INIT(64'hF444444444444444)) 
    ctl_fetch0_fl_i_20
       (.I0(ctl_fetch0_fl_i_32_n_0),
        .I1(ctl_fetch0_fl_i_33_n_0),
        .I2(ctl_fetch0_fl_reg[3]),
        .I3(ctl_fetch0_fl_reg[7]),
        .I4(ctl_fetch0_fl_i_34_n_0),
        .I5(\stat_reg[1]_2 ),
        .O(ctl_fetch0_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEEFEE)) 
    ctl_fetch0_fl_i_21
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ctl_fetch0_fl_i_8_0),
        .I2(\sr_reg[15]_0 [6]),
        .I3(ctl_fetch0_fl_reg[13]),
        .I4(ctl_fetch0_fl_reg[12]),
        .I5(ctl_fetch0_fl_i_36_n_0),
        .O(ctl_fetch0_fl_i_21_n_0));
  LUT6 #(
    .INIT(64'h770F770000000000)) 
    ctl_fetch0_fl_i_22
       (.I0(ctl_fetch0_fl_i_37_n_0),
        .I1(ctl_fetch0_fl_reg[5]),
        .I2(ctl_fetch0_fl_i_38_n_0),
        .I3(ctl_fetch0_fl_reg[6]),
        .I4(ctl_fetch0_fl_reg[10]),
        .I5(ctl_fetch0_fl_reg[9]),
        .O(ctl_fetch0_fl_i_22_n_0));
  LUT5 #(
    .INIT(32'hFF0A3000)) 
    ctl_fetch0_fl_i_23
       (.I0(ctl_fetch0_fl_reg[7]),
        .I1(ctl_fetch0_fl_reg[6]),
        .I2(ctl_fetch0_fl_reg[9]),
        .I3(ctl_fetch0_fl_reg[8]),
        .I4(ctl_fetch0_fl_reg[10]),
        .O(ctl_fetch0_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'hE0E0FFFFFFFFFFE0)) 
    ctl_fetch0_fl_i_24
       (.I0(ctl_fetch0_fl_reg[3]),
        .I1(ctl_fetch0_fl_reg[1]),
        .I2(ctl_fetch0_fl_reg_0[1]),
        .I3(ctl_fetch0_fl_reg[7]),
        .I4(ctl_fetch0_fl_reg[12]),
        .I5(ctl_fetch0_fl_reg[13]),
        .O(ctl_fetch0_fl_i_24_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    ctl_fetch0_fl_i_25
       (.I0(ctl_fetch0_fl_reg[9]),
        .I1(ctl_fetch0_fl_reg[8]),
        .I2(crdy),
        .O(ctl_fetch0_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFEFEFEFFFFFEFEF)) 
    ctl_fetch0_fl_i_26
       (.I0(ctl_fetch0_fl_reg_4),
        .I1(ctl_fetch0_fl_reg_0[1]),
        .I2(ctl_fetch0_fl_i_39_n_0),
        .I3(\sr_reg[15]_0 [11]),
        .I4(ctl_fetch0_fl_reg[8]),
        .I5(crdy),
        .O(ctl_fetch0_fl_i_26_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4447)) 
    ctl_fetch0_fl_i_27
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ctl_fetch0_fl_reg[1]),
        .I2(ctl_fetch0_fl_reg[3]),
        .I3(ctl_fetch0_fl_reg[0]),
        .I4(ctl_fetch0_fl_i_40_n_0),
        .I5(ctl_fetch0_fl_i_41_n_0),
        .O(ctl_fetch0_fl_i_27_n_0));
  LUT6 #(
    .INIT(64'hA0FFFFFFA0FFFFE0)) 
    ctl_fetch0_fl_i_28
       (.I0(ctl_fetch0_fl_reg[10]),
        .I1(ctl_fetch0_fl_i_15_0),
        .I2(ctl_fetch0_fl_reg[12]),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_reg_4),
        .I5(\sr[13]_i_13 ),
        .O(ctl_fetch0_fl_i_28_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF4F)) 
    ctl_fetch0_fl_i_29
       (.I0(ctl_fetch0_fl_i_16_0),
        .I1(ctl_fetch0_fl_i_43_n_0),
        .I2(ctl_fetch0_fl_i_16_1),
        .I3(ctl_fetch0_fl_reg_0[1]),
        .I4(ctl_fetch0_fl_reg[1]),
        .I5(ctl_fetch0_fl_reg[2]),
        .O(ctl_fetch0_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    ctl_fetch0_fl_i_3
       (.I0(ctl_fetch0_fl_i_11_n_0),
        .I1(ctl_fetch0_fl_i_12_n_0),
        .I2(ctl_fetch0_fl_reg_0[0]),
        .I3(ctl_fetch0_fl_i_13_n_0),
        .I4(ctl_fetch0_fl_i_14_n_0),
        .I5(ctl_fetch0_fl_i_15_n_0),
        .O(ctl_fetch0_fl_i_3_n_0));
  LUT4 #(
    .INIT(16'hB888)) 
    ctl_fetch0_fl_i_30
       (.I0(ctl_fetch0_fl_reg[3]),
        .I1(\sr_reg[15]_0 [10]),
        .I2(ctl_fetch0_fl_reg[2]),
        .I3(ctl_fetch0_fl_reg[1]),
        .O(ctl_fetch0_fl_i_30_n_0));
  LUT4 #(
    .INIT(16'hE000)) 
    ctl_fetch0_fl_i_31
       (.I0(\sr[13]_i_13 ),
        .I1(\sr_reg[15]_0 [10]),
        .I2(crdy),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .O(ctl_fetch0_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFBBBBBBEFEFEFCF)) 
    ctl_fetch0_fl_i_32
       (.I0(ctl_fetch0_fl_reg_0[1]),
        .I1(ctl_fetch0_fl_reg[8]),
        .I2(ctl_fetch0_fl_i_45_n_0),
        .I3(ctl_fetch0_fl_reg_0[0]),
        .I4(ctl_fetch0_fl_reg[6]),
        .I5(ctl_fetch0_fl_reg[9]),
        .O(ctl_fetch0_fl_i_32_n_0));
  LUT6 #(
    .INIT(64'hE6666666FFFFFFFF)) 
    ctl_fetch0_fl_i_33
       (.I0(ctl_fetch0_fl_reg[10]),
        .I1(ctl_fetch0_fl_reg[11]),
        .I2(ctl_fetch0_fl_reg[7]),
        .I3(ctl_fetch0_fl_reg[6]),
        .I4(ctl_fetch0_fl_reg[5]),
        .I5(ctl_fetch0_fl_reg[8]),
        .O(ctl_fetch0_fl_i_33_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_34
       (.I0(ctl_fetch0_fl_reg[6]),
        .I1(ctl_fetch0_fl_reg[5]),
        .O(ctl_fetch0_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'h04FF040404040404)) 
    ctl_fetch0_fl_i_36
       (.I0(\sr_reg[15]_0 [5]),
        .I1(ctl_fetch0_fl_reg[14]),
        .I2(ctl_fetch0_fl_reg[12]),
        .I3(ctl_fetch0_fl_reg[8]),
        .I4(ctl_fetch0_fl_reg[6]),
        .I5(ctl_fetch0_fl_reg_0[0]),
        .O(ctl_fetch0_fl_i_36_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_37
       (.I0(ctl_fetch0_fl_reg[7]),
        .I1(ctl_fetch0_fl_reg[3]),
        .O(ctl_fetch0_fl_i_37_n_0));
  LUT3 #(
    .INIT(8'h02)) 
    ctl_fetch0_fl_i_38
       (.I0(ctl_fetch0_fl_reg[7]),
        .I1(ctl_fetch0_fl_reg[4]),
        .I2(ctl_fetch0_fl_reg[5]),
        .O(ctl_fetch0_fl_i_38_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_39
       (.I0(ctl_fetch0_fl_reg[12]),
        .I1(ctl_fetch0_fl_reg[10]),
        .O(ctl_fetch0_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'h00FD00CD00310001)) 
    ctl_fetch0_fl_i_4
       (.I0(ctl_fetch0_fl_i_16_n_0),
        .I1(ctl_fetch0_fl_reg[13]),
        .I2(ctl_fetch0_fl_reg[14]),
        .I3(ctl_fetch0_fl_reg[12]),
        .I4(\sr_reg[15]_0 [5]),
        .I5(\sr_reg[15]_0 [6]),
        .O(ctl_fetch0_fl_i_4_n_0));
  LUT5 #(
    .INIT(32'hFFAAFFA8)) 
    ctl_fetch0_fl_i_40
       (.I0(ctl_fetch0_fl_reg_0[2]),
        .I1(ctl_fetch0_fl_reg[10]),
        .I2(ctl_fetch0_fl_reg[3]),
        .I3(ctl_fetch0_fl_reg[15]),
        .I4(ctl_fetch0_fl_reg_0[1]),
        .O(ctl_fetch0_fl_i_40_n_0));
  LUT5 #(
    .INIT(32'hFFAFEFFF)) 
    ctl_fetch0_fl_i_41
       (.I0(ctl_fetch0_fl_reg[9]),
        .I1(ctl_fetch0_fl_reg[3]),
        .I2(ctl_fetch0_fl_i_27_0),
        .I3(ctl_fetch0_fl_reg[0]),
        .I4(ctl_fetch0_fl_reg[2]),
        .O(ctl_fetch0_fl_i_41_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_43
       (.I0(ctl_fetch0_fl_reg[0]),
        .I1(ctl_fetch0_fl_reg[3]),
        .O(ctl_fetch0_fl_i_43_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch0_fl_i_45
       (.I0(ctl_fetch0_fl_reg[10]),
        .I1(ctl_fetch0_fl_reg[11]),
        .I2(ctl_fetch0_fl_reg[7]),
        .O(ctl_fetch0_fl_i_45_n_0));
  LUT6 #(
    .INIT(64'h3333BBBBFFFFFBFF)) 
    ctl_fetch0_fl_i_5
       (.I0(ctl_fetch0_fl_i_17_n_0),
        .I1(ctl_fetch0_fl_reg[12]),
        .I2(crdy_0),
        .I3(ctl_fetch0_fl_reg[8]),
        .I4(ctl_fetch0_fl_reg_4),
        .I5(ctl_fetch0_fl_i_19_n_0),
        .O(ctl_fetch0_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    ctl_fetch0_fl_i_6
       (.I0(ctl_fetch0_fl_i_20_n_0),
        .I1(brdy),
        .I2(ctl_fetch0_fl_reg[14]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(ctl_fetch0_fl_reg[15]),
        .I5(ctl_fetch0_fl_reg_5),
        .O(ctl_fetch0_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEF000000)) 
    ctl_fetch0_fl_i_8
       (.I0(ctl_fetch0_fl_i_2_0),
        .I1(ctl_fetch0_fl_reg[4]),
        .I2(ctl_fetch0_fl_reg[10]),
        .I3(ctl_fetch0_fl_reg[9]),
        .I4(ctl_fetch0_fl_reg_0[0]),
        .I5(ctl_fetch0_fl_i_21_n_0),
        .O(ctl_fetch0_fl_i_8_n_0));
  LUT5 #(
    .INIT(32'hF800F8F8)) 
    ctl_fetch0_fl_i_9
       (.I0(ctl_fetch0_fl_reg[13]),
        .I1(ctl_fetch0_fl_reg[14]),
        .I2(ctl_fetch0_fl_reg_0[2]),
        .I3(ctl_fetch0_fl_i_22_n_0),
        .I4(ctl_fetch0_fl_i_23_n_0),
        .O(ctl_fetch0_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'h5555555504550404)) 
    ctl_fetch1_fl_i_1
       (.I0(ctl_fetch1_fl_i_2_n_0),
        .I1(brdy),
        .I2(\stat_reg[0]_3 ),
        .I3(ctl_fetch1_fl_i_3_n_0),
        .I4(ctl_fetch1_fl_i_4_n_0),
        .I5(ctl_fetch1_fl_i_5_n_0),
        .O(ctl_fetch1));
  LUT6 #(
    .INIT(64'h00000000003E0000)) 
    ctl_fetch1_fl_i_10
       (.I0(ctl_fetch1_fl_i_21_0[1]),
        .I1(ctl_fetch1_fl_i_21_0[3]),
        .I2(ctl_fetch1_fl_i_21_0[0]),
        .I3(ctl_fetch1_fl_i_21_0[9]),
        .I4(ctl_fetch1_fl_i_2_5),
        .I5(ctl_fetch1_fl_i_21_n_0),
        .O(ctl_fetch1_fl_i_10_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch1_fl_i_11
       (.I0(ctl_fetch1_fl_i_21_0[9]),
        .I1(ctl_fetch1_fl_i_21_0[11]),
        .I2(ctl_fetch1_fl_i_21_0[10]),
        .O(rst_n_fl_reg_2));
  LUT2 #(
    .INIT(4'h7)) 
    ctl_fetch1_fl_i_12
       (.I0(ctl_fetch1_fl_i_21_0[6]),
        .I1(ctl_fetch1_fl_i_21_0[3]),
        .O(ctl_fetch1_fl_i_12_n_0));
  LUT6 #(
    .INIT(64'h7F0055FF00FF00FF)) 
    ctl_fetch1_fl_i_13
       (.I0(ctl_fetch1_fl_i_21_0[7]),
        .I1(ctl_fetch1_fl_i_21_0[6]),
        .I2(ctl_fetch1_fl_i_21_0[5]),
        .I3(ctl_fetch1_fl_i_21_0[11]),
        .I4(ctl_fetch1_fl_i_21_0[8]),
        .I5(ctl_fetch1_fl_i_21_0[10]),
        .O(ctl_fetch1_fl_i_13_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch1_fl_i_14
       (.I0(ctl_fetch1_fl_i_21_0[6]),
        .I1(ctl_fetch1_fl_reg[0]),
        .O(ctl_fetch1_fl_i_14_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFB0B0B000)) 
    ctl_fetch1_fl_i_15
       (.I0(ctl_fetch1_fl_i_22_n_0),
        .I1(ctl_fetch1_fl_reg_i_6_2),
        .I2(ctl_fetch1_fl_i_21_0[12]),
        .I3(ctl_fetch1_fl_i_2_0),
        .I4(ctl_fetch1_fl_i_24_n_0),
        .I5(ctl_fetch1_fl_i_25_n_0),
        .O(ctl_fetch1_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'hFFFFFDFF00000100)) 
    ctl_fetch1_fl_i_16
       (.I0(ctl_fetch1_fl_reg_i_6_0),
        .I1(ctl_fetch1_fl_i_21_0[13]),
        .I2(ctl_fetch1_fl_i_21_0[14]),
        .I3(\sr_reg[15]_0 [4]),
        .I4(ctl_fetch1_fl_reg_i_6_1),
        .I5(ctl_fetch1_fl_i_27_n_0),
        .O(ctl_fetch1_fl_i_16_n_0));
  LUT6 #(
    .INIT(64'h4040404340434043)) 
    ctl_fetch1_fl_i_17
       (.I0(ctl_fetch1_fl_reg[1]),
        .I1(ctl_fetch1_fl_i_21_0[12]),
        .I2(ctl_fetch1_fl_i_21_0[14]),
        .I3(ctl_fetch1_fl_i_28_n_0),
        .I4(ctl_fetch1_fl_i_21_0[2]),
        .I5(ctl_fetch1_fl_i_29_n_0),
        .O(ctl_fetch1_fl_i_17_n_0));
  LUT5 #(
    .INIT(32'h30202023)) 
    ctl_fetch1_fl_i_18
       (.I0(ctl_fetch1_fl_i_21_0[3]),
        .I1(ctl_fetch1_fl_i_21_0[12]),
        .I2(ctl_fetch1_fl_i_21_0[0]),
        .I3(ctl_fetch1_fl_i_21_0[2]),
        .I4(ctl_fetch1_fl_i_21_0[1]),
        .O(ctl_fetch1_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0FFE0E0)) 
    ctl_fetch1_fl_i_19
       (.I0(ctl_fetch1_fl_i_21_0[3]),
        .I1(ctl_fetch1_fl_i_21_0[1]),
        .I2(ctl_fetch1_fl_reg[1]),
        .I3(\sr_reg[15]_0 [10]),
        .I4(ctl_fetch1_fl_i_21_0[8]),
        .I5(ctl_fetch1_fl_i_21_0[9]),
        .O(ctl_fetch1_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'h1011101100001011)) 
    ctl_fetch1_fl_i_2
       (.I0(ctl_fetch1_fl_reg_i_6_n_0),
        .I1(ctl_fetch1_fl_i_7_n_0),
        .I2(ctl_fetch1_fl_i_8_n_0),
        .I3(ctl_fetch1_fl_reg[0]),
        .I4(ctl_fetch1_fl_i_9_n_0),
        .I5(ctl_fetch1_fl_i_10_n_0),
        .O(ctl_fetch1_fl_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFBABAFF)) 
    ctl_fetch1_fl_i_21
       (.I0(ctl_fetch1_fl_i_30_n_0),
        .I1(ctl_fetch1_fl_reg[1]),
        .I2(ctl_fetch1_fl_i_21_0[1]),
        .I3(ctl_fetch1_fl_i_21_0[0]),
        .I4(ctl_fetch1_fl_i_21_0[2]),
        .O(ctl_fetch1_fl_i_21_n_0));
  LUT6 #(
    .INIT(64'h8BB8FF338BB8CC00)) 
    ctl_fetch1_fl_i_22
       (.I0(ctl_fetch1_fl_i_21_0[8]),
        .I1(ctl_fetch1_fl_i_21_0[13]),
        .I2(\sr_reg[15]_0 [5]),
        .I3(\sr_reg[15]_0 [7]),
        .I4(ctl_fetch1_fl_i_21_0[14]),
        .I5(\sr_reg[15]_0 [4]),
        .O(ctl_fetch1_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFEFFFEFFF00FF0)) 
    ctl_fetch1_fl_i_24
       (.I0(\sr_reg[15]_0 [10]),
        .I1(ctl_fetch1_fl_i_2_4),
        .I2(ctl_fetch1_fl_i_21_0[10]),
        .I3(ctl_fetch1_fl_i_21_0[9]),
        .I4(ctl_fetch1_fl_i_21_0[6]),
        .I5(ctl_fetch1_fl_reg[0]),
        .O(ctl_fetch1_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'h00FD00CD00310001)) 
    ctl_fetch1_fl_i_25
       (.I0(ctl_fetch1_fl_i_31_n_0),
        .I1(ctl_fetch1_fl_i_21_0[13]),
        .I2(ctl_fetch1_fl_i_21_0[14]),
        .I3(ctl_fetch1_fl_i_21_0[12]),
        .I4(\sr_reg[15]_0 [5]),
        .I5(\sr_reg[15]_0 [6]),
        .O(ctl_fetch1_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFBAAAFFFFFFFF)) 
    ctl_fetch1_fl_i_27
       (.I0(ctl_fetch1_fl_i_32_n_0),
        .I1(ctl_fetch1_fl_i_21_0[8]),
        .I2(ctl_fetch1_fl_i_21_0[6]),
        .I3(ctl_fetch1_fl_reg[0]),
        .I4(ctl_fetch1_fl_i_16_0),
        .I5(ctl_fetch1_fl_i_34_n_0),
        .O(ctl_fetch1_fl_i_27_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_28
       (.I0(ctl_fetch1_fl_i_21_0[3]),
        .I1(\sr_reg[15]_0 [10]),
        .O(ctl_fetch1_fl_i_28_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_29
       (.I0(ctl_fetch1_fl_i_21_0[1]),
        .I1(\sr_reg[15]_0 [10]),
        .O(ctl_fetch1_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    ctl_fetch1_fl_i_3
       (.I0(rst_n_fl_reg_2),
        .I1(ctl_fetch1_fl_i_12_n_0),
        .I2(ctl_fetch1_fl_i_21_0[7]),
        .I3(ctl_fetch1_fl_i_21_0[5]),
        .I4(ctl_fetch1_fl_reg[1]),
        .I5(ctl_fetch1_fl_i_21_0[8]),
        .O(ctl_fetch1_fl_i_3_n_0));
  LUT5 #(
    .INIT(32'hFFAAFFA8)) 
    ctl_fetch1_fl_i_30
       (.I0(ctl_fetch1_fl_reg[2]),
        .I1(ctl_fetch1_fl_i_21_0[10]),
        .I2(ctl_fetch1_fl_i_21_0[3]),
        .I3(ctl_fetch1_fl_i_21_0[15]),
        .I4(ctl_fetch1_fl_reg[1]),
        .O(ctl_fetch1_fl_i_30_n_0));
  LUT6 #(
    .INIT(64'h00000000000077F7)) 
    ctl_fetch1_fl_i_31
       (.I0(ctl_fetch1_fl_reg_i_6_0),
        .I1(rst_n_fl_reg_1),
        .I2(ctl_fetch1_fl_i_25_0),
        .I3(ctl_fetch0_fl_i_16_0),
        .I4(ctl_fetch1_fl_i_35_n_0),
        .I5(ctl_fetch1_fl_i_25_1),
        .O(ctl_fetch1_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFD000FF00)) 
    ctl_fetch1_fl_i_32
       (.I0(ctl_fetch1_fl_i_37_n_0),
        .I1(ctl_fetch1_fl_i_27_2),
        .I2(ctl_fetch1_fl_i_21_0[9]),
        .I3(ctl_fetch1_fl_reg[0]),
        .I4(ctl_fetch1_fl_i_21_0[7]),
        .I5(ctl_fetch1_fl_reg[1]),
        .O(ctl_fetch1_fl_i_32_n_0));
  LUT6 #(
    .INIT(64'h4F444F4F4F444F44)) 
    ctl_fetch1_fl_i_34
       (.I0(ctl_fetch1_fl_reg[2]),
        .I1(ctl_fetch1_fl_i_2_0),
        .I2(ctl_fetch1_fl_i_39_n_0),
        .I3(ctl_fetch1_fl_i_27_0),
        .I4(ctl_fetch1_fl_i_27_1),
        .I5(ctl_fetch1_fl_i_2_1),
        .O(ctl_fetch1_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'hFEFEFAFABAAAAAAA)) 
    ctl_fetch1_fl_i_35
       (.I0(ctl_fetch1_fl_i_21_0[6]),
        .I1(\sr_reg[15]_0 [10]),
        .I2(ctl_fetch1_fl_i_21_0[1]),
        .I3(ctl_fetch1_fl_i_21_0[2]),
        .I4(ctl_fetch1_fl_i_21_0[0]),
        .I5(ctl_fetch1_fl_i_21_0[3]),
        .O(ctl_fetch1_fl_i_35_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_37
       (.I0(ctl_fetch1_fl_i_21_0[10]),
        .I1(ctl_fetch1_fl_i_21_0[3]),
        .O(ctl_fetch1_fl_i_37_n_0));
  LUT6 #(
    .INIT(64'h005500550055FCFF)) 
    ctl_fetch1_fl_i_39
       (.I0(ctl_fetch1_fl_i_21_0[8]),
        .I1(ctl_fetch1_fl_i_21_0[4]),
        .I2(ctl_fetch1_fl_i_21_0[5]),
        .I3(ctl_fetch1_fl_i_21_0[7]),
        .I4(ctl_fetch1_fl_i_21_0[6]),
        .I5(ctl_fetch1_fl_i_34_0),
        .O(ctl_fetch1_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEF676767)) 
    ctl_fetch1_fl_i_4
       (.I0(ctl_fetch1_fl_i_21_0[9]),
        .I1(ctl_fetch1_fl_i_21_0[8]),
        .I2(ctl_fetch1_fl_i_21_0[10]),
        .I3(ctl_fetch1_fl_reg[0]),
        .I4(ctl_fetch1_fl_i_21_0[6]),
        .I5(ctl_fetch1_fl_i_13_n_0),
        .O(ctl_fetch1_fl_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFD0FFFFFFFF)) 
    ctl_fetch1_fl_i_5
       (.I0(ctl_fetch1_fl_i_14_n_0),
        .I1(ctl_fetch1_fl_i_21_0[8]),
        .I2(ctl_fetch1_fl_reg[1]),
        .I3(ctl_fetch1_fl_reg[2]),
        .I4(ctl_fetch1_fl_reg_0),
        .I5(ctl_fetch1_fl_reg_1),
        .O(ctl_fetch1_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'h000001BA00000000)) 
    ctl_fetch1_fl_i_7
       (.I0(ctl_fetch1_fl_i_21_0[9]),
        .I1(ctl_fetch1_fl_i_21_0[7]),
        .I2(\sr_reg[15]_0 [11]),
        .I3(ctl_fetch1_fl_i_21_0[8]),
        .I4(ctl_fetch1_fl_i_2_2),
        .I5(ctl_fetch1_fl_i_2_3),
        .O(ctl_fetch1_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000000020000002)) 
    ctl_fetch1_fl_i_8
       (.I0(ctl_fetch1_fl_i_17_n_0),
        .I1(ctl_fetch1_fl_i_18_n_0),
        .I2(ctl_fetch1_fl_i_21_0[13]),
        .I3(ctl_fetch1_fl_i_21_0[12]),
        .I4(ctl_fetch1_fl_i_21_0[7]),
        .I5(ctl_fetch1_fl_i_19_n_0),
        .O(ctl_fetch1_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'h00015555FFFFFFFF)) 
    ctl_fetch1_fl_i_9
       (.I0(ctl_fetch1_fl_i_2_0),
        .I1(ctl_fetch1_fl_i_2_1),
        .I2(ctl_fetch1_fl_i_21_0[10]),
        .I3(ctl_fetch1_fl_i_2_4),
        .I4(ctl_fetch1_fl_i_21_0[12]),
        .I5(ctl_fetch1_fl_i_2_6),
        .O(ctl_fetch1_fl_i_9_n_0));
  MUXF7 ctl_fetch1_fl_reg_i_6
       (.I0(ctl_fetch1_fl_i_15_n_0),
        .I1(ctl_fetch1_fl_i_16_n_0),
        .O(ctl_fetch1_fl_reg_i_6_n_0),
        .S(ctl_fetch1_fl_i_21_0[11]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_1
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [15]),
        .I2(eir_inferred_i_17_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [15]),
        .O(eir[15]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_10
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [6]),
        .I2(eir_inferred_i_26_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [6]),
        .O(eir[6]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_11
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [5]),
        .I2(eir_inferred_i_27_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [5]),
        .O(eir[5]));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_12
       (.I0(rst_n_fl),
        .I1(eir_inferred_i_28_n_0),
        .I2(ctl_fetch_ext_fl),
        .I3(fch_leir_nir),
        .I4(\eir_fl_reg[15] [4]),
        .I5(\eir_fl_reg[15]_0 [4]),
        .O(eir[4]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_13
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [3]),
        .I2(eir_inferred_i_29_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [3]),
        .O(eir[3]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_14
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [2]),
        .I2(eir_inferred_i_30_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [2]),
        .O(eir[2]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_15
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [1]),
        .I2(eir_inferred_i_31_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [1]),
        .O(eir[1]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_16
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [0]),
        .I2(eir_inferred_i_32_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [0]),
        .O(eir[0]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_17
       (.I0(fdat[15]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [15]),
        .I3(fch_leir_hir),
        .I4(fdatx[15]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_18
       (.I0(fdat[14]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [14]),
        .I3(fch_leir_hir),
        .I4(fdatx[14]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_19
       (.I0(fdat[13]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [13]),
        .I3(fdatx[13]),
        .I4(fch_leir_hir),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_2
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [14]),
        .I2(eir_inferred_i_18_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [14]),
        .O(eir[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_20
       (.I0(fdat[12]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [12]),
        .I3(fdatx[12]),
        .I4(fch_leir_hir),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_21
       (.I0(fdat[11]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [11]),
        .I3(fch_leir_hir),
        .I4(fdatx[11]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_22
       (.I0(fdat[10]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [10]),
        .I3(fch_leir_hir),
        .I4(fdatx[10]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_23
       (.I0(fdat[9]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [9]),
        .I3(fch_leir_hir),
        .I4(fdatx[9]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_24
       (.I0(fdat[8]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [8]),
        .I3(fch_leir_hir),
        .I4(fdatx[8]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_25
       (.I0(fdat[7]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [7]),
        .I3(fch_leir_hir),
        .I4(fdatx[7]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_26
       (.I0(fdat[6]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [6]),
        .I3(fch_leir_hir),
        .I4(fdatx[6]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_27
       (.I0(fdat[5]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [5]),
        .I3(fch_leir_hir),
        .I4(fdatx[5]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_28
       (.I0(fdat[4]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [4]),
        .I3(fdatx[4]),
        .I4(fch_leir_hir),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_29
       (.I0(fdat[3]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [3]),
        .I3(fch_leir_hir),
        .I4(fdatx[3]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_3
       (.I0(rst_n_fl),
        .I1(eir_inferred_i_19_n_0),
        .I2(ctl_fetch_ext_fl),
        .I3(fch_leir_nir),
        .I4(\eir_fl_reg[15] [13]),
        .I5(\eir_fl_reg[15]_0 [13]),
        .O(eir[13]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_30
       (.I0(fdat[2]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [2]),
        .I3(fch_leir_hir),
        .I4(fdatx[2]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_31
       (.I0(fdat[1]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [1]),
        .I3(fch_leir_hir),
        .I4(fdatx[1]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_32
       (.I0(fdat[0]),
        .I1(fch_leir_lir),
        .I2(\eir_fl_reg[15]_0 [0]),
        .I3(fch_leir_hir),
        .I4(fdatx[0]),
        .I5(fch_leir_nir),
        .O(eir_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_4
       (.I0(rst_n_fl),
        .I1(eir_inferred_i_20_n_0),
        .I2(ctl_fetch_ext_fl),
        .I3(fch_leir_nir),
        .I4(\eir_fl_reg[15] [12]),
        .I5(\eir_fl_reg[15]_0 [12]),
        .O(eir[12]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_5
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [11]),
        .I2(eir_inferred_i_21_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [11]),
        .O(eir[11]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_6
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [10]),
        .I2(eir_inferred_i_22_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [10]),
        .O(eir[10]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_7
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [9]),
        .I2(eir_inferred_i_23_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [9]),
        .O(eir[9]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_8
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [8]),
        .I2(eir_inferred_i_24_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [8]),
        .O(eir[8]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_9
       (.I0(fch_leir_nir),
        .I1(\eir_fl_reg[15] [7]),
        .I2(eir_inferred_i_25_n_0),
        .I3(rst_n_fl),
        .I4(ctl_fetch_ext_fl),
        .I5(\eir_fl_reg[15]_0 [7]),
        .O(eir[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \fadr[0]_INST_0 
       (.I0(p_2_in_0[0]),
        .I1(\stat_reg[0]_0 ),
        .I2(\pc0_reg[12] [0]),
        .O(fadr[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[10]_INST_0 
       (.I0(p_2_in_0[10]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[12] [1]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [10]),
        .O(fadr[10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[11]_INST_0 
       (.I0(p_2_in_0[11]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[12] [2]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [11]),
        .O(fadr[11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[12]_INST_0 
       (.I0(p_2_in_0[12]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[12] [3]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [12]),
        .O(fadr[12]));
  LUT6 #(
    .INIT(64'h000000000000002F)) 
    \fadr[15]_INST_0_i_1 
       (.I0(brdy_0),
        .I1(\stat_reg[0]_2 ),
        .I2(\fadr[15]_INST_0_i_4_n_0 ),
        .I3(stat[0]),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(stat[1]),
        .O(\stat_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \fadr[15]_INST_0_i_10 
       (.I0(ctl_fetch1_fl_i_21_0[8]),
        .I1(ctl_fetch1_fl_i_21_0[6]),
        .I2(\fch_irq_lev[1]_i_2 ),
        .I3(\fch_irq_lev[1]_i_2_0 ),
        .I4(ctl_fetch1_fl_i_21_0[10]),
        .I5(ctl_fetch1_fl_i_21_0[9]),
        .O(rst_n_fl_reg_0));
  LUT4 #(
    .INIT(16'h0004)) 
    \fadr[15]_INST_0_i_12 
       (.I0(ctl_fetch0_fl_reg[2]),
        .I1(ctl_fetch0_fl_reg[0]),
        .I2(ctl_fetch0_fl_reg[15]),
        .I3(ctl_fetch0_fl_reg[14]),
        .O(\fadr[15]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \fadr[15]_INST_0_i_15 
       (.I0(ctl_fetch1_fl_i_21_0[0]),
        .I1(ctl_fetch1_fl_i_21_0[1]),
        .O(\fadr[15]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \fadr[15]_INST_0_i_2 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(stat[1]),
        .I2(\fadr[15]_INST_0_i_6_n_0 ),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h5555555455555555)) 
    \fadr[15]_INST_0_i_4 
       (.I0(ctl_fetch_ext0),
        .I1(\fadr[15]_INST_0_i_9_n_0 ),
        .I2(ctl_fetch1_fl_i_21_0[12]),
        .I3(ctl_fetch1_fl_i_21_0[11]),
        .I4(ctl_fetch1_fl_i_21_0[13]),
        .I5(rst_n_fl_reg_0),
        .O(\fadr[15]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h04FF)) 
    \fadr[15]_INST_0_i_5 
       (.I0(fch_leir_lir_reg_0),
        .I1(fch_leir_lir_reg_1),
        .I2(\fadr[15]_INST_0_i_4_n_0 ),
        .I3(rst_n_fl),
        .O(\fadr[15]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFFDF0FFFF)) 
    \fadr[15]_INST_0_i_6 
       (.I0(brdy_0),
        .I1(\stat_reg[0]_2 ),
        .I2(stat[0]),
        .I3(\stat_reg[2]_0 ),
        .I4(fch_issu1_ir),
        .I5(stat[2]),
        .O(\fadr[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \fadr[15]_INST_0_i_8 
       (.I0(\stat[2]_i_4_0 ),
        .I1(\fadr[15]_INST_0_i_12_n_0 ),
        .I2(ctl_fetch0_fl_reg[1]),
        .I3(ctl_fetch0_fl_reg_0[2]),
        .I4(\stat[2]_i_4_1 ),
        .I5(\stat[2]_i_4_2 ),
        .O(ctl_fetch_ext0));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFFFF)) 
    \fadr[15]_INST_0_i_9 
       (.I0(fch_leir_nir_reg_0),
        .I1(ctl_fetch1_fl_i_21_0[4]),
        .I2(ctl_fetch1_fl_i_21_0[3]),
        .I3(ctl_fetch1_fl_reg[2]),
        .I4(ctl_fetch1_fl_i_21_0[2]),
        .I5(\fadr[15]_INST_0_i_15_n_0 ),
        .O(\fadr[15]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[1]_INST_0 
       (.I0(p_2_in_0[1]),
        .I1(\stat_reg[0]_0 ),
        .I2(O[0]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [1]),
        .O(fadr[1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[2]_INST_0 
       (.I0(p_2_in_0[2]),
        .I1(\stat_reg[0]_0 ),
        .I2(O[1]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [2]),
        .O(fadr[2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[3]_INST_0 
       (.I0(p_2_in_0[3]),
        .I1(\stat_reg[0]_0 ),
        .I2(O[2]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [3]),
        .O(fadr[3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[4]_INST_0 
       (.I0(p_2_in_0[4]),
        .I1(\stat_reg[0]_0 ),
        .I2(O[3]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [4]),
        .O(fadr[4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[5]_INST_0 
       (.I0(p_2_in_0[5]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[8] [0]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [5]),
        .O(fadr[5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[6]_INST_0 
       (.I0(p_2_in_0[6]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[8] [1]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [6]),
        .O(fadr[6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[7]_INST_0 
       (.I0(p_2_in_0[7]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[8] [2]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [7]),
        .O(fadr[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[8]_INST_0 
       (.I0(p_2_in_0[8]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[8] [3]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [8]),
        .O(fadr[8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[9]_INST_0 
       (.I0(p_2_in_0[9]),
        .I1(\stat_reg[0]_0 ),
        .I2(\fadr[12] [0]),
        .I3(\stat_reg[1]_1 ),
        .I4(\pc0_reg[12] [9]),
        .O(fadr[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    fch_issu1_fl_i_1
       (.I0(out),
        .I1(fch_term_fl),
        .I2(fch_issu1_fl),
        .O(fch_issu1_ir));
  LUT6 #(
    .INIT(64'hAA82AA82A0800A02)) 
    fch_issu1_inferred_i_1
       (.I0(fch_issu1_inferred_i_2_n_0),
        .I1(fch_issu1_inferred_i_3_n_0),
        .I2(fch_issu1_inferred_i_4_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_6_n_0),
        .I5(fch_issu1_inferred_i_7_n_0),
        .O(fch_issu1));
  LUT6 #(
    .INIT(64'h35353F3F3535303F)) 
    fch_issu1_inferred_i_10
       (.I0(\ir1_id_fl_reg[21]_0 [3]),
        .I1(fch_issu1_inferred_i_11_0[7]),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fch_issu1_inferred_i_2_1),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_2_2),
        .O(fch_issu1_inferred_i_10_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00AB)) 
    fch_issu1_inferred_i_11
       (.I0(fch_issu1_inferred_i_38_n_0),
        .I1(fdatx[15]),
        .I2(fch_issu1_inferred_i_2_0),
        .I3(fch_issu1_inferred_i_40_n_0),
        .I4(\sr_reg[15]_0 [9]),
        .I5(fch_issu1_inferred_i_41_n_0),
        .O(fch_issu1_inferred_i_11_n_0));
  LUT4 #(
    .INIT(16'h0D00)) 
    fch_issu1_inferred_i_112
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(fadr_1_fl),
        .I3(fdat[8]),
        .O(fch_issu1_inferred_i_112_n_0));
  LUT5 #(
    .INIT(32'h00000990)) 
    fch_issu1_inferred_i_12
       (.I0(fch_issu1_inferred_i_28_n_0),
        .I1(fch_issu1_inferred_i_34_n_0),
        .I2(fch_issu1_inferred_i_29_n_0),
        .I3(fch_issu1_inferred_i_33_n_0),
        .I4(fch_issu1_inferred_i_42_n_0),
        .O(fch_issu1_inferred_i_12_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_13
       (.I0(stat[1]),
        .I1(stat[0]),
        .O(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'h444F444F444F4444)) 
    fch_issu1_inferred_i_144
       (.I0(stat[0]),
        .I1(stat[1]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[12]),
        .O(fch_issu1_inferred_i_144_n_0));
  LUT6 #(
    .INIT(64'h0700F7FFF7FFF7FF)) 
    fch_issu1_inferred_i_18
       (.I0(fch_issu1_inferred_i_5_0),
        .I1(fdatx[0]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdat[0]),
        .I5(fch_issu1_inferred_i_5_1),
        .O(fch_issu1_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000FF0FBB0BBB0B)) 
    fch_issu1_inferred_i_19
       (.I0(fch_issu1_inferred_i_8_0),
        .I1(fadr_1_fl),
        .I2(fch_issu1_inferred_i_48_n_0),
        .I3(fch_issu1_inferred_i_8_1),
        .I4(fch_issu1_inferred_i_11_0[0]),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h000000000000A88A)) 
    fch_issu1_inferred_i_2
       (.I0(fch_issu1_inferred_i_8_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_3_n_0),
        .I4(fch_issu1_inferred_i_11_n_0),
        .I5(fch_issu1_inferred_i_12_n_0),
        .O(fch_issu1_inferred_i_2_n_0));
  LUT6 #(
    .INIT(64'h0B0B000F0B0B0B0B)) 
    fch_issu1_inferred_i_20
       (.I0(fch_issu1_inferred_i_8_2),
        .I1(fadr_1_fl),
        .I2(fch_issu1_inferred_i_50_n_0),
        .I3(fch_issu1_inferred_i_11_0[2]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hBFBBB0BBBFBBBFBB)) 
    fch_issu1_inferred_i_21
       (.I0(fdat[2]),
        .I1(fch_issu1_inferred_i_5_1),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_5_0),
        .O(fch_issu1_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h0FBB0FBB00000FBB)) 
    fch_issu1_inferred_i_22
       (.I0(fch_issu1_inferred_i_8_9),
        .I1(fadr_1_fl),
        .I2(fch_issu1_inferred_i_11_0[1]),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_48_n_0),
        .I5(fch_issu1_inferred_i_8_10),
        .O(fch_issu1_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hF0BBF0F0FFBBFFFF)) 
    fch_issu1_inferred_i_23
       (.I0(fdatx[1]),
        .I1(fch_issu1_inferred_i_5_0),
        .I2(fdat[1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_5_1),
        .O(fch_issu1_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hD0D0D0D0D000D0D0)) 
    fch_issu1_inferred_i_24
       (.I0(fch_issu1_inferred_i_6_1),
        .I1(fch_issu1_inferred_i_6_2),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fch_issu1_inferred_i_6_3),
        .I4(fch_issu1_inferred_i_6_0),
        .I5(fch_issu1_inferred_i_6_4),
        .O(fch_issu1_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h0001010101010101)) 
    fch_issu1_inferred_i_28
       (.I0(fch_issu1_inferred_i_59_n_0),
        .I1(fch_issu1_inferred_i_60_n_0),
        .I2(fch_issu1_inferred_i_61_n_0),
        .I3(fch_issu1_inferred_i_7_0),
        .I4(fch_issu1_inferred_i_6_0),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hACACACACAFAFACAF)) 
    fch_issu1_inferred_i_29
       (.I0(fch_issu1_inferred_i_7_1),
        .I1(fch_issu1_inferred_i_7_2),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fch_issu1_inferred_i_7_3),
        .I4(fdat[10]),
        .I5(fch_issu1_inferred_i_7_4),
        .O(fch_issu1_inferred_i_29_n_0));
  MUXF7 fch_issu1_inferred_i_3
       (.I0(fch_issu1_inferred_i_1_3),
        .I1(fch_issu1_inferred_i_1_4),
        .O(fch_issu1_inferred_i_3_n_0),
        .S(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'h0300AAAAFFFFAAAA)) 
    fch_issu1_inferred_i_30
       (.I0(fch_issu1_inferred_i_7_5),
        .I1(fdatx[9]),
        .I2(fch_issu1_inferred_i_33_3),
        .I3(fch_issu1_inferred_i_6_1),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fch_issu1_inferred_i_7_6),
        .O(fch_issu1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h00000000EEEEEE0E)) 
    fch_issu1_inferred_i_31
       (.I0(fch_issu1_inferred_i_70_n_0),
        .I1(fch_issu1_inferred_i_8_3),
        .I2(fch_issu1_inferred_i_8_4),
        .I3(fch_issu1_inferred_i_8_5),
        .I4(fch_issu1_inferred_i_74_n_0),
        .I5(fch_issu1_inferred_i_75_n_0),
        .O(fch_issu1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    fch_issu1_inferred_i_32
       (.I0(fch_issu1_inferred_i_74_n_0),
        .I1(fch_issu1_inferred_i_8_6),
        .I2(fch_issu1_inferred_i_8_7),
        .I3(fch_issu1_inferred_i_8_8),
        .I4(fch_issu1_inferred_i_79_n_0),
        .I5(fch_issu1_inferred_i_75_n_0),
        .O(fch_issu1_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h00000000770F7777)) 
    fch_issu1_inferred_i_33
       (.I0(fadr_1_fl),
        .I1(\ir1_id_fl_reg[21]_0 [2]),
        .I2(fch_issu1_inferred_i_11_0[6]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fch_issu1_inferred_i_80_n_0),
        .O(fch_issu1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h35353F3F3535303F)) 
    fch_issu1_inferred_i_34
       (.I0(\ir1_id_fl_reg[21]_0 [0]),
        .I1(fch_issu1_inferred_i_11_0[4]),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fch_issu1_inferred_i_41_2),
        .I4(fadr_1_fl),
        .I5(fch_issu1_inferred_i_41_3),
        .O(fch_issu1_inferred_i_34_n_0));
  LUT6 #(
    .INIT(64'h005F005CFF5FFF5C)) 
    fch_issu1_inferred_i_35
       (.I0(\ir1_id_fl_reg[21]_0 [1]),
        .I1(fch_issu1_inferred_i_41_0),
        .I2(fadr_1_fl),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_41_1),
        .I5(fch_issu1_inferred_i_11_0[5]),
        .O(fch_issu1_inferred_i_35_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF0D)) 
    fch_issu1_inferred_i_38
       (.I0(fch_issu1_inferred_i_11_3),
        .I1(fch_issu1_inferred_i_11_4),
        .I2(fdat[15]),
        .I3(fadr_1_fl),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fch_issu1_inferred_i_11_5),
        .O(fch_issu1_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hF3A200A2FFAE0CAE)) 
    fch_issu1_inferred_i_4
       (.I0(fch_issu1_inferred_i_1_5),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fch_issu1_inferred_i_1_6),
        .I5(fch_issu1_inferred_i_11_0[3]),
        .O(fch_issu1_inferred_i_4_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB80000)) 
    fch_issu1_inferred_i_40
       (.I0(fch_issu1_inferred_i_11_1),
        .I1(fdatx[12]),
        .I2(fch_issu1_inferred_i_11_2),
        .I3(fdatx[15]),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fch_issu1_inferred_i_11_0[10]),
        .O(fch_issu1_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'h0900000000000900)) 
    fch_issu1_inferred_i_41
       (.I0(fch_issu1_inferred_i_32_n_0),
        .I1(fch_issu1_inferred_i_35_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_34_n_0),
        .I4(fch_issu1_inferred_i_33_n_0),
        .I5(fch_issu1_inferred_i_31_n_0),
        .O(fch_issu1_inferred_i_41_n_0));
  LUT4 #(
    .INIT(16'hF66F)) 
    fch_issu1_inferred_i_42
       (.I0(fch_issu1_inferred_i_35_n_0),
        .I1(fch_issu1_inferred_i_30_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_6_n_0),
        .O(fch_issu1_inferred_i_42_n_0));
  LUT6 #(
    .INIT(64'h82AAA2AA80AA80AA)) 
    fch_issu1_inferred_i_48
       (.I0(fch_issu1_inferred_i_98_n_0),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .I3(fdatx[15]),
        .I4(fdatx[11]),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_48_n_0));
  LUT6 #(
    .INIT(64'hFFFFF66FF66FFFFF)) 
    fch_issu1_inferred_i_5
       (.I0(fch_issu1_inferred_i_18_n_0),
        .I1(fch_issu1_inferred_i_19_n_0),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(fch_issu1_inferred_i_21_n_0),
        .I4(fch_issu1_inferred_i_22_n_0),
        .I5(fch_issu1_inferred_i_23_n_0),
        .O(fch_issu1_inferred_i_5_n_0));
  LUT5 #(
    .INIT(32'h8000AAAA)) 
    fch_issu1_inferred_i_50
       (.I0(fch_issu1_inferred_i_48_n_0),
        .I1(fch_issu1_inferred_i_20_0),
        .I2(fch_issu1_inferred_i_20_1),
        .I3(fdatx[14]),
        .I4(fch_issu1_inferred_i_20_2),
        .O(fch_issu1_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'h0000000022F20000)) 
    fch_issu1_inferred_i_59
       (.I0(fch_issu1_inferred_i_28_0),
        .I1(fch_issu1_inferred_i_28_1),
        .I2(fdat[3]),
        .I3(fch_issu1_inferred_i_28_2),
        .I4(fch_issu1_inferred_i_98_n_0),
        .I5(fch_issu1_inferred_i_28_3),
        .O(fch_issu1_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFAAFB)) 
    fch_issu1_inferred_i_6
       (.I0(fch_issu1_inferred_i_24_n_0),
        .I1(fch_issu1_inferred_i_1_0),
        .I2(fch_issu1_inferred_i_1_1),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_1_2),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'h0080808080808080)) 
    fch_issu1_inferred_i_60
       (.I0(fch_issu1_inferred_i_6_1),
        .I1(fdatx[8]),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .I5(fdatx[13]),
        .O(fch_issu1_inferred_i_60_n_0));
  LUT6 #(
    .INIT(64'h2AAA22AA00000000)) 
    fch_issu1_inferred_i_61
       (.I0(fch_issu1_inferred_i_112_n_0),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fdat[11]),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_61_n_0));
  LUT6 #(
    .INIT(64'hF66FFFFFFFFFF66F)) 
    fch_issu1_inferred_i_7
       (.I0(fch_issu1_inferred_i_28_n_0),
        .I1(fch_issu1_inferred_i_19_n_0),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(fch_issu1_inferred_i_29_n_0),
        .I4(fch_issu1_inferred_i_22_n_0),
        .I5(fch_issu1_inferred_i_30_n_0),
        .O(fch_issu1_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'hF0F0F0FFF0F0F0FE)) 
    fch_issu1_inferred_i_70
       (.I0(fdat[12]),
        .I1(fdat[14]),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fdat[15]),
        .I4(fdat[13]),
        .I5(fch_issu1_inferred_i_31_0),
        .O(fch_issu1_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'hFFFF1110FFFFFFFF)) 
    fch_issu1_inferred_i_74
       (.I0(fdatx[13]),
        .I1(fdatx[15]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(fch_issu1_inferred_i_74_n_0));
  LUT3 #(
    .INIT(8'h8A)) 
    fch_issu1_inferred_i_75
       (.I0(fadr_1_fl),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(fch_issu1_inferred_i_75_n_0));
  LUT6 #(
    .INIT(64'hAEAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_79
       (.I0(fch_issu1_inferred_i_144_n_0),
        .I1(fdat[12]),
        .I2(fdat[15]),
        .I3(fch_issu1_inferred_i_32_0),
        .I4(fch_issu1_inferred_i_32_1),
        .I5(fch_issu1_inferred_i_32_2),
        .O(fch_issu1_inferred_i_79_n_0));
  LUT6 #(
    .INIT(64'hF6FFFFFFFFFFF6FF)) 
    fch_issu1_inferred_i_8
       (.I0(fch_issu1_inferred_i_31_n_0),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(fch_issu1_inferred_i_4_n_0),
        .I3(fch_issu1_inferred_i_19_n_0),
        .I4(fch_issu1_inferred_i_22_n_0),
        .I5(fch_issu1_inferred_i_32_n_0),
        .O(fch_issu1_inferred_i_8_n_0));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E000E0)) 
    fch_issu1_inferred_i_80
       (.I0(fch_issu1_inferred_i_33_0),
        .I1(fch_issu1_inferred_i_33_1),
        .I2(fch_issu1_inferred_i_98_n_0),
        .I3(fch_issu1_inferred_i_33_2),
        .I4(fch_issu1_inferred_i_33_3),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_80_n_0));
  LUT6 #(
    .INIT(64'hFFFF9FF99FF9FFFF)) 
    fch_issu1_inferred_i_9
       (.I0(fch_issu1_inferred_i_21_n_0),
        .I1(fch_issu1_inferred_i_33_n_0),
        .I2(fch_issu1_inferred_i_34_n_0),
        .I3(fch_issu1_inferred_i_18_n_0),
        .I4(fch_issu1_inferred_i_35_n_0),
        .I5(fch_issu1_inferred_i_23_n_0),
        .O(fch_issu1_inferred_i_9_n_0));
  LUT3 #(
    .INIT(8'h45)) 
    fch_issu1_inferred_i_98
       (.I0(fadr_1_fl),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(fch_issu1_inferred_i_98_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF55150000)) 
    fch_leir_hir_i_1
       (.I0(\pc0_reg[12] [1]),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(stat[2]),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(fch_leir_hir_i_2_n_0),
        .O(fch_leir_hir_t));
  LUT6 #(
    .INIT(64'h0000000008020828)) 
    fch_leir_hir_i_2
       (.I0(\stat[2]_i_3_n_0 ),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(stat[2]),
        .I4(fch_issu1_ir),
        .I5(\fadr[15]_INST_0_i_4_n_0 ),
        .O(fch_leir_hir_i_2_n_0));
  FDRE fch_leir_hir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_hir_t),
        .Q(fch_leir_hir),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'h8AAA0000)) 
    fch_leir_lir_i_1
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(stat[2]),
        .I2(stat[1]),
        .I3(stat[0]),
        .I4(\pc0_reg[12] [1]),
        .O(fch_leir_lir_i_1_n_0));
  FDRE fch_leir_lir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_lir_i_1_n_0),
        .Q(fch_leir_lir),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001100101)) 
    fch_leir_nir_i_1
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(stat[2]),
        .I4(fch_issu1_ir),
        .I5(\stat_reg[2]_0 ),
        .O(fch_leir_nir_t));
  FDRE fch_leir_nir_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_leir_nir_t),
        .Q(fch_leir_nir),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    fch_term_fl_i_1
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .O(brdy_0));
  LUT4 #(
    .INIT(16'hAAAE)) 
    \grn[15]_i_1 
       (.I0(\rgf/bank02/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_20 ));
  LUT4 #(
    .INIT(16'hEAAA)) 
    \grn[15]_i_1__0 
       (.I0(\rgf/bank13/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_21 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1__1 
       (.I0(\rgf/bank13/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_22 ));
  LUT5 #(
    .INIT(32'hF0F0F0F1)) 
    \grn[15]_i_1__10 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn03/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__11 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn22/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__12 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn02/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_5 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__13 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn22/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_6 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__14 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn02/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_7 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__15 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn21/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_2 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__16 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn01/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_8 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__17 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn21/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_9 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__18 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn01/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_10 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__19 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn26/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_3 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1__2 
       (.I0(\rgf/bank02/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_6 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__20 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn06/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_11 ));
  LUT6 #(
    .INIT(64'hFF40FF00FF00FF00)) 
    \grn[15]_i_1__21 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn26/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_12 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF40)) 
    \grn[15]_i_1__22 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn06/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_13 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__23 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn24/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_4 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__24 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn04/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_14 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__25 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn24/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_15 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__26 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn04/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_16 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF01FF00)) 
    \grn[15]_i_1__27 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank13/grn00/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_17 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF01FF00)) 
    \grn[15]_i_1__28 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank02/grn20/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_5 ));
  LUT6 #(
    .INIT(64'hFF01FF00FF00FF00)) 
    \grn[15]_i_1__29 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank13/grn20/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_18 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn27/grn1 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF01)) 
    \grn[15]_i_1__30 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank02/grn00/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_19 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__4 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn07/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFF02FF00FF00FF00)) 
    \grn[15]_i_1__5 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn27/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF02)) 
    \grn[15]_i_1__6 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn07/grn1 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__7 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn23/grn1 ),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\sr_reg[15]_0 [0]),
        .O(\sr_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__8 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn03/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_2 ));
  LUT5 #(
    .INIT(32'hF1F0F0F0)) 
    \grn[15]_i_1__9 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn23/grn1 ),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\sr_reg[15]_0 [1]),
        .O(\sr_reg[0]_3 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .O(\grn[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_3__0 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [1]),
        .O(\rgf/rctl/p_0_in [1]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_3__1 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .O(\grn[15]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__10 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__11 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn04/grn1 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \grn[15]_i_3__12 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \grn[15]_i_3__13 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__14 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__15 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \grn[15]_i_3__16 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \grn[15]_i_3__17 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn20/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__18 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn20/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__19 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn00/grn1 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \grn[15]_i_3__2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__20 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__21 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn03/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__22 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__23 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank02/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__24 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank13/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__25 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [0]),
        .I3(\sr_reg[15]_0 [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__26 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__27 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank13/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__28 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__29 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank02/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__30 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h1B1F5F1FFFFFFFFF)) 
    \grn[15]_i_3__5 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn[15]_i_3__5_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_3__5_1 [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\grn[15]_i_3__5_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__6 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [0]),
        .I5(\sr_reg[15]_0 [1]),
        .O(\rgf/bank02/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__7 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn05/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__8 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank13/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_3__9 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn05/grn1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4 
       (.I0(\grn[15]_i_3__5_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/rctl/p_0_in [2]),
        .O(\rgf/c0bus_sel_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__0 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [0]),
        .O(\rgf/rctl/p_0_in [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__1 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn_reg[15]_0 [2]),
        .I3(rgf_selc0_stat),
        .I4(\grn_reg[15]_1 [2]),
        .O(\rgf/rctl/p_0_in [2]));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \grn[15]_i_4__2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_4__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn03/grn1 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_5 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn[15]_i_3__5_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_3__5_1 [1]),
        .O(\rgf/rctl/p_0_in [4]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_5__0 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .O(\grn[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_5__1 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [1]),
        .I3(\sr_reg[15]_0 [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn04/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \grn[15]_i_6 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr_reg[15]_0 [1]),
        .I5(\sr_reg[15]_0 [0]),
        .O(\rgf/bank02/grn00/grn1 ));
  LUT6 #(
    .INIT(64'h1B1F5F1FFFFFFFFF)) 
    \grn[15]_i_7 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[13]_i_5_2 [1]),
        .I3(rgf_selc1_stat),
        .I4(\sr[13]_i_5_3 [1]),
        .I5(\rgf/rctl/rgf_selc1 ),
        .O(\grn[15]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h8880)) 
    \ir0_id_fl[20]_i_1 
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl),
        .I3(\ir0_id_fl_reg[21] [0]),
        .O(rst_n_fl_reg_3[0]));
  LUT6 #(
    .INIT(64'hFFCFFCCCFDCDFDCD)) 
    \ir0_id_fl[20]_i_2 
       (.I0(\ir1_id_fl_reg[20] ),
        .I1(\ir0_id_fl_reg[20] ),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fch_issu1_inferred_i_11_0[8]),
        .I4(\ir1_id_fl_reg[21]_0 [4]),
        .I5(fadr_1_fl),
        .O(\ir0_id_fl[20]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8880)) 
    \ir0_id_fl[21]_i_1 
       (.I0(\ir0_id_fl[21]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl),
        .I3(\ir0_id_fl_reg[21] [1]),
        .O(rst_n_fl_reg_3[1]));
  LUT6 #(
    .INIT(64'hFFCFFCCCFDCDFDCD)) 
    \ir0_id_fl[21]_i_2 
       (.I0(\ir1_id_fl_reg[21]_1 ),
        .I1(\ir0_id_fl_reg[20] ),
        .I2(fch_issu1_inferred_i_13_n_0),
        .I3(fch_issu1_inferred_i_11_0[9]),
        .I4(\ir1_id_fl_reg[21]_0 [5]),
        .I5(fadr_1_fl),
        .O(\ir0_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_1
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_17_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [15]),
        .O(in0[15]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_10
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_26_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [6]),
        .O(in0[6]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_11
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_27_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [5]),
        .O(in0[5]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_12
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_28_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [4]),
        .O(in0[4]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_13
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_29_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [3]),
        .O(in0[3]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_30_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [2]),
        .O(in0[2]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_31_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [1]),
        .O(in0[1]));
  LUT6 #(
    .INIT(64'hAA08AA08AA080008)) 
    ir0_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\ir0_fl_reg[15] [0]),
        .I2(ctl_fetch0_fl),
        .I3(fch_term_fl),
        .I4(ir0_inferred_i_32_n_0),
        .I5(\ir0_fl_reg[0] ),
        .O(in0[0]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_17
       (.I0(\eir_fl_reg[15] [15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[15]),
        .I4(fadr_1_fl),
        .I5(fdatx[15]),
        .O(ir0_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_18
       (.I0(\eir_fl_reg[15] [14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[14]),
        .I4(fadr_1_fl),
        .I5(fdatx[14]),
        .O(ir0_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_19
       (.I0(\eir_fl_reg[15] [13]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[13]),
        .I4(fadr_1_fl),
        .I5(fdatx[13]),
        .O(ir0_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_2
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_18_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [14]),
        .O(in0[14]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_20
       (.I0(\eir_fl_reg[15] [12]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[12]),
        .I4(fadr_1_fl),
        .I5(fdatx[12]),
        .O(ir0_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_21
       (.I0(\eir_fl_reg[15] [11]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[11]),
        .I4(fadr_1_fl),
        .I5(fdatx[11]),
        .O(ir0_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_22
       (.I0(\eir_fl_reg[15] [10]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[10]),
        .I4(fadr_1_fl),
        .I5(fdatx[10]),
        .O(ir0_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_23
       (.I0(\eir_fl_reg[15] [9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[9]),
        .I4(fadr_1_fl),
        .I5(fdatx[9]),
        .O(ir0_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_24
       (.I0(\eir_fl_reg[15] [8]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[8]),
        .I4(fadr_1_fl),
        .I5(fdatx[8]),
        .O(ir0_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_25
       (.I0(\eir_fl_reg[15] [7]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[7]),
        .I4(fadr_1_fl),
        .I5(fdatx[7]),
        .O(ir0_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_26
       (.I0(\eir_fl_reg[15] [6]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[6]),
        .I4(fadr_1_fl),
        .I5(fdatx[6]),
        .O(ir0_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_27
       (.I0(\eir_fl_reg[15] [5]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[5]),
        .I4(fadr_1_fl),
        .I5(fdatx[5]),
        .O(ir0_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_28
       (.I0(\eir_fl_reg[15] [4]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[4]),
        .I4(fadr_1_fl),
        .I5(fdatx[4]),
        .O(ir0_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_29
       (.I0(\eir_fl_reg[15] [3]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[3]),
        .I4(fadr_1_fl),
        .I5(fdatx[3]),
        .O(ir0_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_3
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_19_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [13]),
        .O(in0[13]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_30
       (.I0(\eir_fl_reg[15] [2]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[2]),
        .I4(fadr_1_fl),
        .I5(fdatx[2]),
        .O(ir0_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_31
       (.I0(\eir_fl_reg[15] [1]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[1]),
        .I4(fadr_1_fl),
        .I5(fdatx[1]),
        .O(ir0_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_32
       (.I0(\eir_fl_reg[15] [0]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[0]),
        .I4(fadr_1_fl),
        .I5(fdatx[0]),
        .O(ir0_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_4
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_20_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [12]),
        .O(in0[12]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_5
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_21_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [11]),
        .O(in0[11]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_6
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_22_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [10]),
        .O(in0[10]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_7
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_23_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [9]),
        .O(in0[9]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_8
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_24_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [8]),
        .O(in0[8]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_9
       (.I0(rst_n_fl),
        .I1(ir0_inferred_i_25_n_0),
        .I2(fch_term_fl),
        .I3(\ir0_fl_reg[0] ),
        .I4(ctl_fetch0_fl),
        .I5(\ir0_fl_reg[15] [7]),
        .O(in0[7]));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[20]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [0]),
        .I2(fch_term_fl),
        .I3(\ir1_id_fl[20]_i_2_n_0 ),
        .I4(\ir0_fl_reg[0] ),
        .I5(out),
        .O(fch_wrbufn1));
  LUT5 #(
    .INIT(32'hCACCFAFF)) 
    \ir1_id_fl[20]_i_2 
       (.I0(\ir1_id_fl_reg[20] ),
        .I1(fadr_1_fl),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\ir1_id_fl_reg[21]_0 [4]),
        .O(\ir1_id_fl[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[21]_i_1 
       (.I0(rst_n_fl),
        .I1(\ir1_id_fl_reg[21] [1]),
        .I2(fch_term_fl),
        .I3(\ir1_id_fl[21]_i_2_n_0 ),
        .I4(\ir0_fl_reg[0] ),
        .I5(out),
        .O(fch_memacc1));
  LUT5 #(
    .INIT(32'hDDDDF0DD)) 
    \ir1_id_fl[21]_i_2 
       (.I0(\ir1_id_fl_reg[21]_0 [5]),
        .I1(fadr_1_fl),
        .I2(\ir1_id_fl_reg[21]_1 ),
        .I3(stat[1]),
        .I4(stat[0]),
        .O(\ir1_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_1
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_18_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [15]),
        .O(ir1[15]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_10
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_27_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [6]),
        .O(ir1[6]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_11
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_28_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [5]),
        .O(ir1[5]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_12
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_29_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [4]),
        .O(ir1[4]));
  LUT6 #(
    .INIT(64'h808080AA80808080)) 
    ir1_inferred_i_13
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_30_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [3]),
        .O(ir1[3]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_31_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl),
        .I4(\ir1_fl_reg[15] [2]),
        .O(ir1[2]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir1_inferred_i_32_n_0),
        .I2(ctl_fetch1_fl),
        .I3(fch_term_fl),
        .I4(\ir1_fl_reg[15] [1]),
        .O(ir1[1]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_33_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [0]),
        .O(ir1[0]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_18
       (.I0(fdatx[15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[15]),
        .O(ir1_inferred_i_18_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_19
       (.I0(fdatx[14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[14]),
        .O(ir1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_2
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_19_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [14]),
        .O(ir1[14]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_20
       (.I0(fdatx[13]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[13]),
        .O(ir1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_21
       (.I0(fdatx[12]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[12]),
        .O(ir1_inferred_i_21_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_22
       (.I0(fdatx[11]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[11]),
        .O(ir1_inferred_i_22_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_23
       (.I0(fdatx[10]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[10]),
        .O(ir1_inferred_i_23_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_24
       (.I0(fdatx[9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[9]),
        .O(ir1_inferred_i_24_n_0));
  LUT5 #(
    .INIT(32'hF355F3F3)) 
    ir1_inferred_i_25
       (.I0(fdatx[8]),
        .I1(fdat[8]),
        .I2(fadr_1_fl),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(ir1_inferred_i_25_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_26
       (.I0(fdatx[7]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[7]),
        .O(ir1_inferred_i_26_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_27
       (.I0(fdatx[6]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[6]),
        .O(ir1_inferred_i_27_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_28
       (.I0(fdatx[5]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[5]),
        .O(ir1_inferred_i_28_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_29
       (.I0(fdatx[4]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fadr_1_fl),
        .I4(fdat[4]),
        .O(ir1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_3
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_20_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [13]),
        .O(ir1[13]));
  LUT5 #(
    .INIT(32'h0808FB08)) 
    ir1_inferred_i_30
       (.I0(fdatx[3]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(fdat[3]),
        .I4(fadr_1_fl),
        .O(ir1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h4C4440440C000000)) 
    ir1_inferred_i_31
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(fdatx[2]),
        .I5(fdat[2]),
        .O(ir1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h40CC404040004040)) 
    ir1_inferred_i_32
       (.I0(fadr_1_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(fdat[1]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(fdatx[1]),
        .O(ir1_inferred_i_32_n_0));
  LUT5 #(
    .INIT(32'hF355F3F3)) 
    ir1_inferred_i_33
       (.I0(fdatx[0]),
        .I1(fdat[0]),
        .I2(fadr_1_fl),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(ir1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_4
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_21_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [12]),
        .O(ir1[12]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_5
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_22_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [11]),
        .O(ir1[11]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_6
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_23_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [10]),
        .O(ir1[10]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_7
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_24_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [9]),
        .O(ir1[9]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_8
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_25_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [8]),
        .O(ir1[8]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_9
       (.I0(rst_n_fl),
        .I1(\ir1_fl_reg[0] ),
        .I2(ir1_inferred_i_26_n_0),
        .I3(ctl_fetch1_fl),
        .I4(fch_term_fl),
        .I5(\ir1_fl_reg[15] [7]),
        .O(ir1[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [0]),
        .O(\iv_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [10]),
        .O(\iv_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [11]),
        .O(\iv_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [12]),
        .O(\iv_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [13]),
        .O(\iv_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [14]),
        .O(\iv_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [15]),
        .O(\iv_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0008)) 
    \iv[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_3 
       (.I0(\grn[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\sr[15]_i_4_n_0 ),
        .O(\rgf/c0bus_sel_cr [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [1]),
        .O(\iv_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [2]),
        .O(\iv_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [3]),
        .O(\iv_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [4]),
        .O(\iv_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [5]),
        .O(\iv_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [6]),
        .O(\iv_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [7]),
        .O(\iv_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [8]),
        .O(\iv_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\iv_reg[15]_0 [9]),
        .O(\iv_reg[15] [9]));
  LUT6 #(
    .INIT(64'h00EB00EB000000FB)) 
    \nir_id[24]_i_1 
       (.I0(stat[2]),
        .I1(fch_issu1_ir),
        .I2(stat[1]),
        .I3(\nir_id[24]_i_3_n_0 ),
        .I4(\nir_id[24]_i_4_n_0 ),
        .I5(brdy_0),
        .O(E));
  LUT5 #(
    .INIT(32'hFFFFBEEE)) 
    \nir_id[24]_i_3 
       (.I0(\stat[1]_i_4_n_0 ),
        .I1(stat[0]),
        .I2(stat[2]),
        .I3(stat[1]),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\nir_id[24]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_4 
       (.I0(stat[0]),
        .I1(\stat_reg[2]_0 ),
        .O(\nir_id[24]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    \pc0[0]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(fch_irq_req),
        .I2(p_2_in_0[0]),
        .I3(\stat_reg[1]_0 ),
        .I4(\pc0_reg[12] [0]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[10]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [10]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[10]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [1]),
        .O(D[10]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[11]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [11]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[11]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [2]),
        .O(D[11]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[12]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [12]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[12]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [3]),
        .O(D[12]));
  LUT4 #(
    .INIT(16'hFBFA)) 
    \pc0[15]_i_3 
       (.I0(\fadr[15]_INST_0_i_6_n_0 ),
        .I1(stat[1]),
        .I2(\fadr[15]_INST_0_i_5_n_0 ),
        .I3(stat[0]),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hF0E2F0E2FFE200E2)) 
    \pc0[1]_i_1 
       (.I0(O[0]),
        .I1(\stat_reg[1]_0 ),
        .I2(p_2_in_0[1]),
        .I3(fch_irq_req),
        .I4(\pc0_reg[12] [1]),
        .I5(\pc0_reg[3] ),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[2]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [2]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[2]),
        .I4(\stat_reg[1]_0 ),
        .I5(O[1]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[3]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [3]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[3]),
        .I4(\stat_reg[1]_0 ),
        .I5(O[2]),
        .O(D[3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[4]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [4]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[4]),
        .I4(\stat_reg[1]_0 ),
        .I5(O[3]),
        .O(D[4]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[5]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [5]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[5]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [0]),
        .O(D[5]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[6]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [6]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[6]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [1]),
        .O(D[6]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[7]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [7]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[7]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [2]),
        .O(D[7]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[8]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [8]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[8]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [3]),
        .O(D[8]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[9]_i_1 
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [9]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[9]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [0]),
        .O(D[9]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_1
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [7]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[7]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [2]),
        .O(\pc_reg[7] [3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_2
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [6]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[6]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [1]),
        .O(\pc_reg[7] [2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_3
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [5]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[5]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [0]),
        .O(\pc_reg[7] [1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_4
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [4]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[4]),
        .I4(\stat_reg[1]_0 ),
        .I5(O[3]),
        .O(\pc_reg[7] [0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_1
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [11]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[11]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [2]),
        .O(\pc_reg[11] [3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_2
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [10]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[10]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [1]),
        .O(\pc_reg[11] [2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_3
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [9]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[9]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [0]),
        .O(\pc_reg[11] [1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_4
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [8]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[8]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[8] [3]),
        .O(\pc_reg[11] [0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_4
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [12]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[12]),
        .I4(\stat_reg[1]_0 ),
        .I5(\fadr[12] [3]),
        .O(\pc_reg[12] ));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry_i_1
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [3]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[3]),
        .I4(\stat_reg[1]_0 ),
        .I5(O[2]),
        .O(S[3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry_i_2
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [2]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[2]),
        .I4(\stat_reg[1]_0 ),
        .I5(O[1]),
        .O(S[2]));
  LUT6 #(
    .INIT(64'h10BF10B010BF1FBF)) 
    pc10_carry_i_3
       (.I0(\pc0_reg[3] ),
        .I1(\pc0_reg[12] [1]),
        .I2(fch_irq_req),
        .I3(p_2_in_0[1]),
        .I4(\stat_reg[1]_0 ),
        .I5(O[0]),
        .O(S[1]));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    pc10_carry_i_4
       (.I0(\pc0_reg[3] ),
        .I1(fch_irq_req),
        .I2(p_2_in_0[0]),
        .I3(\stat_reg[1]_0 ),
        .I4(\pc0_reg[12] [0]),
        .O(S[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[0]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[0]));
  LUT6 #(
    .INIT(64'hF4F7FFFFB0800000)) 
    \pc[0]_i_2 
       (.I0(\pc0_reg[3] ),
        .I1(fch_irq_req),
        .I2(p_2_in_0[0]),
        .I3(\stat_reg[1]_0 ),
        .I4(\pc_reg[0] ),
        .I5(\pc0_reg[12] [0]),
        .O(\pc[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[10]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[10]_i_2 
       (.I0(D[10]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [10]),
        .O(\pc[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[11]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[11]_i_2 
       (.I0(D[11]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [11]),
        .O(\pc[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[12]_i_4_n_0 ),
        .O(rgf_selc1_stat_reg[12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [12]),
        .I3(rgf_selc1_stat),
        .I4(Q[12]),
        .O(\rgf/rgf_c1bus_0 [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [11]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [12]),
        .O(\rgf/rgf_c0bus_0 [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[12]_i_4 
       (.I0(D[12]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [12]),
        .O(\pc[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[13] ),
        .O(rgf_selc1_stat_reg[13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [13]),
        .I3(rgf_selc1_stat),
        .I4(Q[13]),
        .O(\rgf/rgf_c1bus_0 [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [12]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [13]),
        .O(\rgf/rgf_c0bus_0 [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[14]_1 ),
        .O(rgf_selc1_stat_reg[14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [14]),
        .I3(rgf_selc1_stat),
        .I4(Q[14]),
        .O(\rgf/rgf_c1bus_0 [14]));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \pc[14]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[14] ),
        .I3(\pc_reg[14]_0 ),
        .I4(rgf_selc0_stat),
        .I5(\pc_reg[15]_1 [14]),
        .O(\rgf/rgf_c0bus_0 [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc_reg[15]_2 ),
        .O(rgf_selc1_stat_reg[15]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [15]),
        .I3(rgf_selc1_stat),
        .I4(Q[15]),
        .O(\rgf/rgf_c1bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [13]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [15]),
        .O(\rgf/rgf_c0bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_5 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\sr[15]_i_4_n_0 ),
        .O(\rgf/c0bus_sel_cr [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[1]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[1]_i_2 
       (.I0(D[1]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [1]),
        .O(\pc[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[2]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[2]_i_2 
       (.I0(D[2]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [2]),
        .O(\pc[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[3]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[3]_i_2 
       (.I0(D[3]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [3]),
        .O(\pc[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[4]_i_4_n_0 ),
        .O(rgf_selc1_stat_reg[4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [4]),
        .I3(rgf_selc1_stat),
        .I4(Q[4]),
        .O(\rgf/rgf_c1bus_0 [4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [3]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [4]),
        .O(\rgf/rgf_c0bus_0 [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[4]_i_4 
       (.I0(D[4]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [4]),
        .O(\pc[4]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[5]_i_3_n_0 ),
        .O(rgf_selc1_stat_reg[5]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[5]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [5]),
        .I3(rgf_selc1_stat),
        .I4(Q[5]),
        .O(\rgf/rgf_c1bus_0 [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[5]_i_3 
       (.I0(D[5]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [5]),
        .O(\pc[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[6]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[6]_i_2 
       (.I0(D[6]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [6]),
        .O(\pc[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[7]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[7]_i_2 
       (.I0(D[7]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [7]),
        .O(\pc[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[8]_i_4_n_0 ),
        .O(rgf_selc1_stat_reg[8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_2 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [8]),
        .I3(rgf_selc1_stat),
        .I4(Q[8]),
        .O(\rgf/rgf_c1bus_0 [8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [7]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [8]),
        .O(\rgf/rgf_c0bus_0 [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[8]_i_4 
       (.I0(D[8]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [8]),
        .O(\pc[8]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[9]_i_2_n_0 ),
        .O(rgf_selc1_stat_reg[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[9]_i_2 
       (.I0(D[9]),
        .I1(\pc_reg[0] ),
        .I2(\pc0_reg[12] [9]),
        .O(\pc[9]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc0_stat_i_3
       (.I0(fch_wrbufn0),
        .O(p_2_in));
  LUT5 #(
    .INIT(32'hFFFF8880)) 
    rgf_selc0_stat_i_4
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(rst_n_fl),
        .I2(fch_term_fl),
        .I3(\ir0_id_fl_reg[21] [0]),
        .I4(\ir0_fl_reg[0] ),
        .O(fch_wrbufn0));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc1_stat_i_2
       (.I0(fch_wrbufn1),
        .O(rst_n_fl_reg));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[0]_i_1 
       (.I0(\sp_reg[0] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [0]),
        .I4(\rgf/rgf_c1bus_0 [0]),
        .O(\sp_reg[15] [0]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[10]_i_1 
       (.I0(\sp_reg[10] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [10]),
        .I4(\rgf/rgf_c1bus_0 [10]),
        .O(\sp_reg[15] [10]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[11]_i_1 
       (.I0(\sp_reg[11] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [11]),
        .I4(\rgf/rgf_c1bus_0 [11]),
        .O(\sp_reg[15] [11]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[12]_i_1 
       (.I0(\sp_reg[12] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [12]),
        .I4(\rgf/rgf_c1bus_0 [12]),
        .O(\sp_reg[15] [12]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[13]_i_1 
       (.I0(\sp_reg[13] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [13]),
        .I4(\rgf/rgf_c1bus_0 [13]),
        .O(\sp_reg[15] [13]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[14]_i_1 
       (.I0(\sp_reg[14] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [14]),
        .I4(\rgf/rgf_c1bus_0 [14]),
        .O(\sp_reg[15] [14]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[15]_i_1 
       (.I0(\sp_reg[15]_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [15]),
        .I4(\rgf/rgf_c1bus_0 [15]),
        .O(\sp_reg[15] [15]));
  LUT3 #(
    .INIT(8'h04)) 
    \sp[15]_i_3 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\sr[15]_i_4_n_0 ),
        .O(\rgf/c0bus_sel_cr [2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [2]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[1]_i_1 
       (.I0(\sp_reg[1] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [1]),
        .I4(\rgf/rgf_c1bus_0 [1]),
        .O(\sp_reg[15] [1]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[2]_i_1 
       (.I0(\sp_reg[2] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .O(\sp_reg[15] [2]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[3]_i_1 
       (.I0(\sp_reg[3] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\rgf/rgf_c1bus_0 [3]),
        .O(\sp_reg[15] [3]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[4]_i_1 
       (.I0(\sp_reg[4] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [4]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .O(\sp_reg[15] [4]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[5]_i_1 
       (.I0(\sp_reg[5] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [5]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .O(\sp_reg[15] [5]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[6]_i_1 
       (.I0(\sp_reg[6] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [6]),
        .I4(\rgf/rgf_c1bus_0 [6]),
        .O(\sp_reg[15] [6]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[7]_i_1 
       (.I0(\sp_reg[7] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [7]),
        .I4(\rgf/rgf_c1bus_0 [7]),
        .O(\sp_reg[15] [7]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[8]_i_1 
       (.I0(\sp_reg[8] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [8]),
        .I4(\rgf/rgf_c1bus_0 [8]),
        .O(\sp_reg[15] [8]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[9]_i_1 
       (.I0(\sp_reg[9] ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [9]),
        .I4(\rgf/rgf_c1bus_0 [9]),
        .O(\sp_reg[15] [9]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[0]_i_1 
       (.I0(\sr_reg[15]_0 [0]),
        .I1(\sr[15]_i_2_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\sr[11]_i_2_n_0 ),
        .I4(\rgf/rgf_c1bus_0 [0]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [0]),
        .O(\rgf/rgf_c0bus_0 [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [0]),
        .I3(rgf_selc1_stat),
        .I4(Q[0]),
        .O(\rgf/rgf_c1bus_0 [0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[10]_i_1 
       (.I0(\sr_reg[15]_0 [10]),
        .I1(\sr[15]_i_2_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\sr[11]_i_2_n_0 ),
        .I4(\rgf/rgf_c1bus_0 [10]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [9]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [10]),
        .O(\rgf/rgf_c0bus_0 [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [10]),
        .I3(rgf_selc1_stat),
        .I4(Q[10]),
        .O(\rgf/rgf_c1bus_0 [10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[11]_i_1 
       (.I0(\sr_reg[15]_0 [11]),
        .I1(\sr[15]_i_2_n_0 ),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c0bus_0 [11]),
        .I4(\rgf/rgf_c1bus_0 [11]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_10 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[13]_i_5_2 [0]),
        .I3(rgf_selc1_stat),
        .I4(\sr[13]_i_5_3 [0]),
        .O(\rgf/rctl/rgf_selc1 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \sr[11]_i_2 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\sr[15]_i_4_n_0 ),
        .I3(\sr[13]_i_2_n_0 ),
        .O(\sr[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [10]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [11]),
        .O(\rgf/rgf_c0bus_0 [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_4 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [11]),
        .I3(rgf_selc1_stat),
        .I4(Q[11]),
        .O(\rgf/rgf_c1bus_0 [11]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \sr[11]_i_5 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(rst_n),
        .O(\sr[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_6 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[13]_i_5_0 [2]),
        .I3(rgf_selc1_stat),
        .I4(\sr[13]_i_5_1 [2]),
        .O(\rgf/rctl/rgf_selc1_rn [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_7 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[13]_i_5_0 [0]),
        .I3(rgf_selc1_stat),
        .I4(\sr[13]_i_5_1 [0]),
        .O(\rgf/rctl/rgf_selc1_rn [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_8 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\sr[13]_i_5_0 [1]),
        .I3(rgf_selc1_stat),
        .I4(\sr[13]_i_5_1 [1]),
        .O(\rgf/rctl/rgf_selc1_rn [1]));
  LUT6 #(
    .INIT(64'hAAFFAAFFBABFFFFF)) 
    \sr[11]_i_9 
       (.I0(\rgf/rctl/rgf_selc1 ),
        .I1(\sr[13]_i_5_3 [1]),
        .I2(rgf_selc1_stat),
        .I3(\sr[13]_i_5_2 [1]),
        .I4(\grn_reg[15] ),
        .I5(fch_wrbufn1),
        .O(\sr[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFEFEFF000000)) 
    \sr[12]_i_1 
       (.I0(\sr[13]_i_2_n_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\sr[13]_i_4_n_0 ),
        .I3(\sr_reg[15]_0 [12]),
        .I4(\sr[15]_i_2_n_0 ),
        .I5(cpuid[0]),
        .O(\sr_reg[15] [12]));
  LUT6 #(
    .INIT(64'hFFFEFEFEFF000000)) 
    \sr[13]_i_1 
       (.I0(\sr[13]_i_2_n_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\sr[13]_i_4_n_0 ),
        .I3(\sr_reg[15]_0 [13]),
        .I4(\sr[15]_i_2_n_0 ),
        .I5(cpuid[1]),
        .O(\sr_reg[15] [13]));
  LUT5 #(
    .INIT(32'h0008005D)) 
    \sr[13]_i_10 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\sr[15]_i_4_n_0 ),
        .I4(\sr[15]_i_3_n_0 ),
        .O(\sr[13]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[13]_i_2 
       (.I0(\sr[13]_i_5_n_0 ),
        .I1(ctl_sr_ldie1),
        .O(\sr[13]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[13]_i_4 
       (.I0(ctl_sr_upd0),
        .I1(\sr[13]_i_10_n_0 ),
        .O(\sr[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF555555D7)) 
    \sr[13]_i_5 
       (.I0(rst_n),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\sr[11]_i_9_n_0 ),
        .I5(ctl_sr_upd1),
        .O(\sr[13]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[14]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [14]),
        .O(\sr_reg[15] [14]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[15]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [15]),
        .O(\sr_reg[15] [15]));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \sr[15]_i_2 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\sr[15]_i_4_n_0 ),
        .I3(ctl_sr_ldie1),
        .I4(\sr[15]_i_6_n_0 ),
        .I5(\sr[15]_i_7_n_0 ),
        .O(\sr[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .O(\sr[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hE4E0A0E0FFFFFFFF)) 
    \sr[15]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\grn[15]_i_3__5_0 [0]),
        .I3(rgf_selc0_stat),
        .I4(\grn[15]_i_3__5_1 [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\sr[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hABAAAAAA)) 
    \sr[15]_i_6 
       (.I0(ctl_sr_upd1),
        .I1(\sr[11]_i_9_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\sr[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    \sr[15]_i_7 
       (.I0(\sr[11]_i_9_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(rst_n),
        .O(\sr[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[1]_i_1 
       (.I0(\sr_reg[15]_0 [1]),
        .I1(\sr[15]_i_2_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\sr[11]_i_2_n_0 ),
        .I4(\rgf/rgf_c1bus_0 [1]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [1]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [1]),
        .O(\rgf/rgf_c0bus_0 [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [1]),
        .I3(rgf_selc1_stat),
        .I4(Q[1]),
        .O(\rgf/rgf_c1bus_0 [1]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[2]_i_1 
       (.I0(\sr[2]_i_2_n_0 ),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\sr[11]_i_5_n_0 ),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .O(\sr_reg[15] [2]));
  LUT6 #(
    .INIT(64'h08080808FF080808)) 
    \sr[2]_i_2 
       (.I0(\sr[3]_i_5_n_0 ),
        .I1(\sr_reg[15]_0 [2]),
        .I2(\sr[15]_i_7_n_0 ),
        .I3(\sr[3]_i_6_n_0 ),
        .I4(fch_irq_lev[0]),
        .I5(\sr[13]_i_5_n_0 ),
        .O(\sr[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [2]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [2]),
        .O(\rgf/rgf_c0bus_0 [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_4 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [2]),
        .I3(rgf_selc1_stat),
        .I4(Q[2]),
        .O(\rgf/rgf_c1bus_0 [2]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[3]_i_1 
       (.I0(\sr[3]_i_2_n_0 ),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\sr[11]_i_5_n_0 ),
        .I4(\rgf/rgf_c1bus_0 [3]),
        .O(\sr_reg[15] [3]));
  LUT6 #(
    .INIT(64'h08080808FF080808)) 
    \sr[3]_i_2 
       (.I0(\sr[3]_i_5_n_0 ),
        .I1(\sr_reg[15]_0 [3]),
        .I2(\sr[15]_i_7_n_0 ),
        .I3(\sr[3]_i_6_n_0 ),
        .I4(fch_irq_lev[1]),
        .I5(\sr[13]_i_5_n_0 ),
        .O(\sr[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \sr[3]_i_3 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\sr_reg[3] ),
        .I3(\sr_reg[3]_0 ),
        .I4(rgf_selc0_stat),
        .I5(\pc_reg[15]_1 [3]),
        .O(\rgf/rgf_c0bus_0 [3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[3]_i_4 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [3]),
        .I3(rgf_selc1_stat),
        .I4(Q[3]),
        .O(\rgf/rgf_c1bus_0 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FE00)) 
    \sr[3]_i_5 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\sr[15]_i_4_n_0 ),
        .I3(\sr[3]_i_8_n_0 ),
        .I4(ctl_sr_ldie1),
        .I5(\sr[15]_i_6_n_0 ),
        .O(\sr[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF00FE)) 
    \sr[3]_i_6 
       (.I0(\sr[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\sr[15]_i_4_n_0 ),
        .I3(\sr[3]_i_8_n_0 ),
        .I4(ctl_sr_ldie1),
        .O(\sr[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0008FFFFFFFF)) 
    \sr[3]_i_8 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\sr[15]_i_4_n_0 ),
        .I4(ctl_sr_upd0),
        .I5(ctl_sr_ldie0),
        .O(\sr[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \sr[4]_i_1 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(alu_sr_flag1),
        .I2(\sr[4]_i_4_n_0 ),
        .I3(\sr_reg[4] ),
        .I4(alu_sr_flag0[0]),
        .I5(\sr[4]_i_7_n_0 ),
        .O(\sr_reg[15] [4]));
  LUT6 #(
    .INIT(64'h0000FFF700000000)) 
    \sr[4]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(\sr[15]_i_7_n_0 ),
        .I5(ctl_sr_upd1),
        .O(\sr[4]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[4]_i_4 
       (.I0(\sr[7]_i_4_n_0 ),
        .I1(\rgf/rgf_c1bus_0 [4]),
        .I2(\sr[7]_i_6_n_0 ),
        .I3(\rgf/rgf_c0bus_0 [4]),
        .O(\sr[4]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[4]_i_7 
       (.I0(\sr[13]_i_10_n_0 ),
        .I1(ctl_sr_upd0),
        .I2(ctl_sr_ldie1),
        .I3(\sr[13]_i_5_n_0 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \sr[5]_i_1 
       (.I0(\sr[5]_i_2_n_0 ),
        .I1(\sr[5]_i_3_n_0 ),
        .I2(\sr[7]_i_6_n_0 ),
        .I3(\rgf/rgf_c0bus_0 [5]),
        .I4(\sr_reg[5] ),
        .I5(\sr[5]_i_6_n_0 ),
        .O(\sr_reg[15] [5]));
  LUT6 #(
    .INIT(64'hAAAAAAAA00008828)) 
    \sr[5]_i_2 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr_reg[5]_0 ),
        .I2(\sr_reg[5]_1 ),
        .I3(\sr_reg[5]_2 ),
        .I4(\sr_reg[5]_3 ),
        .I5(\sr_reg[5]_4 ),
        .O(\sr[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0B80000000000)) 
    \sr[5]_i_3 
       (.I0(Q[5]),
        .I1(rgf_selc1_stat),
        .I2(\pc_reg[15] [5]),
        .I3(\grn_reg[15] ),
        .I4(fch_wrbufn1),
        .I5(\sr[7]_i_4_n_0 ),
        .O(\sr[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[5]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [4]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [5]),
        .O(\rgf/rgf_c0bus_0 [5]));
  LUT6 #(
    .INIT(64'hFFFF600000000000)) 
    \sr[5]_i_6 
       (.I0(\sr_reg[5]_5 ),
        .I1(\sr_reg[5]_6 ),
        .I2(\sr_reg[5]_7 ),
        .I3(\sr_reg[5]_8 ),
        .I4(\sr_reg[5]_9 ),
        .I5(\sr[4]_i_7_n_0 ),
        .O(\sr[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \sr[6]_i_1 
       (.I0(\sr[6]_i_2_n_0 ),
        .I1(\sr[7]_i_4_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\sr[7]_i_6_n_0 ),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\sr[6]_i_5_n_0 ),
        .O(\sr_reg[15] [6]));
  LUT5 #(
    .INIT(32'hAAAA0028)) 
    \sr[6]_i_2 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr_reg[6] ),
        .I2(\sr_reg[6]_0 ),
        .I3(\sr_reg[7] ),
        .I4(\sr_reg[5]_0 ),
        .O(\sr[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[6]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [6]),
        .I3(rgf_selc1_stat),
        .I4(Q[6]),
        .O(\rgf/rgf_c1bus_0 [6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[6]_i_4 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [5]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [6]),
        .O(\rgf/rgf_c0bus_0 [6]));
  LUT5 #(
    .INIT(32'hFFA8A8A8)) 
    \sr[6]_i_5 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(\sr_reg[5]_5 ),
        .I2(\sr_reg[6]_1 ),
        .I3(rst_n_0),
        .I4(\sr_reg[15]_0 [6]),
        .O(\sr[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \sr[7]_i_1 
       (.I0(\sr[7]_i_2_n_0 ),
        .I1(\rgf/rgf_c1bus_0 [7]),
        .I2(\sr[7]_i_4_n_0 ),
        .I3(\rgf/rgf_c0bus_0 [7]),
        .I4(\sr[7]_i_6_n_0 ),
        .I5(\sr[7]_i_7_n_0 ),
        .O(\sr_reg[15] [7]));
  LUT6 #(
    .INIT(64'hF4F4FFF400000000)) 
    \sr[7]_i_2 
       (.I0(\sr_reg[5]_2 ),
        .I1(\sr_reg[5]_1 ),
        .I2(\sr_reg[7]_0 ),
        .I3(\sr_reg[7]_1 ),
        .I4(\sr_reg[7] ),
        .I5(\sr[4]_i_2_n_0 ),
        .O(\sr[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[7]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [7]),
        .I3(rgf_selc1_stat),
        .I4(Q[7]),
        .O(\rgf/rgf_c1bus_0 [7]));
  LUT5 #(
    .INIT(32'h00210000)) 
    \sr[7]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(rst_n),
        .O(\sr[7]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[7]_i_5 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [6]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [7]),
        .O(\rgf/rgf_c0bus_0 [7]));
  LUT3 #(
    .INIT(8'h02)) 
    \sr[7]_i_6 
       (.I0(\sr[13]_i_10_n_0 ),
        .I1(ctl_sr_ldie1),
        .I2(\sr[13]_i_5_n_0 ),
        .O(\sr[7]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[7]_i_7 
       (.I0(alu_sr_flag0[1]),
        .I1(\sr[4]_i_7_n_0 ),
        .I2(\sr_reg[15]_0 [7]),
        .I3(rst_n_0),
        .O(\sr[7]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h31)) 
    \sr[7]_i_9 
       (.I0(\sr[13]_i_4_n_0 ),
        .I1(\sr[13]_i_5_n_0 ),
        .I2(ctl_sr_ldie1),
        .O(rst_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[8]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\sr_reg[15]_0 [8]),
        .O(\sr_reg[15] [8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[9]_i_1 
       (.I0(\sr_reg[15]_0 [9]),
        .I1(\sr[15]_i_2_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\sr[11]_i_2_n_0 ),
        .I4(\rgf/rgf_c1bus_0 [9]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\sr_reg[15] [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_2 
       (.I0(fch_wrbufn0),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15]_0 [8]),
        .I3(rgf_selc0_stat),
        .I4(\pc_reg[15]_1 [9]),
        .O(\rgf/rgf_c0bus_0 [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_3 
       (.I0(fch_wrbufn1),
        .I1(\grn_reg[15] ),
        .I2(\pc_reg[15] [9]),
        .I3(rgf_selc1_stat),
        .I4(Q[9]),
        .O(\rgf/rgf_c1bus_0 [9]));
  LUT5 #(
    .INIT(32'hE0F5E0A0)) 
    \stat[0]_i_1__0 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\stat[0]_i_2__2_n_0 ),
        .I3(brdy_0),
        .I4(\stat[0]_i_3_n_0 ),
        .O(stat_nx[0]));
  LUT6 #(
    .INIT(64'h000B0000FFFFFFFF)) 
    \stat[0]_i_1__1 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[0]_5 ),
        .I2(\stat_reg[0]_6 ),
        .I3(\stat_reg[0]_7 ),
        .I4(\stat[0]_i_6__0_n_0 ),
        .I5(\stat_reg[0]_3 ),
        .O(\stat_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hAA2A)) 
    \stat[0]_i_2__2 
       (.I0(\pc0_reg[12] [1]),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(stat[2]),
        .O(\stat[0]_i_2__2_n_0 ));
  LUT4 #(
    .INIT(16'h8808)) 
    \stat[0]_i_3 
       (.I0(\fadr[15]_INST_0_i_4_n_0 ),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(stat[2]),
        .O(\stat[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE0FFE0E0)) 
    \stat[0]_i_6__0 
       (.I0(\ir0_fl_reg[0] ),
        .I1(rst_n_fl_reg_3[1]),
        .I2(fch_memacc1),
        .I3(\stat_reg[0]_8 [0]),
        .I4(\stat_reg[0]_8 [1]),
        .O(\stat[0]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000088888A88)) 
    \stat[1]_i_1 
       (.I0(\stat[1]_i_2_n_0 ),
        .I1(\stat[1]_i_3__1_n_0 ),
        .I2(\stat[1]_i_4_n_0 ),
        .I3(stat[1]),
        .I4(stat[0]),
        .I5(\fadr[15]_INST_0_i_5_n_0 ),
        .O(stat_nx[1]));
  LUT6 #(
    .INIT(64'h7F733F333333737F)) 
    \stat[1]_i_2 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat[1]_i_3__1_n_0 ),
        .I2(brdy_0),
        .I3(\fadr[15]_INST_0_i_4_n_0 ),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(\stat[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hCDCCCDDD)) 
    \stat[1]_i_3__1 
       (.I0(stat[0]),
        .I1(stat[2]),
        .I2(out),
        .I3(fch_term_fl),
        .I4(fch_issu1_fl),
        .O(\stat[1]_i_3__1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[1]_i_4 
       (.I0(brdy_0),
        .I1(\stat_reg[0]_2 ),
        .O(\stat[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h01555555)) 
    \stat[2]_i_18 
       (.I0(\ir0_fl_reg[0] ),
        .I1(\ir0_id_fl_reg[21] [1]),
        .I2(fch_term_fl),
        .I3(rst_n_fl),
        .I4(\ir0_id_fl[21]_i_2_n_0 ),
        .O(fch_irq_req_fl_reg));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1__1 
       (.I0(rst_n_fl),
        .O(\stat[2]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA000002AAAA)) 
    \stat[2]_i_2 
       (.I0(\stat[2]_i_3_n_0 ),
        .I1(fch_issu1_ir),
        .I2(stat[1]),
        .I3(stat[2]),
        .I4(stat[0]),
        .I5(\stat_reg[2]_0 ),
        .O(stat_nx[2]));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_3 
       (.I0(brdy_0),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\stat[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5555515555555555)) 
    \stat[2]_i_4 
       (.I0(ctl_fetch_ext0),
        .I1(fch_leir_nir_reg_0),
        .I2(ctl_fetch1_fl_i_21_0[2]),
        .I3(fch_leir_nir_reg_1),
        .I4(\stat[2]_i_6__1_n_0 ),
        .I5(rst_n_fl_reg_0),
        .O(\stat_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFFFF)) 
    \stat[2]_i_6__1 
       (.I0(ctl_fetch1_fl_i_21_0[12]),
        .I1(ctl_fetch1_fl_i_21_0[11]),
        .I2(ctl_fetch1_fl_i_21_0[13]),
        .I3(ctl_fetch1_fl_reg[2]),
        .I4(ctl_fetch1_fl_i_21_0[0]),
        .I5(ctl_fetch1_fl_i_21_0[1]),
        .O(\stat[2]_i_6__1_n_0 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[0]),
        .Q(stat[0]),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[1]),
        .Q(stat[1]),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx[2]),
        .Q(stat[2]),
        .R(\stat[2]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [0]),
        .O(\tr_reg[15] [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [10]),
        .O(\tr_reg[15] [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [11]),
        .O(\tr_reg[15] [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [12]),
        .O(\tr_reg[15] [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [13]),
        .O(\tr_reg[15] [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [14]),
        .O(\tr_reg[15] [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [15]),
        .O(\tr_reg[15] [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [4]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\sr[15]_i_4_n_0 ),
        .O(\rgf/c0bus_sel_cr [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [1]),
        .O(\tr_reg[15] [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [2]),
        .O(\tr_reg[15] [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [3]),
        .O(\tr_reg[15] [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [4]),
        .O(\tr_reg[15] [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [5]),
        .O(\tr_reg[15] [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [6]),
        .O(\tr_reg[15] [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [7]),
        .O(\tr_reg[15] [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [8]),
        .O(\tr_reg[15] [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\tr_reg[15]_0 [9]),
        .O(\tr_reg[15] [9]));
endmodule

module mcss_fsm
   (\stat_reg[2]_0 ,
    \stat_reg[1]_0 ,
    Q,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    \stat_reg[0]_2 ,
    \stat_reg[0]_3 ,
    \stat_reg[1]_1 ,
    \stat_reg[0]_4 ,
    \stat_reg[1]_2 ,
    \stat_reg[2]_1 ,
    \stat_reg[1]_3 ,
    \stat_reg[1]_4 ,
    \stat_reg[0]_5 ,
    \stat_reg[0]_6 ,
    \stat_reg[0]_7 ,
    \stat_reg[0]_8 ,
    \stat_reg[2]_2 ,
    \stat_reg[2]_3 ,
    \stat_reg[0]_9 ,
    \stat_reg[0]_10 ,
    \stat_reg[0]_11 ,
    \stat_reg[0]_12 ,
    \stat_reg[1]_5 ,
    \stat_reg[1]_6 ,
    \stat_reg[2]_4 ,
    \stat_reg[0]_13 ,
    \stat_reg[0]_14 ,
    \stat_reg[0]_15 ,
    out,
    \stat_reg[1]_7 ,
    \stat_reg[1]_8 ,
    \ccmd[4]_INST_0_i_2 ,
    brdy,
    ctl_bcc_take1_fl,
    ctl_bcc_take0_fl,
    \stat_reg[0]_16 ,
    rgf_sr_dr,
    crdy,
    SR,
    D,
    clk);
  output \stat_reg[2]_0 ;
  output \stat_reg[1]_0 ;
  output [2:0]Q;
  output \stat_reg[0]_0 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[0]_4 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[2]_1 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[1]_4 ;
  output \stat_reg[0]_5 ;
  output \stat_reg[0]_6 ;
  output \stat_reg[0]_7 ;
  output \stat_reg[0]_8 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[2]_3 ;
  output \stat_reg[0]_9 ;
  output \stat_reg[0]_10 ;
  output \stat_reg[0]_11 ;
  output \stat_reg[0]_12 ;
  output \stat_reg[1]_5 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[2]_4 ;
  output \stat_reg[0]_13 ;
  input \stat_reg[0]_14 ;
  input \stat_reg[0]_15 ;
  input [10:0]out;
  input \stat_reg[1]_7 ;
  input \stat_reg[1]_8 ;
  input \ccmd[4]_INST_0_i_2 ;
  input brdy;
  input ctl_bcc_take1_fl;
  input ctl_bcc_take0_fl;
  input \stat_reg[0]_16 ;
  input rgf_sr_dr;
  input crdy;
  input [0:0]SR;
  input [2:0]D;
  input clk;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]Q;
  wire [0:0]SR;
  wire brdy;
  wire \ccmd[4]_INST_0_i_2 ;
  wire clk;
  wire crdy;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take1_fl;
  wire [10:0]out;
  wire rgf_sr_dr;
  wire \stat[0]_i_5__1_n_0 ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_12 ;
  wire \stat_reg[0]_13 ;
  wire \stat_reg[0]_14 ;
  wire \stat_reg[0]_15 ;
  wire \stat_reg[0]_16 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[10]),
        .O(\stat_reg[2]_4 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bcmd[2]_INST_0_i_10 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[9]),
        .I3(out[10]),
        .O(\stat_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hEFF0)) 
    \bdatw[15]_INST_0_i_230 
       (.I0(Q[1]),
        .I1(Q[2]),
        .I2(out[9]),
        .I3(out[8]),
        .O(\stat_reg[1]_2 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(Q[0]),
        .I1(out[2]),
        .O(\stat_reg[0]_11 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(Q[0]),
        .I1(out[7]),
        .I2(Q[1]),
        .O(\stat_reg[0]_12 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0_i_15 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\stat_reg[0]_10 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .O(\stat_reg[0]_3 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_19 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_5 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF0FEFF)) 
    \ccmd[4]_INST_0_i_10 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(out[6]),
        .I4(out[7]),
        .I5(\ccmd[4]_INST_0_i_2 ),
        .O(\stat_reg[0]_4 ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take0_fl_i_1
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(ctl_bcc_take0_fl),
        .O(\stat_reg[0]_13 ));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_35
       (.I0(Q[0]),
        .I1(out[3]),
        .O(\stat_reg[0]_5 ));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch0_fl_i_44
       (.I0(Q[2]),
        .I1(Q[0]),
        .O(\stat_reg[2]_3 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \fadr[15]_INST_0_i_14 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(out[5]),
        .I3(out[4]),
        .O(\stat_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF80)) 
    \fadr[15]_INST_0_i_3 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(ctl_bcc_take1_fl),
        .I4(ctl_bcc_take0_fl),
        .I5(\stat_reg[0]_16 ),
        .O(\stat_reg[0]_6 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[1]_i_9 
       (.I0(Q[1]),
        .I1(out[10]),
        .O(\stat_reg[1]_6 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[2]_i_6 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_1 ));
  LUT3 #(
    .INIT(8'hFD)) 
    \rgf_selc0_wb[1]_i_27 
       (.I0(out[7]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\stat_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \stat[0]_i_12__0 
       (.I0(Q[1]),
        .I1(out[10]),
        .I2(Q[2]),
        .I3(brdy),
        .O(\stat_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h88888888AAAAAAA8)) 
    \stat[0]_i_2 
       (.I0(\stat[0]_i_5__1_n_0 ),
        .I1(\stat_reg[0]_14 ),
        .I2(\stat_reg[1]_0 ),
        .I3(Q[2]),
        .I4(Q[0]),
        .I5(\stat_reg[0]_15 ),
        .O(\stat_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFBF0000FFAF00FF)) 
    \stat[0]_i_29__0 
       (.I0(Q[0]),
        .I1(rgf_sr_dr),
        .I2(crdy),
        .I3(Q[2]),
        .I4(out[2]),
        .I5(out[1]),
        .O(\stat_reg[0]_7 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \stat[0]_i_32 
       (.I0(out[6]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\stat_reg[0]_9 ));
  LUT6 #(
    .INIT(64'hEDEDEDEDEDEDEDFD)) 
    \stat[0]_i_35 
       (.I0(out[0]),
        .I1(Q[2]),
        .I2(out[2]),
        .I3(crdy),
        .I4(Q[1]),
        .I5(Q[0]),
        .O(\stat_reg[2]_2 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_5__1 
       (.I0(\stat_reg[1]_7 ),
        .I1(Q[2]),
        .I2(Q[1]),
        .I3(Q[0]),
        .O(\stat[0]_i_5__1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_7__1 
       (.I0(Q[1]),
        .I1(out[6]),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hBFBFFFCF0033FFFF)) 
    \stat[2]_i_11__0 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(brdy),
        .I3(Q[2]),
        .I4(out[0]),
        .I5(out[1]),
        .O(\stat_reg[0]_8 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8FFFA)) 
    \stat[2]_i_3__0 
       (.I0(\stat_reg[1]_7 ),
        .I1(\stat_reg[1]_8 ),
        .I2(Q[0]),
        .I3(Q[2]),
        .I4(out[6]),
        .I5(Q[1]),
        .O(\stat_reg[0]_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_6 
       (.I0(Q[1]),
        .I1(Q[2]),
        .O(\stat_reg[1]_4 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(Q[2]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_fsm" *) 
module mcss_fsm_1
   (\stat_reg[2]_0 ,
    \stat_reg[2]_1 ,
    Q,
    \stat_reg[2]_2 ,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    \stat_reg[1]_0 ,
    \stat_reg[1]_1 ,
    \stat_reg[1]_2 ,
    \stat_reg[1]_3 ,
    \stat_reg[0]_2 ,
    \stat_reg[1]_4 ,
    \stat_reg[0]_3 ,
    \stat_reg[0]_4 ,
    \stat_reg[1]_5 ,
    \stat_reg[1]_6 ,
    \stat_reg[1]_7 ,
    brdy_0,
    \stat_reg[0]_5 ,
    \stat_reg[2]_3 ,
    \stat_reg[1]_8 ,
    D,
    \stat_reg[2]_4 ,
    \stat_reg[2]_5 ,
    \stat_reg[2]_6 ,
    \stat_reg[2]_7 ,
    \rgf_selc1_rn_wb_reg[0] ,
    out,
    \stat_reg[2]_8 ,
    \sp[15]_i_6 ,
    brdy,
    ctl_bcc_take1_fl,
    SR,
    clk);
  output \stat_reg[2]_0 ;
  output \stat_reg[2]_1 ;
  output [2:0]Q;
  output \stat_reg[2]_2 ;
  output \stat_reg[0]_0 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[1]_0 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[1]_4 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[0]_4 ;
  output \stat_reg[1]_5 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[1]_7 ;
  output brdy_0;
  output \stat_reg[0]_5 ;
  output \stat_reg[2]_3 ;
  output \stat_reg[1]_8 ;
  input [1:0]D;
  input \stat_reg[2]_4 ;
  input \stat_reg[2]_5 ;
  input \stat_reg[2]_6 ;
  input \stat_reg[2]_7 ;
  input \rgf_selc1_rn_wb_reg[0] ;
  input [9:0]out;
  input \stat_reg[2]_8 ;
  input \sp[15]_i_6 ;
  input brdy;
  input ctl_bcc_take1_fl;
  input [0:0]SR;
  input clk;

  wire \<const1> ;
  wire [1:0]D;
  wire [2:0]Q;
  wire [0:0]SR;
  wire brdy;
  wire brdy_0;
  wire clk;
  wire ctl_bcc_take1_fl;
  wire [9:0]out;
  wire \rgf_selc1_rn_wb_reg[0] ;
  wire \sp[15]_i_6 ;
  wire \stat[2]_i_7__0_n_0 ;
  wire [2:2]stat_nx;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire \stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire \stat_reg[2]_7 ;
  wire \stat_reg[2]_8 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[15]_INST_0_i_172 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(out[9]),
        .O(\stat_reg[1]_5 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_228 
       (.I0(Q[0]),
        .I1(out[7]),
        .O(\stat_reg[0]_4 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badrx[15]_INST_0_i_4 
       (.I0(Q[1]),
        .I1(out[4]),
        .O(\stat_reg[1]_3 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(Q[1]),
        .I1(out[9]),
        .I2(Q[2]),
        .O(\stat_reg[1]_1 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[2]_INST_0_i_6 
       (.I0(Q[1]),
        .I1(Q[2]),
        .O(\stat_reg[1]_2 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bdatw[15]_INST_0_i_102 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .O(\stat_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take1_fl_i_1
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(ctl_bcc_take1_fl),
        .O(\stat_reg[0]_5 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_17 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \fadr[15]_INST_0_i_7 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .O(\stat_reg[2]_3 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_2 
       (.I0(Q[2]),
        .I1(\rgf_selc1_rn_wb_reg[0] ),
        .O(\stat_reg[2]_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_4 
       (.I0(Q[1]),
        .I1(out[9]),
        .O(\stat_reg[1]_6 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_17 
       (.I0(Q[1]),
        .I1(out[5]),
        .O(\stat_reg[1]_7 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_selc1_rn_wb[1]_i_18 
       (.I0(Q[1]),
        .I1(out[3]),
        .I2(Q[0]),
        .O(\stat_reg[1]_8 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_wb[0]_i_14 
       (.I0(Q[1]),
        .I1(out[5]),
        .O(\stat_reg[1]_4 ));
  LUT3 #(
    .INIT(8'hFD)) 
    \rgf_selc1_wb[1]_i_27 
       (.I0(out[6]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\stat_reg[0]_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_wb[1]_i_28 
       (.I0(Q[0]),
        .I1(out[6]),
        .I2(Q[1]),
        .O(\stat_reg[0]_2 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \sp[15]_i_12 
       (.I0(\sp[15]_i_6 ),
        .I1(brdy),
        .I2(Q[2]),
        .I3(out[9]),
        .I4(Q[1]),
        .O(brdy_0));
  LUT6 #(
    .INIT(64'hEAEEFFFFEAEEEAEE)) 
    \stat[2]_i_1__0 
       (.I0(\stat_reg[2]_0 ),
        .I1(\stat_reg[2]_1 ),
        .I2(\stat_reg[2]_4 ),
        .I3(\stat_reg[2]_5 ),
        .I4(\stat_reg[2]_6 ),
        .I5(\stat[2]_i_7__0_n_0 ),
        .O(stat_nx));
  LUT4 #(
    .INIT(16'h0001)) 
    \stat[2]_i_2__1 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(Q[0]),
        .I3(\stat_reg[2]_7 ),
        .O(\stat_reg[2]_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \stat[2]_i_3__1 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[8]),
        .I3(out[9]),
        .O(\stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h04003C3C03000000)) 
    \stat[2]_i_7__0 
       (.I0(Q[0]),
        .I1(Q[1]),
        .I2(Q[2]),
        .I3(\stat_reg[2]_8 ),
        .I4(out[1]),
        .I5(out[0]),
        .O(\stat[2]_i_7__0_n_0 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx),
        .Q(Q[2]),
        .R(SR));
  LUT2 #(
    .INIT(4'h7)) 
    tout__1_carry_i_35
       (.I0(Q[0]),
        .I1(out[2]),
        .O(\stat_reg[0]_3 ));
endmodule

module mcss_mem
   (.cbus_i_0_sp_1(cbus_i_0_sn_1),
    \read_cyc_reg[3] ,
    .cbus_i_3_sp_1(cbus_i_3_sn_1),
    \read_cyc_reg[3]_0 ,
    \read_cyc_reg[3]_1 ,
    \read_cyc_reg[3]_2 ,
    \read_cyc_reg[3]_3 ,
    \cbus_i[15] ,
    .bdatr_2_sp_1(bdatr_2_sn_1),
    \read_cyc_reg[2] ,
    .bdatr_6_sp_1(bdatr_6_sn_1),
    \read_cyc_reg[2]_0 ,
    \read_cyc_reg[2]_1 ,
    \read_cyc_reg[2]_2 ,
    \read_cyc_reg[2]_3 ,
    brdy_0,
    Q,
    \stat_reg[1] ,
    .fdatx_8_sp_1(fdatx_8_sn_1),
    \fdatx[8]_0 ,
    \fdat[8] ,
    \stat_reg[1]_0 ,
    .bdatr_15_sp_1(bdatr_15_sn_1),
    \read_cyc_reg[0] ,
    \read_cyc_reg[1] ,
    \read_cyc_reg[0]_0 ,
    \read_cyc_reg[1]_0 ,
    \read_cyc_reg[1]_1 ,
    \read_cyc_reg[1]_2 ,
    \read_cyc_reg[0]_1 ,
    \read_cyc_reg[3]_4 ,
    \read_cyc_reg[0]_2 ,
    \read_cyc_reg[3]_5 ,
    \read_cyc_reg[3]_6 ,
    \read_cyc_reg[3]_7 ,
    \read_cyc_reg[0]_3 ,
    brdy_1,
    brdy_2,
    out,
    clk,
    \rgf_c0bus_wb_reg[15] ,
    cbus_i,
    bdatr,
    \rgf_c1bus_wb_reg[14] ,
    O,
    \rgf_c1bus_wb_reg[6] ,
    \rgf_c1bus_wb_reg[9] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    brdy,
    \stat[2]_i_7__0 ,
    fch_memacc1,
    ir0_id,
    fch_irq_req_fl,
    fdatx,
    \ir0_id_fl[21]_i_5 ,
    \nir_id_reg[21] ,
    fdat,
    \nir_id[21]_i_2 ,
    \stat[0]_i_4 ,
    \stat[0]_i_24__0 ,
    D,
    SR,
    \read_cyc_reg[2]_4 );
  output \read_cyc_reg[3] ;
  output \read_cyc_reg[3]_0 ;
  output \read_cyc_reg[3]_1 ;
  output \read_cyc_reg[3]_2 ;
  output \read_cyc_reg[3]_3 ;
  output \cbus_i[15] ;
  output \read_cyc_reg[2] ;
  output \read_cyc_reg[2]_0 ;
  output \read_cyc_reg[2]_1 ;
  output \read_cyc_reg[2]_2 ;
  output \read_cyc_reg[2]_3 ;
  output brdy_0;
  output [1:0]Q;
  output \stat_reg[1] ;
  output \fdatx[8]_0 ;
  output [0:0]\fdat[8] ;
  output \stat_reg[1]_0 ;
  output \read_cyc_reg[0] ;
  output \read_cyc_reg[1] ;
  output \read_cyc_reg[0]_0 ;
  output \read_cyc_reg[1]_0 ;
  output \read_cyc_reg[1]_1 ;
  output \read_cyc_reg[1]_2 ;
  output \read_cyc_reg[0]_1 ;
  output \read_cyc_reg[3]_4 ;
  output \read_cyc_reg[0]_2 ;
  output \read_cyc_reg[3]_5 ;
  output \read_cyc_reg[3]_6 ;
  output \read_cyc_reg[3]_7 ;
  output \read_cyc_reg[0]_3 ;
  output brdy_1;
  output brdy_2;
  input out;
  input clk;
  input \rgf_c0bus_wb_reg[15] ;
  input [6:0]cbus_i;
  input [15:0]bdatr;
  input \rgf_c1bus_wb_reg[14] ;
  input [0:0]O;
  input [0:0]\rgf_c1bus_wb_reg[6] ;
  input [1:0]\rgf_c1bus_wb_reg[9] ;
  input [1:0]\rgf_c1bus_wb_reg[14]_0 ;
  input brdy;
  input \stat[2]_i_7__0 ;
  input fch_memacc1;
  input [0:0]ir0_id;
  input fch_irq_req_fl;
  input [15:0]fdatx;
  input \ir0_id_fl[21]_i_5 ;
  input \nir_id_reg[21] ;
  input [13:0]fdat;
  input \nir_id[21]_i_2 ;
  input [1:0]\stat[0]_i_4 ;
  input [1:0]\stat[0]_i_24__0 ;
  input [0:0]D;
  input [0:0]SR;
  input [2:0]\read_cyc_reg[2]_4 ;
  output cbus_i_0_sn_1;
  output cbus_i_3_sn_1;
  output bdatr_2_sn_1;
  output bdatr_6_sn_1;
  output fdatx_8_sn_1;
  output bdatr_15_sn_1;

  wire [0:0]D;
  wire [0:0]O;
  wire [1:0]Q;
  wire [0:0]SR;
  wire [15:0]bdatr;
  wire bdatr_15_sn_1;
  wire bdatr_2_sn_1;
  wire bdatr_6_sn_1;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire brdy_2;
  wire [6:0]cbus_i;
  wire \cbus_i[15] ;
  wire cbus_i_0_sn_1;
  wire cbus_i_3_sn_1;
  wire clk;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire [13:0]fdat;
  wire [0:0]\fdat[8] ;
  wire [15:0]fdatx;
  wire \fdatx[8]_0 ;
  wire fdatx_8_sn_1;
  wire [0:0]ir0_id;
  wire \ir0_id_fl[21]_i_5 ;
  wire \nir_id[21]_i_2 ;
  wire \nir_id_reg[21] ;
  wire out;
  wire \read_cyc_reg[0] ;
  wire \read_cyc_reg[0]_0 ;
  wire \read_cyc_reg[0]_1 ;
  wire \read_cyc_reg[0]_2 ;
  wire \read_cyc_reg[0]_3 ;
  wire \read_cyc_reg[1] ;
  wire \read_cyc_reg[1]_0 ;
  wire \read_cyc_reg[1]_1 ;
  wire \read_cyc_reg[1]_2 ;
  wire \read_cyc_reg[2] ;
  wire \read_cyc_reg[2]_0 ;
  wire \read_cyc_reg[2]_1 ;
  wire \read_cyc_reg[2]_2 ;
  wire \read_cyc_reg[2]_3 ;
  wire [2:0]\read_cyc_reg[2]_4 ;
  wire \read_cyc_reg[3] ;
  wire \read_cyc_reg[3]_0 ;
  wire \read_cyc_reg[3]_1 ;
  wire \read_cyc_reg[3]_2 ;
  wire \read_cyc_reg[3]_3 ;
  wire \read_cyc_reg[3]_4 ;
  wire \read_cyc_reg[3]_5 ;
  wire \read_cyc_reg[3]_6 ;
  wire \read_cyc_reg[3]_7 ;
  wire \rgf_c0bus_wb_reg[15] ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire [1:0]\rgf_c1bus_wb_reg[14]_0 ;
  wire [0:0]\rgf_c1bus_wb_reg[6] ;
  wire [1:0]\rgf_c1bus_wb_reg[9] ;
  wire [1:0]\stat[0]_i_24__0 ;
  wire [1:0]\stat[0]_i_4 ;
  wire \stat[2]_i_7__0 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;

  mcss_mem_bctl bctl
       (.D(D),
        .O(O),
        .Q(Q),
        .SR(SR),
        .bdatr(bdatr),
        .bdatr_15_sp_1(bdatr_15_sn_1),
        .bdatr_2_sp_1(bdatr_2_sn_1),
        .bdatr_6_sp_1(bdatr_6_sn_1),
        .brdy(brdy),
        .brdy_0(brdy_0),
        .brdy_1(brdy_1),
        .brdy_2(brdy_2),
        .cbus_i(cbus_i),
        .\cbus_i[15] (\cbus_i[15] ),
        .cbus_i_0_sp_1(cbus_i_0_sn_1),
        .cbus_i_3_sp_1(cbus_i_3_sn_1),
        .clk(clk),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_memacc1(fch_memacc1),
        .fdat(fdat),
        .\fdat[8] (\fdat[8] ),
        .fdatx(fdatx),
        .\fdatx[8]_0 (\fdatx[8]_0 ),
        .fdatx_8_sp_1(fdatx_8_sn_1),
        .ir0_id(ir0_id),
        .\ir0_id_fl[21]_i_5 (\ir0_id_fl[21]_i_5 ),
        .\nir_id[21]_i_2 (\nir_id[21]_i_2 ),
        .\nir_id_reg[21] (\nir_id_reg[21] ),
        .out(out),
        .\read_cyc_reg[0]_0 (\read_cyc_reg[0] ),
        .\read_cyc_reg[0]_1 (\read_cyc_reg[0]_0 ),
        .\read_cyc_reg[0]_2 (\read_cyc_reg[0]_1 ),
        .\read_cyc_reg[0]_3 (\read_cyc_reg[0]_2 ),
        .\read_cyc_reg[0]_4 (\read_cyc_reg[0]_3 ),
        .\read_cyc_reg[1]_0 (\read_cyc_reg[1] ),
        .\read_cyc_reg[1]_1 (\read_cyc_reg[1]_0 ),
        .\read_cyc_reg[1]_2 (\read_cyc_reg[1]_1 ),
        .\read_cyc_reg[1]_3 (\read_cyc_reg[1]_2 ),
        .\read_cyc_reg[2]_0 (\read_cyc_reg[2] ),
        .\read_cyc_reg[2]_1 (\read_cyc_reg[2]_0 ),
        .\read_cyc_reg[2]_2 (\read_cyc_reg[2]_1 ),
        .\read_cyc_reg[2]_3 (\read_cyc_reg[2]_2 ),
        .\read_cyc_reg[2]_4 (\read_cyc_reg[2]_3 ),
        .\read_cyc_reg[2]_5 (\read_cyc_reg[2]_4 ),
        .\read_cyc_reg[3]_0 (\read_cyc_reg[3] ),
        .\read_cyc_reg[3]_1 (\read_cyc_reg[3]_0 ),
        .\read_cyc_reg[3]_2 (\read_cyc_reg[3]_1 ),
        .\read_cyc_reg[3]_3 (\read_cyc_reg[3]_2 ),
        .\read_cyc_reg[3]_4 (\read_cyc_reg[3]_3 ),
        .\read_cyc_reg[3]_5 (\read_cyc_reg[3]_4 ),
        .\read_cyc_reg[3]_6 (\read_cyc_reg[3]_5 ),
        .\read_cyc_reg[3]_7 (\read_cyc_reg[3]_6 ),
        .\read_cyc_reg[3]_8 (\read_cyc_reg[3]_7 ),
        .\rgf_c0bus_wb_reg[15] (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[14] (\rgf_c1bus_wb_reg[14] ),
        .\rgf_c1bus_wb_reg[14]_0 (\rgf_c1bus_wb_reg[14]_0 ),
        .\rgf_c1bus_wb_reg[6] (\rgf_c1bus_wb_reg[6] ),
        .\rgf_c1bus_wb_reg[9] (\rgf_c1bus_wb_reg[9] ),
        .\stat[0]_i_24__0 (\stat[0]_i_24__0 ),
        .\stat[0]_i_4 (\stat[0]_i_4 ),
        .\stat[2]_i_7__0 (\stat[2]_i_7__0 ),
        .\stat_reg[1] (\stat_reg[1] ),
        .\stat_reg[1]_0 (\stat_reg[1]_0 ));
endmodule

module mcss_mem_bctl
   (.cbus_i_0_sp_1(cbus_i_0_sn_1),
    \read_cyc_reg[3]_0 ,
    .cbus_i_3_sp_1(cbus_i_3_sn_1),
    \read_cyc_reg[3]_1 ,
    \read_cyc_reg[3]_2 ,
    \read_cyc_reg[3]_3 ,
    \read_cyc_reg[3]_4 ,
    \cbus_i[15] ,
    .bdatr_2_sp_1(bdatr_2_sn_1),
    \read_cyc_reg[2]_0 ,
    .bdatr_6_sp_1(bdatr_6_sn_1),
    \read_cyc_reg[2]_1 ,
    \read_cyc_reg[2]_2 ,
    \read_cyc_reg[2]_3 ,
    \read_cyc_reg[2]_4 ,
    brdy_0,
    Q,
    \stat_reg[1] ,
    .fdatx_8_sp_1(fdatx_8_sn_1),
    \fdatx[8]_0 ,
    \fdat[8] ,
    \stat_reg[1]_0 ,
    .bdatr_15_sp_1(bdatr_15_sn_1),
    \read_cyc_reg[0]_0 ,
    \read_cyc_reg[1]_0 ,
    \read_cyc_reg[0]_1 ,
    \read_cyc_reg[1]_1 ,
    \read_cyc_reg[1]_2 ,
    \read_cyc_reg[1]_3 ,
    \read_cyc_reg[0]_2 ,
    \read_cyc_reg[3]_5 ,
    \read_cyc_reg[0]_3 ,
    \read_cyc_reg[3]_6 ,
    \read_cyc_reg[3]_7 ,
    \read_cyc_reg[3]_8 ,
    \read_cyc_reg[0]_4 ,
    brdy_1,
    brdy_2,
    out,
    clk,
    \rgf_c0bus_wb_reg[15] ,
    cbus_i,
    bdatr,
    \rgf_c1bus_wb_reg[14] ,
    O,
    \rgf_c1bus_wb_reg[6] ,
    \rgf_c1bus_wb_reg[9] ,
    \rgf_c1bus_wb_reg[14]_0 ,
    brdy,
    \stat[2]_i_7__0 ,
    fch_memacc1,
    ir0_id,
    fch_irq_req_fl,
    fdatx,
    \ir0_id_fl[21]_i_5 ,
    \nir_id_reg[21] ,
    fdat,
    \nir_id[21]_i_2 ,
    \stat[0]_i_4 ,
    \stat[0]_i_24__0 ,
    SR,
    D,
    \read_cyc_reg[2]_5 );
  output \read_cyc_reg[3]_0 ;
  output \read_cyc_reg[3]_1 ;
  output \read_cyc_reg[3]_2 ;
  output \read_cyc_reg[3]_3 ;
  output \read_cyc_reg[3]_4 ;
  output \cbus_i[15] ;
  output \read_cyc_reg[2]_0 ;
  output \read_cyc_reg[2]_1 ;
  output \read_cyc_reg[2]_2 ;
  output \read_cyc_reg[2]_3 ;
  output \read_cyc_reg[2]_4 ;
  output brdy_0;
  output [1:0]Q;
  output \stat_reg[1] ;
  output \fdatx[8]_0 ;
  output [0:0]\fdat[8] ;
  output \stat_reg[1]_0 ;
  output \read_cyc_reg[0]_0 ;
  output \read_cyc_reg[1]_0 ;
  output \read_cyc_reg[0]_1 ;
  output \read_cyc_reg[1]_1 ;
  output \read_cyc_reg[1]_2 ;
  output \read_cyc_reg[1]_3 ;
  output \read_cyc_reg[0]_2 ;
  output \read_cyc_reg[3]_5 ;
  output \read_cyc_reg[0]_3 ;
  output \read_cyc_reg[3]_6 ;
  output \read_cyc_reg[3]_7 ;
  output \read_cyc_reg[3]_8 ;
  output \read_cyc_reg[0]_4 ;
  output brdy_1;
  output brdy_2;
  input out;
  input clk;
  input \rgf_c0bus_wb_reg[15] ;
  input [6:0]cbus_i;
  input [15:0]bdatr;
  input \rgf_c1bus_wb_reg[14] ;
  input [0:0]O;
  input [0:0]\rgf_c1bus_wb_reg[6] ;
  input [1:0]\rgf_c1bus_wb_reg[9] ;
  input [1:0]\rgf_c1bus_wb_reg[14]_0 ;
  input brdy;
  input \stat[2]_i_7__0 ;
  input fch_memacc1;
  input [0:0]ir0_id;
  input fch_irq_req_fl;
  input [15:0]fdatx;
  input \ir0_id_fl[21]_i_5 ;
  input \nir_id_reg[21] ;
  input [13:0]fdat;
  input \nir_id[21]_i_2 ;
  input [1:0]\stat[0]_i_4 ;
  input [1:0]\stat[0]_i_24__0 ;
  input [0:0]SR;
  input [0:0]D;
  input [2:0]\read_cyc_reg[2]_5 ;
  output cbus_i_0_sn_1;
  output cbus_i_3_sn_1;
  output bdatr_2_sn_1;
  output bdatr_6_sn_1;
  output fdatx_8_sn_1;
  output bdatr_15_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]D;
  wire [0:0]O;
  wire [1:0]Q;
  wire [0:0]SR;
  wire [15:0]bdatr;
  wire bdatr_15_sn_1;
  wire bdatr_2_sn_1;
  wire bdatr_6_sn_1;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire brdy_2;
  wire [6:0]cbus_i;
  wire \cbus_i[15] ;
  wire cbus_i_0_sn_1;
  wire cbus_i_3_sn_1;
  wire clk;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire fch_term_fl;
  wire [13:0]fdat;
  wire [0:0]\fdat[8] ;
  wire [15:0]fdatx;
  wire \fdatx[8]_0 ;
  wire fdatx_8_sn_1;
  wire [0:0]ir0_id;
  wire \ir0_id_fl[21]_i_5 ;
  wire mem_accslot;
  wire \nir_id[21]_i_2 ;
  wire \nir_id_reg[21] ;
  wire out;
  wire [3:0]read_cyc;
  wire \read_cyc_reg[0]_0 ;
  wire \read_cyc_reg[0]_1 ;
  wire \read_cyc_reg[0]_2 ;
  wire \read_cyc_reg[0]_3 ;
  wire \read_cyc_reg[0]_4 ;
  wire \read_cyc_reg[1]_0 ;
  wire \read_cyc_reg[1]_1 ;
  wire \read_cyc_reg[1]_2 ;
  wire \read_cyc_reg[1]_3 ;
  wire \read_cyc_reg[2]_0 ;
  wire \read_cyc_reg[2]_1 ;
  wire \read_cyc_reg[2]_2 ;
  wire \read_cyc_reg[2]_3 ;
  wire \read_cyc_reg[2]_4 ;
  wire [2:0]\read_cyc_reg[2]_5 ;
  wire \read_cyc_reg[3]_0 ;
  wire \read_cyc_reg[3]_1 ;
  wire \read_cyc_reg[3]_2 ;
  wire \read_cyc_reg[3]_3 ;
  wire \read_cyc_reg[3]_4 ;
  wire \read_cyc_reg[3]_5 ;
  wire \read_cyc_reg[3]_6 ;
  wire \read_cyc_reg[3]_7 ;
  wire \read_cyc_reg[3]_8 ;
  wire \rgf_c0bus_wb[0]_i_10_n_0 ;
  wire \rgf_c0bus_wb[3]_i_8_n_0 ;
  wire \rgf_c0bus_wb[3]_i_9_n_0 ;
  wire \rgf_c0bus_wb_reg[15] ;
  wire \rgf_c1bus_wb[2]_i_13_n_0 ;
  wire \rgf_c1bus_wb[6]_i_13_n_0 ;
  wire \rgf_c1bus_wb[6]_i_14_n_0 ;
  wire \rgf_c1bus_wb_reg[14] ;
  wire [1:0]\rgf_c1bus_wb_reg[14]_0 ;
  wire [0:0]\rgf_c1bus_wb_reg[6] ;
  wire [1:0]\rgf_c1bus_wb_reg[9] ;
  wire [1:0]\stat[0]_i_24__0 ;
  wire [1:0]\stat[0]_i_4 ;
  wire \stat[2]_i_7__0 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  mcss_mem_fsm ctl
       (.D(mem_accslot),
        .Q(Q),
        .SR(SR),
        .brdy(brdy),
        .brdy_0(brdy_0),
        .brdy_1(brdy_1),
        .brdy_2(brdy_2),
        .clk(clk),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_memacc1(fch_memacc1),
        .fch_term_fl(fch_term_fl),
        .fdat(fdat),
        .\fdat[8] (\fdat[8] ),
        .fdatx(fdatx),
        .\fdatx[8]_0 (\fdatx[8]_0 ),
        .fdatx_8_sp_1(fdatx_8_sn_1),
        .ir0_id(ir0_id),
        .\ir0_id_fl[21]_i_5_0 (\ir0_id_fl[21]_i_5 ),
        .\nir_id[21]_i_2_0 (\nir_id[21]_i_2 ),
        .\nir_id_reg[21] (\nir_id_reg[21] ),
        .\stat[0]_i_24__0 (\stat[0]_i_24__0 ),
        .\stat[0]_i_4 (\stat[0]_i_4 ),
        .\stat[2]_i_7__0 (\stat[2]_i_7__0 ),
        .\stat_reg[0]_0 (D),
        .\stat_reg[1]_0 (\stat_reg[1] ),
        .\stat_reg[1]_1 (\stat_reg[1]_0 ));
  FDRE fch_term_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(out),
        .Q(fch_term_fl),
        .R(\<const0> ));
  FDRE \read_cyc_reg[0] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_5 [0]),
        .Q(read_cyc[0]),
        .R(SR));
  FDRE \read_cyc_reg[1] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_5 [1]),
        .Q(read_cyc[1]),
        .R(SR));
  FDRE \read_cyc_reg[2] 
       (.C(clk),
        .CE(brdy),
        .D(\read_cyc_reg[2]_5 [2]),
        .Q(read_cyc[2]),
        .R(SR));
  FDRE \read_cyc_reg[3] 
       (.C(clk),
        .CE(brdy),
        .D(mem_accslot),
        .Q(read_cyc[3]),
        .R(SR));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[0]_i_10 
       (.I0(bdatr[0]),
        .I1(read_cyc[0]),
        .I2(bdatr[8]),
        .O(\rgf_c0bus_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[0]_i_3 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[0]),
        .I2(\rgf_c0bus_wb[0]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .I4(bdatr[0]),
        .I5(\read_cyc_reg[3]_0 ),
        .O(cbus_i_0_sn_1));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[10]_i_18 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[10]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[3]),
        .O(\read_cyc_reg[3]_2 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[11]_i_20 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[11]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[4]),
        .O(\read_cyc_reg[3]_3 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[13]_i_15 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .O(\read_cyc_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[14]_i_3 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[14]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[5]),
        .O(\read_cyc_reg[3]_4 ));
  LUT6 #(
    .INIT(64'h88888F8888888888)) 
    \rgf_c0bus_wb[15]_i_5 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[6]),
        .I2(read_cyc[3]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(bdatr[15]),
        .O(\cbus_i[15] ));
  LUT6 #(
    .INIT(64'h0E000F0004000000)) 
    \rgf_c0bus_wb[1]_i_12 
       (.I0(read_cyc[0]),
        .I1(bdatr[9]),
        .I2(read_cyc[3]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(bdatr[1]),
        .O(\read_cyc_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h5000504050001000)) 
    \rgf_c0bus_wb[2]_i_14 
       (.I0(read_cyc[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(bdatr[2]),
        .I4(read_cyc[0]),
        .I5(bdatr[10]),
        .O(\read_cyc_reg[3]_5 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[3]_i_3 
       (.I0(\rgf_c0bus_wb_reg[15] ),
        .I1(cbus_i[1]),
        .I2(bdatr[3]),
        .I3(\read_cyc_reg[3]_0 ),
        .I4(\rgf_c0bus_wb[3]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .O(cbus_i_3_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[3]_i_8 
       (.I0(bdatr[3]),
        .I1(read_cyc[0]),
        .I2(bdatr[11]),
        .O(\rgf_c0bus_wb[3]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c0bus_wb[3]_i_9 
       (.I0(read_cyc[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .O(\rgf_c0bus_wb[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5000504050001000)) 
    \rgf_c0bus_wb[4]_i_34 
       (.I0(read_cyc[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(bdatr[4]),
        .I4(read_cyc[0]),
        .I5(bdatr[12]),
        .O(\read_cyc_reg[3]_6 ));
  LUT6 #(
    .INIT(64'h5000504050001000)) 
    \rgf_c0bus_wb[5]_i_14 
       (.I0(read_cyc[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(bdatr[5]),
        .I4(read_cyc[0]),
        .I5(bdatr[13]),
        .O(\read_cyc_reg[3]_7 ));
  LUT6 #(
    .INIT(64'h5000504050001000)) 
    \rgf_c0bus_wb[6]_i_12 
       (.I0(read_cyc[3]),
        .I1(read_cyc[1]),
        .I2(read_cyc[2]),
        .I3(bdatr[6]),
        .I4(read_cyc[0]),
        .I5(bdatr[14]),
        .O(\read_cyc_reg[3]_8 ));
  LUT6 #(
    .INIT(64'h0E000F0004000000)) 
    \rgf_c0bus_wb[7]_i_12 
       (.I0(read_cyc[0]),
        .I1(bdatr[15]),
        .I2(read_cyc[3]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(bdatr[7]),
        .O(\read_cyc_reg[0]_4 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[8]_i_14 
       (.I0(read_cyc[3]),
        .I1(read_cyc[2]),
        .I2(read_cyc[1]),
        .I3(bdatr[8]),
        .I4(\rgf_c0bus_wb_reg[15] ),
        .I5(cbus_i[2]),
        .O(\read_cyc_reg[3]_1 ));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[0]_i_5 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .I3(bdatr[0]),
        .I4(read_cyc[0]),
        .I5(bdatr[8]),
        .O(\read_cyc_reg[1]_3 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[12]_i_16 
       (.I0(read_cyc[2]),
        .I1(read_cyc[1]),
        .I2(read_cyc[3]),
        .O(\read_cyc_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h44F4444444444444)) 
    \rgf_c1bus_wb[13]_i_4 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(\rgf_c1bus_wb_reg[14]_0 [0]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[13]),
        .O(\read_cyc_reg[2]_3 ));
  LUT6 #(
    .INIT(64'h44F4444444444444)) 
    \rgf_c1bus_wb[14]_i_2 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(\rgf_c1bus_wb_reg[14]_0 [1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[14]),
        .O(\read_cyc_reg[2]_4 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[15]_i_6 
       (.I0(bdatr[15]),
        .I1(read_cyc[3]),
        .I2(read_cyc[1]),
        .I3(read_cyc[2]),
        .O(bdatr_15_sn_1));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[1]_i_16 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .I3(bdatr[1]),
        .I4(read_cyc[0]),
        .I5(bdatr[9]),
        .O(\read_cyc_reg[1]_2 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[2]_i_13 
       (.I0(bdatr[2]),
        .I1(read_cyc[0]),
        .I2(bdatr[10]),
        .O(\rgf_c1bus_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[2]_i_4 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(O),
        .I2(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .I4(bdatr[2]),
        .I5(\read_cyc_reg[2]_0 ),
        .O(bdatr_2_sn_1));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[3]_i_14 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .I3(bdatr[3]),
        .I4(read_cyc[0]),
        .I5(bdatr[11]),
        .O(\read_cyc_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[4]_i_17 
       (.I0(read_cyc[0]),
        .I1(bdatr[12]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[4]),
        .O(\read_cyc_reg[0]_1 ));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[5]_i_11 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .I3(bdatr[5]),
        .I4(read_cyc[0]),
        .I5(bdatr[13]),
        .O(\read_cyc_reg[1]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[6]_i_13 
       (.I0(bdatr[6]),
        .I1(read_cyc[0]),
        .I2(bdatr[14]),
        .O(\rgf_c1bus_wb[6]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c1bus_wb[6]_i_14 
       (.I0(read_cyc[1]),
        .I1(read_cyc[2]),
        .I2(read_cyc[3]),
        .O(\rgf_c1bus_wb[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[6]_i_4 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(\rgf_c1bus_wb_reg[6] ),
        .I2(bdatr[6]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\rgf_c1bus_wb[6]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .O(bdatr_6_sn_1));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[7]_i_14 
       (.I0(read_cyc[0]),
        .I1(bdatr[15]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[7]),
        .O(\read_cyc_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h2000FFFF20002000)) 
    \rgf_c1bus_wb[8]_i_4 
       (.I0(read_cyc[2]),
        .I1(read_cyc[1]),
        .I2(read_cyc[3]),
        .I3(bdatr[8]),
        .I4(\rgf_c1bus_wb_reg[14] ),
        .I5(\rgf_c1bus_wb_reg[9] [0]),
        .O(\read_cyc_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h44F4444444444444)) 
    \rgf_c1bus_wb[9]_i_4 
       (.I0(\rgf_c1bus_wb_reg[14] ),
        .I1(\rgf_c1bus_wb_reg[9] [1]),
        .I2(read_cyc[2]),
        .I3(read_cyc[1]),
        .I4(read_cyc[3]),
        .I5(bdatr[9]),
        .O(\read_cyc_reg[2]_2 ));
  LUT6 #(
    .INIT(64'h0E000F0004000000)) 
    \sr[3]_i_9 
       (.I0(read_cyc[0]),
        .I1(bdatr[11]),
        .I2(read_cyc[3]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(bdatr[3]),
        .O(\read_cyc_reg[0]_3 ));
endmodule

module mcss_mem_fsm
   (brdy_0,
    Q,
    D,
    \stat_reg[1]_0 ,
    .fdatx_8_sp_1(fdatx_8_sn_1),
    \fdatx[8]_0 ,
    \fdat[8] ,
    \stat_reg[1]_1 ,
    brdy_1,
    brdy_2,
    brdy,
    fch_term_fl,
    \stat[2]_i_7__0 ,
    fch_memacc1,
    ir0_id,
    fch_irq_req_fl,
    fdatx,
    \ir0_id_fl[21]_i_5_0 ,
    \nir_id_reg[21] ,
    fdat,
    \nir_id[21]_i_2_0 ,
    \stat[0]_i_4 ,
    \stat[0]_i_24__0 ,
    SR,
    clk,
    \stat_reg[0]_0 );
  output brdy_0;
  output [1:0]Q;
  output [0:0]D;
  output \stat_reg[1]_0 ;
  output \fdatx[8]_0 ;
  output [0:0]\fdat[8] ;
  output \stat_reg[1]_1 ;
  output brdy_1;
  output brdy_2;
  input brdy;
  input fch_term_fl;
  input \stat[2]_i_7__0 ;
  input fch_memacc1;
  input [0:0]ir0_id;
  input fch_irq_req_fl;
  input [15:0]fdatx;
  input \ir0_id_fl[21]_i_5_0 ;
  input \nir_id_reg[21] ;
  input [13:0]fdat;
  input \nir_id[21]_i_2_0 ;
  input [1:0]\stat[0]_i_4 ;
  input [1:0]\stat[0]_i_24__0 ;
  input [0:0]SR;
  input clk;
  input [0:0]\stat_reg[0]_0 ;
  output fdatx_8_sn_1;

  wire \<const1> ;
  wire [0:0]D;
  wire [1:0]Q;
  wire [0:0]SR;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire brdy_2;
  wire clk;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire fch_term_fl;
  wire [13:0]fdat;
  wire [0:0]\fdat[8] ;
  wire [15:0]fdatx;
  wire \fdatx[8]_0 ;
  wire fdatx_8_sn_1;
  wire [0:0]ir0_id;
  wire \ir0_id_fl[21]_i_10_n_0 ;
  wire \ir0_id_fl[21]_i_11_n_0 ;
  wire \ir0_id_fl[21]_i_5_0 ;
  wire \ir0_id_fl[21]_i_5_n_0 ;
  wire \ir0_id_fl[21]_i_6_n_0 ;
  wire \ir0_id_fl[21]_i_7_n_0 ;
  wire \ir0_id_fl[21]_i_8_n_0 ;
  wire \ir0_id_fl[21]_i_9_n_0 ;
  wire \nir_id[21]_i_2_0 ;
  wire \nir_id[21]_i_2_n_0 ;
  wire \nir_id[21]_i_4_n_0 ;
  wire \nir_id[21]_i_5_n_0 ;
  wire \nir_id[21]_i_6_n_0 ;
  wire \nir_id[21]_i_7_n_0 ;
  wire \nir_id[21]_i_8_n_0 ;
  wire \nir_id[21]_i_9_n_0 ;
  wire \nir_id_reg[21] ;
  wire [1:0]\stat[0]_i_24__0 ;
  wire [1:0]\stat[0]_i_4 ;
  wire \stat[2]_i_7__0 ;
  wire [1:1]stat_nx;
  wire [0:0]\stat_reg[0]_0 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;

  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'hFFF30000FFFBFFFF)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(Q[1]),
        .I1(fch_memacc1),
        .I2(ir0_id),
        .I3(fch_irq_req_fl),
        .I4(fch_term_fl),
        .I5(Q[0]),
        .O(\stat_reg[1]_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_166
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(\fdatx[8]_0 ));
  LUT6 #(
    .INIT(64'hF600000000000000)) 
    \ir0_id_fl[21]_i_10 
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(\ir0_id_fl[21]_i_11_n_0 ),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(\ir0_id_fl[21]_i_5_0 ),
        .O(\ir0_id_fl[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hC1C0000000000000)) 
    \ir0_id_fl[21]_i_11 
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[6]),
        .I3(fdatx[3]),
        .I4(fdatx[7]),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[21]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAEAAAA)) 
    \ir0_id_fl[21]_i_3 
       (.I0(\ir0_id_fl[21]_i_5_n_0 ),
        .I1(\ir0_id_fl[21]_i_6_n_0 ),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(\ir0_id_fl[21]_i_7_n_0 ),
        .I5(fdatx[15]),
        .O(fdatx_8_sn_1));
  LUT6 #(
    .INIT(64'h00000000FFFFFF76)) 
    \ir0_id_fl[21]_i_5 
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .I2(fdatx[4]),
        .I3(\ir0_id_fl[21]_i_8_n_0 ),
        .I4(\ir0_id_fl[21]_i_9_n_0 ),
        .I5(\ir0_id_fl[21]_i_10_n_0 ),
        .O(\ir0_id_fl[21]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[21]_i_6 
       (.I0(fdatx[3]),
        .I1(fdatx[5]),
        .O(\ir0_id_fl[21]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[21]_i_7 
       (.I0(fdatx[0]),
        .I1(fdatx[1]),
        .O(\ir0_id_fl[21]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h3FFF3FFE)) 
    \ir0_id_fl[21]_i_8 
       (.I0(fdatx[5]),
        .I1(fdatx[12]),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .I4(fdatx[6]),
        .O(\ir0_id_fl[21]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5FFF5FFFFFFFFFFD)) 
    \ir0_id_fl[21]_i_9 
       (.I0(\fdatx[8]_0 ),
        .I1(fdatx[2]),
        .I2(fdatx[11]),
        .I3(fdatx[7]),
        .I4(fdatx[3]),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAAA2)) 
    \nir_id[21]_i_1 
       (.I0(\nir_id[21]_i_2_n_0 ),
        .I1(\nir_id_reg[21] ),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(\nir_id[21]_i_4_n_0 ),
        .I5(fdat[13]),
        .O(\fdat[8] ));
  LUT6 #(
    .INIT(64'hAAAAEAEBAAAAAAAA)) 
    \nir_id[21]_i_2 
       (.I0(\nir_id[21]_i_5_n_0 ),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(fdat[4]),
        .I4(\nir_id[21]_i_6_n_0 ),
        .I5(\nir_id[21]_i_7_n_0 ),
        .O(\nir_id[21]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[21]_i_4 
       (.I0(fdat[1]),
        .I1(fdat[3]),
        .O(\nir_id[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF600000000000000)) 
    \nir_id[21]_i_5 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .I2(\nir_id[21]_i_8_n_0 ),
        .I3(\nir_id[21]_i_2_0 ),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[21]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h5FFF5FFE)) 
    \nir_id[21]_i_6 
       (.I0(fdat[11]),
        .I1(fdat[3]),
        .I2(fdat[10]),
        .I3(fdat[9]),
        .I4(fdat[2]),
        .O(\nir_id[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hA000A00000000002)) 
    \nir_id[21]_i_7 
       (.I0(\nir_id[21]_i_9_n_0 ),
        .I1(fdat[0]),
        .I2(fdat[9]),
        .I3(fdat[5]),
        .I4(fdat[1]),
        .I5(fdat[8]),
        .O(\nir_id[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAA04000000000000)) 
    \nir_id[21]_i_8 
       (.I0(fdat[4]),
        .I1(fdat[1]),
        .I2(fdat[2]),
        .I3(fdat[3]),
        .I4(fdat[5]),
        .I5(fdat[8]),
        .O(\nir_id[21]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[21]_i_9 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[21]_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \read_cyc[3]_i_1 
       (.I0(\stat_reg[1]_0 ),
        .O(D));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[2]_i_9 
       (.I0(\stat_reg[1]_0 ),
        .I1(brdy),
        .I2(\stat[0]_i_24__0 [1]),
        .O(brdy_1));
  LUT3 #(
    .INIT(8'h40)) 
    \sr[15]_i_8 
       (.I0(\stat_reg[1]_0 ),
        .I1(brdy),
        .I2(\stat[0]_i_24__0 [0]),
        .O(brdy_2));
  LUT4 #(
    .INIT(16'h1FF1)) 
    \stat[0]_i_9__1 
       (.I0(Q[1]),
        .I1(fch_term_fl),
        .I2(\stat[0]_i_4 [0]),
        .I3(\stat[0]_i_4 [1]),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hF2F2F222AAAAAAAA)) 
    \stat[1]_i_1__2 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(fch_memacc1),
        .I3(ir0_id),
        .I4(fch_irq_req_fl),
        .I5(fch_term_fl),
        .O(stat_nx));
  LUT6 #(
    .INIT(64'h88080808A8080808)) 
    \stat[2]_i_16 
       (.I0(brdy),
        .I1(Q[0]),
        .I2(fch_term_fl),
        .I3(\stat[2]_i_7__0 ),
        .I4(fch_memacc1),
        .I5(Q[1]),
        .O(brdy_0));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat_reg[0]_0 ),
        .Q(Q[0]),
        .R(SR));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(stat_nx),
        .Q(Q[1]),
        .R(SR));
endmodule

module mcss_rgf
   (rgf_selc0_stat,
    rgf_selc1_stat,
    out,
    \grn_reg[15] ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[4]_2 ,
    \grn_reg[4]_3 ,
    \grn_reg[15]_0 ,
    \grn_reg[4]_4 ,
    \grn_reg[4]_5 ,
    \grn_reg[4]_6 ,
    \grn_reg[4]_7 ,
    \sr_reg[15] ,
    \pc_reg[15] ,
    \sp_reg[0] ,
    \iv_reg[15] ,
    \tr_reg[15] ,
    \sr_reg[4] ,
    \sr_reg[5] ,
    \pc_reg[15]_0 ,
    D,
    \pc_reg[14] ,
    \pc_reg[13] ,
    SR,
    \sp_reg[1] ,
    \sp_reg[15] ,
    \sp_reg[1]_0 ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[5] ,
    \sp_reg[6] ,
    \sp_reg[7] ,
    \sp_reg[8] ,
    \sp_reg[9] ,
    \sp_reg[10] ,
    \sp_reg[11] ,
    \sp_reg[12] ,
    \sp_reg[13] ,
    \sp_reg[14] ,
    bdatw,
    \tr_reg[14] ,
    \tr_reg[14]_0 ,
    \stat_reg[1] ,
    \tr_reg[13] ,
    \tr_reg[13]_0 ,
    \stat_reg[1]_0 ,
    \tr_reg[12] ,
    \tr_reg[11] ,
    \tr_reg[10] ,
    \tr_reg[9] ,
    \tr_reg[8] ,
    \stat_reg[1]_1 ,
    \tr_reg[7] ,
    \tr_reg[7]_0 ,
    \stat_reg[2] ,
    \tr_reg[6] ,
    a1bus_0,
    \badr[6]_INST_0_i_1 ,
    \tr_reg[6]_0 ,
    \stat_reg[2]_0 ,
    \tr_reg[5] ,
    \badr[5]_INST_0_i_1 ,
    \tr_reg[5]_0 ,
    \rgf_c1bus_wb[13]_i_9 ,
    \rgf_c1bus_wb[14]_i_30 ,
    \sr_reg[6] ,
    \badr[15]_INST_0_i_1 ,
    \sr_reg[6]_0 ,
    \sr_reg[6]_1 ,
    \badr[3]_INST_0_i_1 ,
    \sr[4]_i_156 ,
    \tr_reg[11]_0 ,
    \tr_reg[13]_1 ,
    \badr[15]_INST_0_i_1_0 ,
    \badr[1]_INST_0_i_1 ,
    \sr_reg[6]_2 ,
    \badr[9]_INST_0_i_1 ,
    \sr_reg[6]_3 ,
    \rgf_c1bus_wb[15]_i_14 ,
    \badr[10]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1_0 ,
    \badr[2]_INST_0_i_1 ,
    \rgf_c1bus_wb[11]_i_13 ,
    \badr[10]_INST_0_i_1_0 ,
    \badr[14]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_14_0 ,
    \badr[3]_INST_0_i_1_0 ,
    \badr[7]_INST_0_i_1 ,
    \badr[15]_INST_0_i_1_1 ,
    \sr_reg[6]_4 ,
    \badr[6]_INST_0_i_1_1 ,
    \sr_reg[6]_5 ,
    \rgf_c1bus_wb[12]_i_20 ,
    \rgf_c1bus_wb[11]_i_10 ,
    \badr[15]_INST_0_i_1_2 ,
    \rgf_c1bus_wb[14]_i_28 ,
    \rgf_c1bus_wb[15]_i_14_1 ,
    \rgf_c1bus_wb[14]_i_28_0 ,
    \rgf_c1bus_wb[7]_i_4 ,
    \badr[5]_INST_0_i_1_0 ,
    \sr[4]_i_219 ,
    \tr_reg[12]_0 ,
    \rgf_c1bus_wb[11]_i_10_0 ,
    \rgf_c1bus_wb[4]_i_9 ,
    \badr[12]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_28_1 ,
    \sr_reg[6]_6 ,
    \badr[0]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_28_2 ,
    \rgf_c1bus_wb[14]_i_28_3 ,
    \rgf_c1bus_wb[9]_i_17 ,
    \badr[10]_INST_0_i_1_1 ,
    \rgf_c1bus_wb[14]_i_28_4 ,
    \rgf_c1bus_wb[13]_i_16 ,
    \rgf_c1bus_wb[14]_i_28_5 ,
    \rgf_c1bus_wb[4]_i_9_0 ,
    \sr_reg[6]_7 ,
    \tr_reg[1] ,
    \sr_reg[6]_8 ,
    \tr_reg[14]_1 ,
    \sr_reg[6]_9 ,
    \sr_reg[6]_10 ,
    \rgf_c1bus_wb[15]_i_14_2 ,
    \badr[11]_INST_0_i_1 ,
    \sr_reg[6]_11 ,
    \sr_reg[6]_12 ,
    \badr[2]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[15]_i_14_3 ,
    \rgf_c1bus_wb[14]_i_28_6 ,
    \badr[9]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[14]_i_28_7 ,
    \rgf_c1bus_wb[14]_i_32 ,
    \badr[13]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1_1 ,
    \rgf_c1bus_wb[14]_i_32_0 ,
    \sr_reg[6]_13 ,
    \sr_reg[6]_14 ,
    \badr[14]_INST_0_i_1_0 ,
    \stat_reg[2]_1 ,
    \sr_reg[6]_15 ,
    \rgf_c1bus_wb[11]_i_10_1 ,
    \rgf_c1bus_wb[1]_i_14 ,
    \badr[6]_INST_0_i_1_2 ,
    \rgf_c1bus_wb[11]_i_10_2 ,
    \sr_reg[6]_16 ,
    \sr_reg[6]_17 ,
    \rgf_c1bus_wb[4]_i_28 ,
    \tr_reg[12]_1 ,
    \sr[4]_i_220 ,
    \tr_reg[3] ,
    \rgf_c1bus_wb[11]_i_10_3 ,
    \rgf_c1bus_wb[11]_i_10_4 ,
    \rgf_c1bus_wb[15]_i_27 ,
    \sr_reg[6]_18 ,
    \grn_reg[15]_1 ,
    \tr_reg[15]_0 ,
    \sr_reg[15]_0 ,
    \sp_reg[15]_0 ,
    \tr_reg[1]_0 ,
    \tr_reg[14]_2 ,
    \stat_reg[2]_2 ,
    \stat_reg[2]_3 ,
    \tr_reg[15]_1 ,
    \grn_reg[4]_8 ,
    \grn_reg[4]_9 ,
    \tr_reg[12]_2 ,
    \tr_reg[11]_1 ,
    \tr_reg[10]_0 ,
    \tr_reg[9]_0 ,
    \tr_reg[8]_0 ,
    \rgf_c0bus_wb[15]_i_18 ,
    \rgf_c0bus_wb[11]_i_3 ,
    a0bus_0,
    \rgf_c0bus_wb[11]_i_3_0 ,
    \badr[6]_INST_0_i_2 ,
    \sr[4]_i_133 ,
    \rgf_c0bus_wb[4]_i_26 ,
    \rgf_c0bus_wb[11]_i_9 ,
    \sr[4]_i_200 ,
    \sr[4]_i_195 ,
    \rgf_c0bus_wb[11]_i_9_0 ,
    \rgf_c0bus_wb[4]_i_32 ,
    \rgf_c0bus_wb[13]_i_27 ,
    \sr_reg[6]_19 ,
    \rgf_c0bus_wb[11]_i_11 ,
    \badr[5]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \badr[13]_INST_0_i_2 ,
    \badr[9]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_11_0 ,
    \rgf_c0bus_wb[11]_i_22 ,
    \badr[8]_INST_0_i_2 ,
    \badr[3]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_9_1 ,
    \badr[10]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2_0 ,
    \badr[2]_INST_0_i_2 ,
    \rgf_c0bus_wb[15]_i_25 ,
    \rgf_c0bus_wb[11]_i_8 ,
    \badr[4]_INST_0_i_2 ,
    \rgf_c0bus_wb[0]_i_14 ,
    \sr_reg[6]_20 ,
    \sr_reg[6]_21 ,
    \badr[10]_INST_0_i_2_0 ,
    \badr[14]_INST_0_i_2 ,
    \rgf_c0bus_wb[13]_i_29 ,
    \badr[4]_INST_0_i_2_0 ,
    \badr[12]_INST_0_i_2 ,
    \badr[8]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[7]_i_7 ,
    \rgf_c0bus_wb[7]_i_7_0 ,
    \sr_reg[6]_22 ,
    \sr_reg[6]_23 ,
    \badr[14]_INST_0_i_2_0 ,
    \sr_reg[6]_24 ,
    \rgf_c0bus_wb[11]_i_11_1 ,
    \badr[6]_INST_0_i_2_1 ,
    \rgf_c0bus_wb[11]_i_11_2 ,
    \badr[13]_INST_0_i_2_0 ,
    \badr[5]_INST_0_i_2_0 ,
    \badr[9]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[15]_i_26 ,
    \sr_reg[6]_25 ,
    \sp_reg[2]_0 ,
    \rgf_c0bus_wb[13]_i_30 ,
    \sr_reg[6]_26 ,
    \sr_reg[6]_27 ,
    \sp_reg[13]_0 ,
    \sp_reg[11]_0 ,
    \sr_reg[6]_28 ,
    \rgf_c0bus_wb[4]_i_29 ,
    \badr[3]_INST_0_i_2_0 ,
    \sr_reg[6]_29 ,
    \rgf_c0bus_wb[4]_i_33 ,
    \rgf_c0bus_wb[4]_i_31 ,
    \badr[11]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_22_0 ,
    \sr[4]_i_232 ,
    \sp_reg[1]_1 ,
    \badr[2]_INST_0_i_2_0 ,
    \sr_reg[6]_30 ,
    \rgf_c0bus_wb[12]_i_24 ,
    \sp_reg[4]_0 ,
    \sr_reg[14] ,
    \sr_reg[6]_31 ,
    \sr_reg[6]_32 ,
    \rgf_c0bus_wb[10]_i_8 ,
    \rgf_c0bus_wb[11]_i_9_2 ,
    \badr[1]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[13]_i_28 ,
    \sr_reg[6]_33 ,
    \badr[14]_INST_0_i_2_1 ,
    \rgf_c0bus_wb[8]_i_6 ,
    \rgf_c0bus_wb[12]_i_25 ,
    \sr_reg[6]_34 ,
    \sr_reg[6]_35 ,
    \sr_reg[6]_36 ,
    \sr_reg[6]_37 ,
    \badr[8]_INST_0_i_2_1 ,
    \badr[12]_INST_0_i_2_0 ,
    \sr_reg[6]_38 ,
    \badr[15]_INST_0_i_2 ,
    \sp_reg[0]_0 ,
    \sr_reg[0] ,
    \rgf_c0bus_wb[11]_i_3_1 ,
    \sr_reg[6]_39 ,
    fadr,
    fch_irq_req,
    badrx,
    \sr_reg[4]_0 ,
    \sr_reg[5]_0 ,
    \sr_reg[7] ,
    \sr_reg[5]_1 ,
    \sr_reg[6]_40 ,
    \sr_reg[5]_2 ,
    \sr_reg[6]_41 ,
    irq_0,
    \sr_reg[10] ,
    \sr_reg[4]_1 ,
    \fdatx[15] ,
    .fdat_12_sp_1(fdat_12_sn_1),
    S,
    \pc_reg[1] ,
    \pc_reg[15]_1 ,
    \rgf_c1bus_wb[7]_i_4_0 ,
    \sr_reg[6]_42 ,
    \rgf_c1bus_wb[11]_i_10_5 ,
    \rgf_c0bus_wb[15]_i_6 ,
    \rgf_c0bus_wb[15]_i_6_0 ,
    \rgf_c0bus_wb[15]_i_6_1 ,
    bbus_o,
    \rgf_c0bus_wb[11]_i_3_2 ,
    \rgf_c0bus_wb[11]_i_9_3 ,
    \rgf_c0bus_wb[11]_i_9_4 ,
    \rgf_c0bus_wb[11]_i_3_3 ,
    \sr_reg[5]_3 ,
    \sr_reg[5]_4 ,
    \sr_reg[5]_5 ,
    \fdat[15] ,
    \sr_reg[0]_0 ,
    \badr[14]_INST_0_i_1_1 ,
    \badr[13]_INST_0_i_1_0 ,
    \badr[14]_INST_0_i_2_2 ,
    \badr[6]_INST_0_i_1_3 ,
    tout__1_carry__0_i_1__0,
    \badr[10]_INST_0_i_1_2 ,
    tout__1_carry__1_i_1__0,
    \sr_reg[0]_1 ,
    \rgf_selc0_rn_wb_reg[2] ,
    \rgf_selc0_wb_reg[1] ,
    \rgf_selc1_rn_wb_reg[2] ,
    \rgf_selc1_wb_reg[1] ,
    \rgf_c0bus_wb_reg[15] ,
    \rgf_c1bus_wb_reg[15] ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \sp_reg[4]_1 ,
    \sp_reg[3]_0 ,
    \sp_reg[2]_1 ,
    \sp_reg[1]_2 ,
    \sp_reg[0]_1 ,
    \tr_reg[0] ,
    \tr_reg[1]_1 ,
    \tr_reg[2] ,
    \tr_reg[3]_0 ,
    \tr_reg[4] ,
    \iv_reg[15]_0 ,
    \sr_reg[15]_1 ,
    \sr_reg[4]_2 ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sr_reg[0]_2 ,
    \tr_reg[0]_0 ,
    \tr_reg[1]_2 ,
    \tr_reg[2]_0 ,
    \tr_reg[3]_1 ,
    \tr_reg[4]_0 ,
    \sp_reg[0]_2 ,
    \sp_reg[1]_3 ,
    \sp_reg[2]_2 ,
    \sp_reg[3]_1 ,
    \sp_reg[4]_2 ,
    b1bus_b02,
    E,
    p_2_in,
    clk,
    \rgf_selc1_wb_reg[0] ,
    rgf_selc1_stat_reg,
    \rgf_c1bus_wb_reg[0] ,
    rst_n,
    \sr_reg[5]_6 ,
    \pc_reg[13]_0 ,
    \sp_reg[14]_0 ,
    \sp_reg[14]_1 ,
    \bdatw[13] ,
    \bdatw[13]_0 ,
    \bdatw[13]_1 ,
    \bdatw[14] ,
    \bdatw[14]_0 ,
    \bdatw[13]_2 ,
    \bdatw[13]_3 ,
    \bdatw[12] ,
    \bdatw[12]_0 ,
    \bdatw[11] ,
    \bdatw[11]_0 ,
    \bdatw[10] ,
    \bdatw[10]_0 ,
    \bdatw[9] ,
    \bdatw[9]_0 ,
    \bdatw[8] ,
    \bdatw[8]_0 ,
    \rgf_c1bus_wb[15]_i_19 ,
    \rgf_c1bus_wb[15]_i_19_0 ,
    \rgf_c1bus_wb_reg[5] ,
    \sr[6]_i_15 ,
    \rgf_c1bus_wb[5]_i_10 ,
    \rgf_c1bus_wb[14]_i_11 ,
    \rgf_c1bus_wb[14]_i_11_0 ,
    tout__1_carry__0_i_7__0,
    tout__1_carry__0_i_7__0_0,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[5]_1 ,
    \rgf_c1bus_wb_reg[7] ,
    \sr[6]_i_11 ,
    \sr[6]_i_11_0 ,
    \sr[4]_i_27 ,
    \sr[6]_i_11_1 ,
    \sr[4]_i_30 ,
    \rgf_c1bus_wb[12]_i_2 ,
    \rgf_c1bus_wb_reg[3] ,
    \sr[4]_i_38 ,
    \rgf_c1bus_wb_reg[4] ,
    \sr[4]_i_44 ,
    \rgf_c1bus_wb_reg[10] ,
    \sr[4]_i_84 ,
    \bdatw[15] ,
    \bdatw[15]_0 ,
    \bdatw[14]_1 ,
    \bdatw[14]_2 ,
    \bdatw[13]_4 ,
    \bdatw[13]_5 ,
    \bdatw[12]_1 ,
    \bdatw[12]_2 ,
    \bdatw[11]_1 ,
    \bdatw[11]_2 ,
    \bdatw[10]_1 ,
    \bdatw[10]_2 ,
    \bdatw[9]_1 ,
    \bdatw[9]_2 ,
    \bdatw[8]_1 ,
    \bdatw[8]_2 ,
    \rgf_c0bus_wb_reg[7]_i_11 ,
    \sr[4]_i_67 ,
    \rgf_c0bus_wb[6]_i_11 ,
    \rgf_c0bus_wb[14]_i_2 ,
    \bbus_o[7] ,
    \bbus_o[7]_0 ,
    \bbus_o[6] ,
    \bbus_o[6]_0 ,
    \bbus_o[5] ,
    \bbus_o[5]_0 ,
    \sr[4]_i_15 ,
    \sr[4]_i_15_0 ,
    \sr[4]_i_15_1 ,
    \rgf_c0bus_wb_reg[10] ,
    \sr[4]_i_66 ,
    \rgf_c0bus_wb_reg[10]_0 ,
    \rgf_c0bus_wb_reg[10]_1 ,
    \rgf_c0bus_wb[12]_i_2 ,
    \sr[4]_i_55 ,
    \rgf_c0bus_wb[13]_i_4 ,
    \rgf_c0bus_wb[10]_i_4 ,
    \rgf_c0bus_wb[3]_i_7 ,
    \rgf_c0bus_wb[3]_i_7_0 ,
    \sr[4]_i_129 ,
    \rgf_c0bus_wb[15]_i_14 ,
    \pc0_reg[15] ,
    \fadr[15] ,
    O,
    \fadr[15]_0 ,
    \pc0_reg[15]_0 ,
    \pc0_reg[15]_1 ,
    .badrx_15_sp_1(badrx_15_sn_1),
    \badr[15]_INST_0_i_208 ,
    \rgf_selc1_wb[1]_i_16 ,
    irq,
    irq_lev,
    Q,
    ctl_fetch1_fl_i_15,
    fdatx,
    \ir0_id_fl[20]_i_4 ,
    fdat,
    \nir_id_reg[20] ,
    \bbus_o[5]_1 ,
    b0bus_sel_0,
    a1bus_sel_0,
    tout__1_carry__2,
    tout__1_carry__2_0,
    tout__1_carry__2_1,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \rgf_c1bus_wb_reg[15]_0 ,
    a0bus_sel_0,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_43 ,
    ctl_sela0,
    \i_/badr[15]_INST_0_i_43_0 ,
    \i_/bdatw[15]_INST_0_i_9 ,
    \i_/bdatw[15]_INST_0_i_9_0 ,
    \i_/bdatw[15]_INST_0_i_9_1 ,
    \i_/bdatw[15]_INST_0_i_9_2 ,
    ctl_selb0_0,
    \i_/bdatw[15]_INST_0_i_24 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_77 ,
    \i_/bdatw[15]_INST_0_i_9_3 ,
    \i_/bdatw[15]_INST_0_i_24_0 ,
    \i_/badr[15]_INST_0_i_19 ,
    \i_/badr[15]_INST_0_i_19_0 ,
    \i_/badr[15]_INST_0_i_19_1 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_113 ,
    \i_/bdatw[15]_INST_0_i_44 ,
    \i_/bdatw[15]_INST_0_i_112 ,
    \i_/bdatw[15]_INST_0_i_112_0 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_112_1 ,
    \rgf_c1bus_wb[4]_i_47 ,
    \rgf_c1bus_wb[4]_i_41 ,
    \rgf_c1bus_wb[4]_i_51 ,
    \sr[4]_i_235 ,
    \rgf_c1bus_wb[4]_i_65 ,
    \sr[4]_i_237 ,
    \rgf_c1bus_wb[4]_i_61 ,
    \rgf_c1bus_wb[4]_i_57 ,
    \sr[4]_i_245 ,
    \rgf_c1bus_wb[4]_i_53 ,
    \sr[4]_i_243 ,
    \rgf_c1bus_wb[4]_i_33 ,
    \rgf_c1bus_wb[4]_i_67 ,
    \rgf_c1bus_wb[4]_i_37 ,
    \sr[4]_i_240 ,
    \bbus_o[4]_INST_0_i_7 ,
    \bbus_o[4]_INST_0_i_7_0 ,
    \bbus_o[3]_INST_0_i_7 ,
    \bbus_o[3]_INST_0_i_7_0 ,
    \bbus_o[2]_INST_0_i_7 ,
    \bbus_o[2]_INST_0_i_7_0 ,
    \bbus_o[1]_INST_0_i_7 ,
    \bbus_o[1]_INST_0_i_7_0 ,
    \bbus_o[0]_INST_0_i_7 ,
    \bbus_o[0]_INST_0_i_7_0 ,
    \bbus_o[4]_INST_0_i_7_1 ,
    \bbus_o[4]_INST_0_i_7_2 ,
    \bbus_o[3]_INST_0_i_7_1 ,
    \bbus_o[3]_INST_0_i_7_2 ,
    \bbus_o[2]_INST_0_i_7_1 ,
    \bbus_o[2]_INST_0_i_7_2 ,
    \bbus_o[1]_INST_0_i_7_1 ,
    \bbus_o[1]_INST_0_i_7_2 ,
    \bbus_o[0]_INST_0_i_7_1 ,
    \bbus_o[0]_INST_0_i_7_2 ,
    \i_/bbus_o[4]_INST_0_i_20 ,
    \i_/bbus_o[4]_INST_0_i_20_0 ,
    \rgf_c1bus_wb[4]_i_40 ,
    \rgf_c1bus_wb[4]_i_42 ,
    \rgf_c1bus_wb[4]_i_50 ,
    \rgf_c1bus_wb[4]_i_48 ,
    \rgf_c1bus_wb[4]_i_64 ,
    \rgf_c1bus_wb[4]_i_62 ,
    \rgf_c1bus_wb[4]_i_60 ,
    \rgf_c1bus_wb[4]_i_58 ,
    \rgf_c1bus_wb[4]_i_56 ,
    \rgf_c1bus_wb[4]_i_54 ,
    \rgf_c1bus_wb[4]_i_52 ,
    \rgf_c1bus_wb[4]_i_32 ,
    \rgf_c1bus_wb[4]_i_34 ,
    \rgf_c1bus_wb[4]_i_36 ,
    \rgf_c1bus_wb[4]_i_38 ,
    \sr[4]_i_239 ,
    \bbus_o[4]_INST_0_i_7_3 ,
    \bbus_o[4]_INST_0_i_7_4 ,
    \bbus_o[3]_INST_0_i_7_3 ,
    \bbus_o[3]_INST_0_i_7_4 ,
    \bbus_o[2]_INST_0_i_7_3 ,
    \bbus_o[2]_INST_0_i_7_4 ,
    \bbus_o[1]_INST_0_i_7_3 ,
    \bbus_o[1]_INST_0_i_7_4 ,
    \bbus_o[0]_INST_0_i_7_3 ,
    \bbus_o[0]_INST_0_i_7_4 ,
    \bbus_o[4]_INST_0_i_7_5 ,
    \bbus_o[4]_INST_0_i_7_6 ,
    \bbus_o[3]_INST_0_i_7_5 ,
    \bbus_o[3]_INST_0_i_7_6 ,
    \bbus_o[2]_INST_0_i_7_5 ,
    \bbus_o[2]_INST_0_i_7_6 ,
    \bbus_o[1]_INST_0_i_7_5 ,
    \bbus_o[1]_INST_0_i_7_6 ,
    \bbus_o[0]_INST_0_i_7_5 ,
    \bbus_o[0]_INST_0_i_7_6 ,
    \rgf_c1bus_wb[4]_i_45 ,
    \rgf_c1bus_wb[4]_i_42_0 ,
    \rgf_c1bus_wb[4]_i_50_0 ,
    \rgf_c1bus_wb[4]_i_48_0 ,
    \rgf_c1bus_wb[4]_i_64_0 ,
    \rgf_c1bus_wb[4]_i_62_0 ,
    \rgf_c1bus_wb[4]_i_60_0 ,
    \rgf_c1bus_wb[4]_i_58_0 ,
    \rgf_c1bus_wb[4]_i_56_0 ,
    \rgf_c1bus_wb[4]_i_54_0 ,
    \rgf_c1bus_wb[4]_i_52_0 ,
    \rgf_c1bus_wb[4]_i_32_0 ,
    \rgf_c1bus_wb[4]_i_34_0 ,
    \rgf_c1bus_wb[4]_i_36_0 ,
    \rgf_c1bus_wb[4]_i_38_0 ,
    \rgf_c1bus_wb[4]_i_44 ,
    \bdatw[12]_INST_0_i_42 ,
    \bdatw[12]_INST_0_i_42_0 ,
    \bdatw[11]_INST_0_i_44 ,
    \bdatw[11]_INST_0_i_44_0 ,
    \bdatw[10]_INST_0_i_43 ,
    \bdatw[10]_INST_0_i_43_0 ,
    \bdatw[9]_INST_0_i_42 ,
    \bdatw[9]_INST_0_i_42_0 ,
    \bdatw[8]_INST_0_i_43 ,
    \bdatw[8]_INST_0_i_43_0 ,
    \sr_reg[15]_2 ,
    \pc_reg[15]_2 ,
    \sp_reg[15]_1 ,
    \iv_reg[15]_1 ,
    \tr_reg[15]_2 ,
    \abus_o[15] ,
    \abus_o[14] ,
    \abus_o[13] ,
    \abus_o[12] ,
    \abus_o[11] ,
    \abus_o[10] ,
    \abus_o[9] ,
    \abus_o[8] ,
    \abus_o[7] ,
    \abus_o[6] ,
    \abus_o[5] ,
    \abus_o[4] ,
    \abus_o[3] ,
    \abus_o[2] ,
    \abus_o[1] ,
    \abus_o[0] ,
    a0bus_sel_cr,
    \rgf_c0bus_wb[4]_i_21 ,
    a1bus_sr,
    a1bus_sel_cr,
    \rgf_c1bus_wb[4]_i_22 ,
    b0bus_sr,
    b0bus_sel_cr,
    b1bus_sel_cr,
    b1bus_sr,
    \grn_reg[15]_2 ,
    \grn_reg[15]_3 ,
    \grn_reg[15]_4 ,
    \grn_reg[15]_5 ,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[15]_10 ,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 ,
    \grn_reg[15]_46 ,
    \grn_reg[15]_47 ,
    \grn_reg[15]_48 ,
    \grn_reg[15]_49 ,
    \grn_reg[15]_50 ,
    \grn_reg[15]_51 ,
    \grn_reg[15]_52 ,
    \grn_reg[15]_53 ,
    \grn_reg[15]_54 ,
    \grn_reg[15]_55 ,
    \grn_reg[15]_56 ,
    \grn_reg[15]_57 ,
    \grn_reg[15]_58 ,
    \grn_reg[15]_59 ,
    \grn_reg[15]_60 ,
    \grn_reg[15]_61 ,
    \grn_reg[15]_62 ,
    \grn_reg[15]_63 ,
    \grn_reg[15]_64 ,
    \grn_reg[15]_65 );
  output rgf_selc0_stat;
  output rgf_selc1_stat;
  output [14:0]out;
  output [15:0]\grn_reg[15] ;
  output [4:0]\grn_reg[4] ;
  output [4:0]\grn_reg[4]_0 ;
  output [4:0]\grn_reg[4]_1 ;
  output [4:0]\grn_reg[4]_2 ;
  output [4:0]\grn_reg[4]_3 ;
  output [15:0]\grn_reg[15]_0 ;
  output [4:0]\grn_reg[4]_4 ;
  output [4:0]\grn_reg[4]_5 ;
  output [4:0]\grn_reg[4]_6 ;
  output [4:0]\grn_reg[4]_7 ;
  output [15:0]\sr_reg[15] ;
  output [15:0]\pc_reg[15] ;
  output [0:0]\sp_reg[0] ;
  output [15:0]\iv_reg[15] ;
  output [15:0]\tr_reg[15] ;
  output \sr_reg[4] ;
  output \sr_reg[5] ;
  output \pc_reg[15]_0 ;
  output [2:0]D;
  output \pc_reg[14] ;
  output \pc_reg[13] ;
  output [0:0]SR;
  output [0:0]\sp_reg[1] ;
  output \sp_reg[15] ;
  output \sp_reg[1]_0 ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  output \sp_reg[5] ;
  output \sp_reg[6] ;
  output \sp_reg[7] ;
  output \sp_reg[8] ;
  output \sp_reg[9] ;
  output \sp_reg[10] ;
  output \sp_reg[11] ;
  output \sp_reg[12] ;
  output \sp_reg[13] ;
  output \sp_reg[14] ;
  output [1:0]bdatw;
  output \tr_reg[14] ;
  output \tr_reg[14]_0 ;
  output \stat_reg[1] ;
  output \tr_reg[13] ;
  output \tr_reg[13]_0 ;
  output \stat_reg[1]_0 ;
  output \tr_reg[12] ;
  output \tr_reg[11] ;
  output \tr_reg[10] ;
  output \tr_reg[9] ;
  output \tr_reg[8] ;
  output \stat_reg[1]_1 ;
  output \tr_reg[7] ;
  output \tr_reg[7]_0 ;
  output \stat_reg[2] ;
  output \tr_reg[6] ;
  output [15:0]a1bus_0;
  output \badr[6]_INST_0_i_1 ;
  output \tr_reg[6]_0 ;
  output \stat_reg[2]_0 ;
  output \tr_reg[5] ;
  output \badr[5]_INST_0_i_1 ;
  output \tr_reg[5]_0 ;
  output \rgf_c1bus_wb[13]_i_9 ;
  output \rgf_c1bus_wb[14]_i_30 ;
  output \sr_reg[6] ;
  output \badr[15]_INST_0_i_1 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[6]_1 ;
  output \badr[3]_INST_0_i_1 ;
  output \sr[4]_i_156 ;
  output \tr_reg[11]_0 ;
  output \tr_reg[13]_1 ;
  output \badr[15]_INST_0_i_1_0 ;
  output \badr[1]_INST_0_i_1 ;
  output \sr_reg[6]_2 ;
  output \badr[9]_INST_0_i_1 ;
  output \sr_reg[6]_3 ;
  output \rgf_c1bus_wb[15]_i_14 ;
  output \badr[10]_INST_0_i_1 ;
  output \badr[6]_INST_0_i_1_0 ;
  output \badr[2]_INST_0_i_1 ;
  output \rgf_c1bus_wb[11]_i_13 ;
  output \badr[10]_INST_0_i_1_0 ;
  output \badr[14]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_14_0 ;
  output \badr[3]_INST_0_i_1_0 ;
  output \badr[7]_INST_0_i_1 ;
  output \badr[15]_INST_0_i_1_1 ;
  output \sr_reg[6]_4 ;
  output \badr[6]_INST_0_i_1_1 ;
  output \sr_reg[6]_5 ;
  output \rgf_c1bus_wb[12]_i_20 ;
  output \rgf_c1bus_wb[11]_i_10 ;
  output \badr[15]_INST_0_i_1_2 ;
  output \rgf_c1bus_wb[14]_i_28 ;
  output \rgf_c1bus_wb[15]_i_14_1 ;
  output \rgf_c1bus_wb[14]_i_28_0 ;
  output \rgf_c1bus_wb[7]_i_4 ;
  output \badr[5]_INST_0_i_1_0 ;
  output \sr[4]_i_219 ;
  output \tr_reg[12]_0 ;
  output \rgf_c1bus_wb[11]_i_10_0 ;
  output \rgf_c1bus_wb[4]_i_9 ;
  output \badr[12]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_28_1 ;
  output \sr_reg[6]_6 ;
  output \badr[0]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_28_2 ;
  output \rgf_c1bus_wb[14]_i_28_3 ;
  output \rgf_c1bus_wb[9]_i_17 ;
  output \badr[10]_INST_0_i_1_1 ;
  output \rgf_c1bus_wb[14]_i_28_4 ;
  output \rgf_c1bus_wb[13]_i_16 ;
  output \rgf_c1bus_wb[14]_i_28_5 ;
  output \rgf_c1bus_wb[4]_i_9_0 ;
  output \sr_reg[6]_7 ;
  output \tr_reg[1] ;
  output \sr_reg[6]_8 ;
  output \tr_reg[14]_1 ;
  output \sr_reg[6]_9 ;
  output \sr_reg[6]_10 ;
  output \rgf_c1bus_wb[15]_i_14_2 ;
  output \badr[11]_INST_0_i_1 ;
  output \sr_reg[6]_11 ;
  output \sr_reg[6]_12 ;
  output \badr[2]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[15]_i_14_3 ;
  output \rgf_c1bus_wb[14]_i_28_6 ;
  output \badr[9]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[14]_i_28_7 ;
  output \rgf_c1bus_wb[14]_i_32 ;
  output \badr[13]_INST_0_i_1 ;
  output \badr[2]_INST_0_i_1_1 ;
  output \rgf_c1bus_wb[14]_i_32_0 ;
  output \sr_reg[6]_13 ;
  output \sr_reg[6]_14 ;
  output \badr[14]_INST_0_i_1_0 ;
  output \stat_reg[2]_1 ;
  output \sr_reg[6]_15 ;
  output \rgf_c1bus_wb[11]_i_10_1 ;
  output \rgf_c1bus_wb[1]_i_14 ;
  output \badr[6]_INST_0_i_1_2 ;
  output \rgf_c1bus_wb[11]_i_10_2 ;
  output \sr_reg[6]_16 ;
  output \sr_reg[6]_17 ;
  output \rgf_c1bus_wb[4]_i_28 ;
  output \tr_reg[12]_1 ;
  output \sr[4]_i_220 ;
  output \tr_reg[3] ;
  output \rgf_c1bus_wb[11]_i_10_3 ;
  output \rgf_c1bus_wb[11]_i_10_4 ;
  output \rgf_c1bus_wb[15]_i_27 ;
  output \sr_reg[6]_18 ;
  output [0:0]\grn_reg[15]_1 ;
  output \tr_reg[15]_0 ;
  output \sr_reg[15]_0 ;
  output \sp_reg[15]_0 ;
  output \tr_reg[1]_0 ;
  output \tr_reg[14]_2 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[2]_3 ;
  output \tr_reg[15]_1 ;
  output [4:0]\grn_reg[4]_8 ;
  output [4:0]\grn_reg[4]_9 ;
  output \tr_reg[12]_2 ;
  output \tr_reg[11]_1 ;
  output \tr_reg[10]_0 ;
  output \tr_reg[9]_0 ;
  output \tr_reg[8]_0 ;
  output \rgf_c0bus_wb[15]_i_18 ;
  output \rgf_c0bus_wb[11]_i_3 ;
  output [15:0]a0bus_0;
  output \rgf_c0bus_wb[11]_i_3_0 ;
  output \badr[6]_INST_0_i_2 ;
  output \sr[4]_i_133 ;
  output \rgf_c0bus_wb[4]_i_26 ;
  output \rgf_c0bus_wb[11]_i_9 ;
  output \sr[4]_i_200 ;
  output \sr[4]_i_195 ;
  output \rgf_c0bus_wb[11]_i_9_0 ;
  output \rgf_c0bus_wb[4]_i_32 ;
  output \rgf_c0bus_wb[13]_i_27 ;
  output \sr_reg[6]_19 ;
  output \rgf_c0bus_wb[11]_i_11 ;
  output \badr[5]_INST_0_i_2 ;
  output \badr[1]_INST_0_i_2 ;
  output \badr[13]_INST_0_i_2 ;
  output \badr[9]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_11_0 ;
  output \rgf_c0bus_wb[11]_i_22 ;
  output \badr[8]_INST_0_i_2 ;
  output \badr[3]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_9_1 ;
  output \badr[10]_INST_0_i_2 ;
  output \badr[6]_INST_0_i_2_0 ;
  output \badr[2]_INST_0_i_2 ;
  output \rgf_c0bus_wb[15]_i_25 ;
  output \rgf_c0bus_wb[11]_i_8 ;
  output \badr[4]_INST_0_i_2 ;
  output \rgf_c0bus_wb[0]_i_14 ;
  output \sr_reg[6]_20 ;
  output \sr_reg[6]_21 ;
  output \badr[10]_INST_0_i_2_0 ;
  output \badr[14]_INST_0_i_2 ;
  output \rgf_c0bus_wb[13]_i_29 ;
  output \badr[4]_INST_0_i_2_0 ;
  output \badr[12]_INST_0_i_2 ;
  output \badr[8]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[7]_i_7 ;
  output \rgf_c0bus_wb[7]_i_7_0 ;
  output \sr_reg[6]_22 ;
  output \sr_reg[6]_23 ;
  output \badr[14]_INST_0_i_2_0 ;
  output \sr_reg[6]_24 ;
  output \rgf_c0bus_wb[11]_i_11_1 ;
  output \badr[6]_INST_0_i_2_1 ;
  output \rgf_c0bus_wb[11]_i_11_2 ;
  output \badr[13]_INST_0_i_2_0 ;
  output \badr[5]_INST_0_i_2_0 ;
  output \badr[9]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[15]_i_26 ;
  output \sr_reg[6]_25 ;
  output \sp_reg[2]_0 ;
  output \rgf_c0bus_wb[13]_i_30 ;
  output \sr_reg[6]_26 ;
  output \sr_reg[6]_27 ;
  output \sp_reg[13]_0 ;
  output \sp_reg[11]_0 ;
  output \sr_reg[6]_28 ;
  output \rgf_c0bus_wb[4]_i_29 ;
  output \badr[3]_INST_0_i_2_0 ;
  output \sr_reg[6]_29 ;
  output \rgf_c0bus_wb[4]_i_33 ;
  output \rgf_c0bus_wb[4]_i_31 ;
  output \badr[11]_INST_0_i_2 ;
  output \badr[7]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_22_0 ;
  output \sr[4]_i_232 ;
  output \sp_reg[1]_1 ;
  output \badr[2]_INST_0_i_2_0 ;
  output \sr_reg[6]_30 ;
  output \rgf_c0bus_wb[12]_i_24 ;
  output \sp_reg[4]_0 ;
  output \sr_reg[14] ;
  output \sr_reg[6]_31 ;
  output \sr_reg[6]_32 ;
  output \rgf_c0bus_wb[10]_i_8 ;
  output \rgf_c0bus_wb[11]_i_9_2 ;
  output \badr[1]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[13]_i_28 ;
  output \sr_reg[6]_33 ;
  output \badr[14]_INST_0_i_2_1 ;
  output \rgf_c0bus_wb[8]_i_6 ;
  output \rgf_c0bus_wb[12]_i_25 ;
  output \sr_reg[6]_34 ;
  output \sr_reg[6]_35 ;
  output \sr_reg[6]_36 ;
  output \sr_reg[6]_37 ;
  output \badr[8]_INST_0_i_2_1 ;
  output \badr[12]_INST_0_i_2_0 ;
  output \sr_reg[6]_38 ;
  output \badr[15]_INST_0_i_2 ;
  output \sp_reg[0]_0 ;
  output \sr_reg[0] ;
  output \rgf_c0bus_wb[11]_i_3_1 ;
  output \sr_reg[6]_39 ;
  output [2:0]fadr;
  output fch_irq_req;
  output [15:0]badrx;
  output \sr_reg[4]_0 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[7] ;
  output \sr_reg[5]_1 ;
  output \sr_reg[6]_40 ;
  output \sr_reg[5]_2 ;
  output \sr_reg[6]_41 ;
  output irq_0;
  output \sr_reg[10] ;
  output \sr_reg[4]_1 ;
  output \fdatx[15] ;
  output [0:0]S;
  output [0:0]\pc_reg[1] ;
  output [2:0]\pc_reg[15]_1 ;
  output \rgf_c1bus_wb[7]_i_4_0 ;
  output \sr_reg[6]_42 ;
  output \rgf_c1bus_wb[11]_i_10_5 ;
  output \rgf_c0bus_wb[15]_i_6 ;
  output \rgf_c0bus_wb[15]_i_6_0 ;
  output \rgf_c0bus_wb[15]_i_6_1 ;
  output [0:0]bbus_o;
  output \rgf_c0bus_wb[11]_i_3_2 ;
  output \rgf_c0bus_wb[11]_i_9_3 ;
  output \rgf_c0bus_wb[11]_i_9_4 ;
  output \rgf_c0bus_wb[11]_i_3_3 ;
  output \sr_reg[5]_3 ;
  output \sr_reg[5]_4 ;
  output \sr_reg[5]_5 ;
  output [0:0]\fdat[15] ;
  output \sr_reg[0]_0 ;
  output [3:0]\badr[14]_INST_0_i_1_1 ;
  output [2:0]\badr[13]_INST_0_i_1_0 ;
  output [0:0]\badr[14]_INST_0_i_2_2 ;
  output [1:0]\badr[6]_INST_0_i_1_3 ;
  output [1:0]tout__1_carry__0_i_1__0;
  output [3:0]\badr[10]_INST_0_i_1_2 ;
  output [3:0]tout__1_carry__1_i_1__0;
  output [0:0]\sr_reg[0]_1 ;
  output [2:0]\rgf_selc0_rn_wb_reg[2] ;
  output [1:0]\rgf_selc0_wb_reg[1] ;
  output [2:0]\rgf_selc1_rn_wb_reg[2] ;
  output [1:0]\rgf_selc1_wb_reg[1] ;
  output [15:0]\rgf_c0bus_wb_reg[15] ;
  output [15:0]\rgf_c1bus_wb_reg[15] ;
  output [0:0]\grn_reg[0] ;
  output [0:0]\grn_reg[0]_0 ;
  output \sp_reg[4]_1 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[2]_1 ;
  output \sp_reg[1]_2 ;
  output \sp_reg[0]_1 ;
  output \tr_reg[0] ;
  output \tr_reg[1]_1 ;
  output \tr_reg[2] ;
  output \tr_reg[3]_0 ;
  output \tr_reg[4] ;
  output \iv_reg[15]_0 ;
  output \sr_reg[15]_1 ;
  output \sr_reg[4]_2 ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sr_reg[0]_2 ;
  output \tr_reg[0]_0 ;
  output \tr_reg[1]_2 ;
  output \tr_reg[2]_0 ;
  output \tr_reg[3]_1 ;
  output \tr_reg[4]_0 ;
  output \sp_reg[0]_2 ;
  output \sp_reg[1]_3 ;
  output \sp_reg[2]_2 ;
  output \sp_reg[3]_1 ;
  output \sp_reg[4]_2 ;
  output [4:0]b1bus_b02;
  input [0:0]E;
  input p_2_in;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0] ;
  input rgf_selc1_stat_reg;
  input \rgf_c1bus_wb_reg[0] ;
  input rst_n;
  input \sr_reg[5]_6 ;
  input \pc_reg[13]_0 ;
  input \sp_reg[14]_0 ;
  input \sp_reg[14]_1 ;
  input \bdatw[13] ;
  input \bdatw[13]_0 ;
  input \bdatw[13]_1 ;
  input \bdatw[14] ;
  input \bdatw[14]_0 ;
  input \bdatw[13]_2 ;
  input \bdatw[13]_3 ;
  input \bdatw[12] ;
  input \bdatw[12]_0 ;
  input \bdatw[11] ;
  input \bdatw[11]_0 ;
  input \bdatw[10] ;
  input \bdatw[10]_0 ;
  input \bdatw[9] ;
  input \bdatw[9]_0 ;
  input \bdatw[8] ;
  input \bdatw[8]_0 ;
  input \rgf_c1bus_wb[15]_i_19 ;
  input \rgf_c1bus_wb[15]_i_19_0 ;
  input \rgf_c1bus_wb_reg[5] ;
  input \sr[6]_i_15 ;
  input \rgf_c1bus_wb[5]_i_10 ;
  input \rgf_c1bus_wb[14]_i_11 ;
  input \rgf_c1bus_wb[14]_i_11_0 ;
  input tout__1_carry__0_i_7__0;
  input tout__1_carry__0_i_7__0_0;
  input \rgf_c1bus_wb_reg[5]_0 ;
  input \rgf_c1bus_wb_reg[5]_1 ;
  input \rgf_c1bus_wb_reg[7] ;
  input \sr[6]_i_11 ;
  input \sr[6]_i_11_0 ;
  input \sr[4]_i_27 ;
  input \sr[6]_i_11_1 ;
  input \sr[4]_i_30 ;
  input \rgf_c1bus_wb[12]_i_2 ;
  input \rgf_c1bus_wb_reg[3] ;
  input \sr[4]_i_38 ;
  input \rgf_c1bus_wb_reg[4] ;
  input \sr[4]_i_44 ;
  input \rgf_c1bus_wb_reg[10] ;
  input \sr[4]_i_84 ;
  input \bdatw[15] ;
  input \bdatw[15]_0 ;
  input \bdatw[14]_1 ;
  input \bdatw[14]_2 ;
  input \bdatw[13]_4 ;
  input \bdatw[13]_5 ;
  input \bdatw[12]_1 ;
  input \bdatw[12]_2 ;
  input \bdatw[11]_1 ;
  input \bdatw[11]_2 ;
  input \bdatw[10]_1 ;
  input \bdatw[10]_2 ;
  input \bdatw[9]_1 ;
  input \bdatw[9]_2 ;
  input \bdatw[8]_1 ;
  input \bdatw[8]_2 ;
  input \rgf_c0bus_wb_reg[7]_i_11 ;
  input \sr[4]_i_67 ;
  input \rgf_c0bus_wb[6]_i_11 ;
  input \rgf_c0bus_wb[14]_i_2 ;
  input \bbus_o[7] ;
  input \bbus_o[7]_0 ;
  input \bbus_o[6] ;
  input \bbus_o[6]_0 ;
  input \bbus_o[5] ;
  input \bbus_o[5]_0 ;
  input \sr[4]_i_15 ;
  input \sr[4]_i_15_0 ;
  input \sr[4]_i_15_1 ;
  input \rgf_c0bus_wb_reg[10] ;
  input \sr[4]_i_66 ;
  input \rgf_c0bus_wb_reg[10]_0 ;
  input \rgf_c0bus_wb_reg[10]_1 ;
  input \rgf_c0bus_wb[12]_i_2 ;
  input \sr[4]_i_55 ;
  input \rgf_c0bus_wb[13]_i_4 ;
  input \rgf_c0bus_wb[10]_i_4 ;
  input \rgf_c0bus_wb[3]_i_7 ;
  input \rgf_c0bus_wb[3]_i_7_0 ;
  input \sr[4]_i_129 ;
  input \rgf_c0bus_wb[15]_i_14 ;
  input [2:0]\pc0_reg[15] ;
  input \fadr[15] ;
  input [2:0]O;
  input \fadr[15]_0 ;
  input \pc0_reg[15]_0 ;
  input \pc0_reg[15]_1 ;
  input [4:0]\badr[15]_INST_0_i_208 ;
  input [3:0]\rgf_selc1_wb[1]_i_16 ;
  input irq;
  input [1:0]irq_lev;
  input [0:0]Q;
  input ctl_fetch1_fl_i_15;
  input [13:0]fdatx;
  input \ir0_id_fl[20]_i_4 ;
  input [13:0]fdat;
  input \nir_id_reg[20] ;
  input \bbus_o[5]_1 ;
  input [1:0]b0bus_sel_0;
  input [3:0]a1bus_sel_0;
  input tout__1_carry__2;
  input tout__1_carry__2_0;
  input tout__1_carry__2_1;
  input [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  input [1:0]\rgf_selc0_wb_reg[1]_0 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  input [1:0]\rgf_selc1_wb_reg[1]_0 ;
  input [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  input [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [3:0]a0bus_sel_0;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_43 ;
  input [0:0]ctl_sela0;
  input \i_/badr[15]_INST_0_i_43_0 ;
  input \i_/bdatw[15]_INST_0_i_9 ;
  input \i_/bdatw[15]_INST_0_i_9_0 ;
  input \i_/bdatw[15]_INST_0_i_9_1 ;
  input \i_/bdatw[15]_INST_0_i_9_2 ;
  input [0:0]ctl_selb0_0;
  input \i_/bdatw[15]_INST_0_i_24 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_77 ;
  input \i_/bdatw[15]_INST_0_i_9_3 ;
  input \i_/bdatw[15]_INST_0_i_24_0 ;
  input \i_/badr[15]_INST_0_i_19 ;
  input \i_/badr[15]_INST_0_i_19_0 ;
  input \i_/badr[15]_INST_0_i_19_1 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_113 ;
  input \i_/bdatw[15]_INST_0_i_44 ;
  input \i_/bdatw[15]_INST_0_i_112 ;
  input \i_/bdatw[15]_INST_0_i_112_0 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_112_1 ;
  input \rgf_c1bus_wb[4]_i_47 ;
  input \rgf_c1bus_wb[4]_i_41 ;
  input \rgf_c1bus_wb[4]_i_51 ;
  input \sr[4]_i_235 ;
  input \rgf_c1bus_wb[4]_i_65 ;
  input \sr[4]_i_237 ;
  input \rgf_c1bus_wb[4]_i_61 ;
  input \rgf_c1bus_wb[4]_i_57 ;
  input \sr[4]_i_245 ;
  input \rgf_c1bus_wb[4]_i_53 ;
  input \sr[4]_i_243 ;
  input \rgf_c1bus_wb[4]_i_33 ;
  input \rgf_c1bus_wb[4]_i_67 ;
  input \rgf_c1bus_wb[4]_i_37 ;
  input \sr[4]_i_240 ;
  input \bbus_o[4]_INST_0_i_7 ;
  input \bbus_o[4]_INST_0_i_7_0 ;
  input \bbus_o[3]_INST_0_i_7 ;
  input \bbus_o[3]_INST_0_i_7_0 ;
  input \bbus_o[2]_INST_0_i_7 ;
  input \bbus_o[2]_INST_0_i_7_0 ;
  input \bbus_o[1]_INST_0_i_7 ;
  input \bbus_o[1]_INST_0_i_7_0 ;
  input \bbus_o[0]_INST_0_i_7 ;
  input \bbus_o[0]_INST_0_i_7_0 ;
  input \bbus_o[4]_INST_0_i_7_1 ;
  input \bbus_o[4]_INST_0_i_7_2 ;
  input \bbus_o[3]_INST_0_i_7_1 ;
  input \bbus_o[3]_INST_0_i_7_2 ;
  input \bbus_o[2]_INST_0_i_7_1 ;
  input \bbus_o[2]_INST_0_i_7_2 ;
  input \bbus_o[1]_INST_0_i_7_1 ;
  input \bbus_o[1]_INST_0_i_7_2 ;
  input \bbus_o[0]_INST_0_i_7_1 ;
  input \bbus_o[0]_INST_0_i_7_2 ;
  input \i_/bbus_o[4]_INST_0_i_20 ;
  input \i_/bbus_o[4]_INST_0_i_20_0 ;
  input \rgf_c1bus_wb[4]_i_40 ;
  input \rgf_c1bus_wb[4]_i_42 ;
  input \rgf_c1bus_wb[4]_i_50 ;
  input \rgf_c1bus_wb[4]_i_48 ;
  input \rgf_c1bus_wb[4]_i_64 ;
  input \rgf_c1bus_wb[4]_i_62 ;
  input \rgf_c1bus_wb[4]_i_60 ;
  input \rgf_c1bus_wb[4]_i_58 ;
  input \rgf_c1bus_wb[4]_i_56 ;
  input \rgf_c1bus_wb[4]_i_54 ;
  input \rgf_c1bus_wb[4]_i_52 ;
  input \rgf_c1bus_wb[4]_i_32 ;
  input \rgf_c1bus_wb[4]_i_34 ;
  input \rgf_c1bus_wb[4]_i_36 ;
  input \rgf_c1bus_wb[4]_i_38 ;
  input \sr[4]_i_239 ;
  input \bbus_o[4]_INST_0_i_7_3 ;
  input \bbus_o[4]_INST_0_i_7_4 ;
  input \bbus_o[3]_INST_0_i_7_3 ;
  input \bbus_o[3]_INST_0_i_7_4 ;
  input \bbus_o[2]_INST_0_i_7_3 ;
  input \bbus_o[2]_INST_0_i_7_4 ;
  input \bbus_o[1]_INST_0_i_7_3 ;
  input \bbus_o[1]_INST_0_i_7_4 ;
  input \bbus_o[0]_INST_0_i_7_3 ;
  input \bbus_o[0]_INST_0_i_7_4 ;
  input \bbus_o[4]_INST_0_i_7_5 ;
  input \bbus_o[4]_INST_0_i_7_6 ;
  input \bbus_o[3]_INST_0_i_7_5 ;
  input \bbus_o[3]_INST_0_i_7_6 ;
  input \bbus_o[2]_INST_0_i_7_5 ;
  input \bbus_o[2]_INST_0_i_7_6 ;
  input \bbus_o[1]_INST_0_i_7_5 ;
  input \bbus_o[1]_INST_0_i_7_6 ;
  input \bbus_o[0]_INST_0_i_7_5 ;
  input \bbus_o[0]_INST_0_i_7_6 ;
  input \rgf_c1bus_wb[4]_i_45 ;
  input \rgf_c1bus_wb[4]_i_42_0 ;
  input \rgf_c1bus_wb[4]_i_50_0 ;
  input \rgf_c1bus_wb[4]_i_48_0 ;
  input \rgf_c1bus_wb[4]_i_64_0 ;
  input \rgf_c1bus_wb[4]_i_62_0 ;
  input \rgf_c1bus_wb[4]_i_60_0 ;
  input \rgf_c1bus_wb[4]_i_58_0 ;
  input \rgf_c1bus_wb[4]_i_56_0 ;
  input \rgf_c1bus_wb[4]_i_54_0 ;
  input \rgf_c1bus_wb[4]_i_52_0 ;
  input \rgf_c1bus_wb[4]_i_32_0 ;
  input \rgf_c1bus_wb[4]_i_34_0 ;
  input \rgf_c1bus_wb[4]_i_36_0 ;
  input \rgf_c1bus_wb[4]_i_38_0 ;
  input \rgf_c1bus_wb[4]_i_44 ;
  input \bdatw[12]_INST_0_i_42 ;
  input \bdatw[12]_INST_0_i_42_0 ;
  input \bdatw[11]_INST_0_i_44 ;
  input \bdatw[11]_INST_0_i_44_0 ;
  input \bdatw[10]_INST_0_i_43 ;
  input \bdatw[10]_INST_0_i_43_0 ;
  input \bdatw[9]_INST_0_i_42 ;
  input \bdatw[9]_INST_0_i_42_0 ;
  input \bdatw[8]_INST_0_i_43 ;
  input \bdatw[8]_INST_0_i_43_0 ;
  input [15:0]\sr_reg[15]_2 ;
  input [15:0]\pc_reg[15]_2 ;
  input [15:0]\sp_reg[15]_1 ;
  input [15:0]\iv_reg[15]_1 ;
  input [15:0]\tr_reg[15]_2 ;
  input \abus_o[15] ;
  input \abus_o[14] ;
  input \abus_o[13] ;
  input \abus_o[12] ;
  input \abus_o[11] ;
  input \abus_o[10] ;
  input \abus_o[9] ;
  input \abus_o[8] ;
  input \abus_o[7] ;
  input \abus_o[6] ;
  input \abus_o[5] ;
  input \abus_o[4] ;
  input \abus_o[3] ;
  input \abus_o[2] ;
  input \abus_o[1] ;
  input \abus_o[0] ;
  input [3:0]a0bus_sel_cr;
  input [15:0]\rgf_c0bus_wb[4]_i_21 ;
  input [15:0]a1bus_sr;
  input [4:0]a1bus_sel_cr;
  input [15:0]\rgf_c1bus_wb[4]_i_22 ;
  input [15:0]b0bus_sr;
  input [4:0]b0bus_sel_cr;
  input [5:0]b1bus_sel_cr;
  input [14:0]b1bus_sr;
  input [0:0]\grn_reg[15]_2 ;
  input [15:0]\grn_reg[15]_3 ;
  input [0:0]\grn_reg[15]_4 ;
  input [15:0]\grn_reg[15]_5 ;
  input [0:0]\grn_reg[15]_6 ;
  input [15:0]\grn_reg[15]_7 ;
  input [0:0]\grn_reg[15]_8 ;
  input [15:0]\grn_reg[15]_9 ;
  input [0:0]\grn_reg[15]_10 ;
  input [15:0]\grn_reg[15]_11 ;
  input [0:0]\grn_reg[15]_12 ;
  input [15:0]\grn_reg[15]_13 ;
  input [0:0]\grn_reg[15]_14 ;
  input [15:0]\grn_reg[15]_15 ;
  input [0:0]\grn_reg[15]_16 ;
  input [15:0]\grn_reg[15]_17 ;
  input [0:0]\grn_reg[15]_18 ;
  input [15:0]\grn_reg[15]_19 ;
  input [0:0]\grn_reg[15]_20 ;
  input [15:0]\grn_reg[15]_21 ;
  input [0:0]\grn_reg[15]_22 ;
  input [15:0]\grn_reg[15]_23 ;
  input [0:0]\grn_reg[15]_24 ;
  input [15:0]\grn_reg[15]_25 ;
  input [0:0]\grn_reg[15]_26 ;
  input [15:0]\grn_reg[15]_27 ;
  input [0:0]\grn_reg[15]_28 ;
  input [15:0]\grn_reg[15]_29 ;
  input [0:0]\grn_reg[15]_30 ;
  input [15:0]\grn_reg[15]_31 ;
  input [0:0]\grn_reg[15]_32 ;
  input [15:0]\grn_reg[15]_33 ;
  input [0:0]\grn_reg[15]_34 ;
  input [15:0]\grn_reg[15]_35 ;
  input [0:0]\grn_reg[15]_36 ;
  input [15:0]\grn_reg[15]_37 ;
  input [0:0]\grn_reg[15]_38 ;
  input [15:0]\grn_reg[15]_39 ;
  input [0:0]\grn_reg[15]_40 ;
  input [15:0]\grn_reg[15]_41 ;
  input [0:0]\grn_reg[15]_42 ;
  input [15:0]\grn_reg[15]_43 ;
  input [0:0]\grn_reg[15]_44 ;
  input [15:0]\grn_reg[15]_45 ;
  input [0:0]\grn_reg[15]_46 ;
  input [15:0]\grn_reg[15]_47 ;
  input [0:0]\grn_reg[15]_48 ;
  input [15:0]\grn_reg[15]_49 ;
  input [0:0]\grn_reg[15]_50 ;
  input [15:0]\grn_reg[15]_51 ;
  input [0:0]\grn_reg[15]_52 ;
  input [15:0]\grn_reg[15]_53 ;
  input [0:0]\grn_reg[15]_54 ;
  input [15:0]\grn_reg[15]_55 ;
  input [0:0]\grn_reg[15]_56 ;
  input [15:0]\grn_reg[15]_57 ;
  input [0:0]\grn_reg[15]_58 ;
  input [15:0]\grn_reg[15]_59 ;
  input [0:0]\grn_reg[15]_60 ;
  input [15:0]\grn_reg[15]_61 ;
  input [0:0]\grn_reg[15]_62 ;
  input [15:0]\grn_reg[15]_63 ;
  input [0:0]\grn_reg[15]_64 ;
  input [15:0]\grn_reg[15]_65 ;
  output fdat_12_sn_1;
  input badrx_15_sn_1;

  wire [2:0]D;
  wire [0:0]E;
  wire [2:0]O;
  wire [0:0]Q;
  wire [0:0]S;
  wire [0:0]SR;
  wire [15:0]a0bus_0;
  wire a0bus_out_n_1;
  wire a0bus_out_n_10;
  wire a0bus_out_n_11;
  wire a0bus_out_n_13;
  wire a0bus_out_n_14;
  wire a0bus_out_n_15;
  wire a0bus_out_n_17;
  wire a0bus_out_n_18;
  wire a0bus_out_n_19;
  wire a0bus_out_n_2;
  wire a0bus_out_n_21;
  wire a0bus_out_n_22;
  wire a0bus_out_n_23;
  wire a0bus_out_n_25;
  wire a0bus_out_n_26;
  wire a0bus_out_n_27;
  wire a0bus_out_n_29;
  wire a0bus_out_n_3;
  wire a0bus_out_n_30;
  wire a0bus_out_n_31;
  wire a0bus_out_n_33;
  wire a0bus_out_n_34;
  wire a0bus_out_n_35;
  wire a0bus_out_n_37;
  wire a0bus_out_n_38;
  wire a0bus_out_n_39;
  wire a0bus_out_n_41;
  wire a0bus_out_n_42;
  wire a0bus_out_n_43;
  wire a0bus_out_n_45;
  wire a0bus_out_n_46;
  wire a0bus_out_n_47;
  wire a0bus_out_n_49;
  wire a0bus_out_n_5;
  wire a0bus_out_n_50;
  wire a0bus_out_n_51;
  wire a0bus_out_n_53;
  wire a0bus_out_n_54;
  wire a0bus_out_n_55;
  wire a0bus_out_n_57;
  wire a0bus_out_n_58;
  wire a0bus_out_n_59;
  wire a0bus_out_n_6;
  wire a0bus_out_n_63;
  wire a0bus_out_n_64;
  wire a0bus_out_n_65;
  wire a0bus_out_n_66;
  wire a0bus_out_n_67;
  wire a0bus_out_n_68;
  wire a0bus_out_n_69;
  wire a0bus_out_n_7;
  wire a0bus_out_n_70;
  wire a0bus_out_n_71;
  wire a0bus_out_n_72;
  wire a0bus_out_n_73;
  wire a0bus_out_n_74;
  wire a0bus_out_n_75;
  wire a0bus_out_n_76;
  wire a0bus_out_n_77;
  wire a0bus_out_n_78;
  wire a0bus_out_n_79;
  wire a0bus_out_n_9;
  wire [3:0]a0bus_sel_0;
  wire [3:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [14:0]a1bus_b02;
  wire [15:0]a1bus_b13;
  wire a1bus_out_n_11;
  wire a1bus_out_n_12;
  wire a1bus_out_n_14;
  wire a1bus_out_n_15;
  wire a1bus_out_n_17;
  wire a1bus_out_n_18;
  wire a1bus_out_n_20;
  wire a1bus_out_n_21;
  wire a1bus_out_n_23;
  wire a1bus_out_n_25;
  wire a1bus_out_n_26;
  wire a1bus_out_n_28;
  wire a1bus_out_n_29;
  wire a1bus_out_n_3;
  wire a1bus_out_n_31;
  wire a1bus_out_n_32;
  wire a1bus_out_n_34;
  wire a1bus_out_n_35;
  wire a1bus_out_n_37;
  wire a1bus_out_n_38;
  wire a1bus_out_n_40;
  wire a1bus_out_n_41;
  wire a1bus_out_n_43;
  wire a1bus_out_n_44;
  wire a1bus_out_n_46;
  wire a1bus_out_n_47;
  wire a1bus_out_n_48;
  wire a1bus_out_n_49;
  wire a1bus_out_n_5;
  wire a1bus_out_n_51;
  wire a1bus_out_n_52;
  wire a1bus_out_n_53;
  wire a1bus_out_n_54;
  wire a1bus_out_n_55;
  wire a1bus_out_n_56;
  wire a1bus_out_n_57;
  wire a1bus_out_n_58;
  wire a1bus_out_n_59;
  wire a1bus_out_n_6;
  wire a1bus_out_n_60;
  wire a1bus_out_n_61;
  wire a1bus_out_n_62;
  wire a1bus_out_n_63;
  wire a1bus_out_n_64;
  wire a1bus_out_n_65;
  wire a1bus_out_n_66;
  wire a1bus_out_n_8;
  wire a1bus_out_n_9;
  wire [3:0]a1bus_sel_0;
  wire [4:0]a1bus_sel_cr;
  wire [15:0]a1bus_sr;
  wire \a1buso/gr6_bus1 ;
  wire \a1buso2l/gr6_bus1 ;
  wire \a1buso2l/gr6_bus1_0 ;
  wire \abus_o[0] ;
  wire \abus_o[10] ;
  wire \abus_o[11] ;
  wire \abus_o[12] ;
  wire \abus_o[13] ;
  wire \abus_o[14] ;
  wire \abus_o[15] ;
  wire \abus_o[1] ;
  wire \abus_o[2] ;
  wire \abus_o[3] ;
  wire \abus_o[4] ;
  wire \abus_o[5] ;
  wire \abus_o[6] ;
  wire \abus_o[7] ;
  wire \abus_o[8] ;
  wire \abus_o[9] ;
  wire b0bus_out_n_0;
  wire b0bus_out_n_1;
  wire b0bus_out_n_10;
  wire b0bus_out_n_2;
  wire b0bus_out_n_21;
  wire b0bus_out_n_22;
  wire b0bus_out_n_23;
  wire b0bus_out_n_24;
  wire b0bus_out_n_25;
  wire b0bus_out_n_26;
  wire b0bus_out_n_27;
  wire b0bus_out_n_28;
  wire b0bus_out_n_29;
  wire b0bus_out_n_3;
  wire b0bus_out_n_30;
  wire b0bus_out_n_31;
  wire b0bus_out_n_4;
  wire b0bus_out_n_5;
  wire b0bus_out_n_6;
  wire b0bus_out_n_7;
  wire b0bus_out_n_8;
  wire b0bus_out_n_9;
  wire [1:0]b0bus_sel_0;
  wire [4:0]b0bus_sel_cr;
  wire [15:0]b0bus_sr;
  wire [4:0]b1bus_b02;
  wire b1bus_out_n_10;
  wire b1bus_out_n_11;
  wire b1bus_out_n_2;
  wire b1bus_out_n_22;
  wire b1bus_out_n_23;
  wire b1bus_out_n_24;
  wire b1bus_out_n_25;
  wire b1bus_out_n_26;
  wire b1bus_out_n_27;
  wire b1bus_out_n_28;
  wire b1bus_out_n_29;
  wire b1bus_out_n_3;
  wire b1bus_out_n_30;
  wire b1bus_out_n_31;
  wire b1bus_out_n_4;
  wire b1bus_out_n_5;
  wire b1bus_out_n_6;
  wire b1bus_out_n_7;
  wire b1bus_out_n_8;
  wire b1bus_out_n_9;
  wire [5:0]b1bus_sel_cr;
  wire [14:0]b1bus_sr;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1_0 ;
  wire \badr[10]_INST_0_i_1_1 ;
  wire [3:0]\badr[10]_INST_0_i_1_2 ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[10]_INST_0_i_2_0 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2_0 ;
  wire \badr[13]_INST_0_i_1 ;
  wire [2:0]\badr[13]_INST_0_i_1_0 ;
  wire \badr[13]_INST_0_i_2 ;
  wire \badr[13]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire [3:0]\badr[14]_INST_0_i_1_1 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_2_1 ;
  wire [0:0]\badr[14]_INST_0_i_2_2 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_1_1 ;
  wire \badr[15]_INST_0_i_1_2 ;
  wire \badr[15]_INST_0_i_2 ;
  wire [4:0]\badr[15]_INST_0_i_208 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2_0 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1_0 ;
  wire \badr[2]_INST_0_i_1_1 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2_0 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1_0 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[3]_INST_0_i_2_0 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_2_0 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_2_0 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1_0 ;
  wire \badr[6]_INST_0_i_1_1 ;
  wire \badr[6]_INST_0_i_1_2 ;
  wire [1:0]\badr[6]_INST_0_i_1_3 ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2_0 ;
  wire \badr[6]_INST_0_i_2_1 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2_0 ;
  wire \badr[8]_INST_0_i_2_1 ;
  wire \badr[9]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1_0 ;
  wire \badr[9]_INST_0_i_2 ;
  wire \badr[9]_INST_0_i_2_0 ;
  wire [15:0]badrx;
  wire badrx_15_sn_1;
  wire bank02_n_15;
  wire bank02_n_16;
  wire bank02_n_17;
  wire bank02_n_18;
  wire bank02_n_19;
  wire bank02_n_20;
  wire bank02_n_21;
  wire bank02_n_22;
  wire bank02_n_23;
  wire bank02_n_24;
  wire bank02_n_25;
  wire bank02_n_26;
  wire bank02_n_264;
  wire bank02_n_27;
  wire bank02_n_28;
  wire bank02_n_281;
  wire bank02_n_29;
  wire bank02_n_30;
  wire bank02_n_31;
  wire bank02_n_32;
  wire bank02_n_33;
  wire bank02_n_330;
  wire bank02_n_331;
  wire bank02_n_332;
  wire bank02_n_333;
  wire bank02_n_334;
  wire bank02_n_335;
  wire bank02_n_336;
  wire bank02_n_337;
  wire bank02_n_338;
  wire bank02_n_339;
  wire bank02_n_34;
  wire bank02_n_340;
  wire bank02_n_341;
  wire bank02_n_342;
  wire bank02_n_343;
  wire bank02_n_344;
  wire bank02_n_345;
  wire bank02_n_346;
  wire bank02_n_347;
  wire bank02_n_348;
  wire bank02_n_349;
  wire bank02_n_35;
  wire bank02_n_350;
  wire bank02_n_351;
  wire bank02_n_352;
  wire bank02_n_353;
  wire bank02_n_354;
  wire bank02_n_355;
  wire bank02_n_356;
  wire bank02_n_357;
  wire bank02_n_358;
  wire bank02_n_359;
  wire bank02_n_36;
  wire bank02_n_361;
  wire bank02_n_362;
  wire bank02_n_37;
  wire bank02_n_38;
  wire bank02_n_384;
  wire bank02_n_385;
  wire bank02_n_386;
  wire bank02_n_387;
  wire bank02_n_388;
  wire bank02_n_389;
  wire bank02_n_39;
  wire bank02_n_390;
  wire bank02_n_391;
  wire bank02_n_392;
  wire bank02_n_393;
  wire bank02_n_394;
  wire bank02_n_395;
  wire bank02_n_396;
  wire bank02_n_397;
  wire bank02_n_398;
  wire bank02_n_399;
  wire bank02_n_40;
  wire bank02_n_400;
  wire bank02_n_401;
  wire bank02_n_402;
  wire bank02_n_403;
  wire bank02_n_404;
  wire bank02_n_405;
  wire bank02_n_406;
  wire bank02_n_407;
  wire bank02_n_408;
  wire bank02_n_409;
  wire bank02_n_41;
  wire bank02_n_410;
  wire bank02_n_411;
  wire bank02_n_412;
  wire bank02_n_413;
  wire bank02_n_414;
  wire bank02_n_42;
  wire bank02_n_43;
  wire bank02_n_430;
  wire bank02_n_431;
  wire bank02_n_432;
  wire bank02_n_433;
  wire bank02_n_434;
  wire bank02_n_435;
  wire bank02_n_436;
  wire bank02_n_437;
  wire bank02_n_438;
  wire bank02_n_439;
  wire bank02_n_44;
  wire bank02_n_440;
  wire bank02_n_441;
  wire bank02_n_442;
  wire bank02_n_443;
  wire bank02_n_444;
  wire bank02_n_446;
  wire bank02_n_447;
  wire bank02_n_448;
  wire bank02_n_449;
  wire bank02_n_45;
  wire bank02_n_450;
  wire bank02_n_451;
  wire bank02_n_452;
  wire bank02_n_453;
  wire bank02_n_454;
  wire bank02_n_455;
  wire bank02_n_456;
  wire bank02_n_457;
  wire bank02_n_458;
  wire bank02_n_459;
  wire bank02_n_46;
  wire bank02_n_460;
  wire bank02_n_461;
  wire bank02_n_462;
  wire bank02_n_47;
  wire bank02_n_48;
  wire bank02_n_484;
  wire bank02_n_485;
  wire bank02_n_486;
  wire bank02_n_487;
  wire bank02_n_488;
  wire bank02_n_489;
  wire bank02_n_49;
  wire bank02_n_490;
  wire bank02_n_491;
  wire bank02_n_492;
  wire bank02_n_493;
  wire bank02_n_494;
  wire bank02_n_495;
  wire bank02_n_496;
  wire bank02_n_497;
  wire bank02_n_498;
  wire bank02_n_499;
  wire bank02_n_50;
  wire bank02_n_501;
  wire bank02_n_502;
  wire bank02_n_503;
  wire bank02_n_504;
  wire bank02_n_505;
  wire bank02_n_506;
  wire bank02_n_507;
  wire bank02_n_508;
  wire bank02_n_509;
  wire bank02_n_51;
  wire bank02_n_510;
  wire bank02_n_511;
  wire bank02_n_512;
  wire bank02_n_513;
  wire bank02_n_514;
  wire bank02_n_515;
  wire bank02_n_52;
  wire bank02_n_53;
  wire bank02_n_54;
  wire bank02_n_55;
  wire bank02_n_56;
  wire bank02_n_57;
  wire bank02_n_58;
  wire bank02_n_59;
  wire bank02_n_60;
  wire bank02_n_61;
  wire bank02_n_62;
  wire bank02_n_63;
  wire bank02_n_64;
  wire bank02_n_65;
  wire bank02_n_66;
  wire bank02_n_67;
  wire bank02_n_68;
  wire bank02_n_69;
  wire bank02_n_70;
  wire bank02_n_71;
  wire bank02_n_72;
  wire bank02_n_73;
  wire bank02_n_74;
  wire bank02_n_75;
  wire bank02_n_76;
  wire bank02_n_77;
  wire bank02_n_78;
  wire bank02_n_79;
  wire bank02_n_80;
  wire bank02_n_81;
  wire bank02_n_82;
  wire bank02_n_83;
  wire bank02_n_84;
  wire bank02_n_85;
  wire bank02_n_86;
  wire bank02_n_87;
  wire bank02_n_88;
  wire bank13_n_105;
  wire bank13_n_106;
  wire bank13_n_107;
  wire bank13_n_108;
  wire bank13_n_109;
  wire bank13_n_110;
  wire bank13_n_111;
  wire bank13_n_112;
  wire bank13_n_113;
  wire bank13_n_114;
  wire bank13_n_115;
  wire bank13_n_116;
  wire bank13_n_117;
  wire bank13_n_118;
  wire bank13_n_119;
  wire bank13_n_120;
  wire bank13_n_130;
  wire bank13_n_138;
  wire bank13_n_156;
  wire bank13_n_164;
  wire bank13_n_168;
  wire bank13_n_169;
  wire bank13_n_170;
  wire bank13_n_171;
  wire bank13_n_172;
  wire bank13_n_173;
  wire bank13_n_174;
  wire bank13_n_175;
  wire bank13_n_176;
  wire bank13_n_177;
  wire bank13_n_178;
  wire bank13_n_179;
  wire bank13_n_180;
  wire bank13_n_181;
  wire bank13_n_182;
  wire bank13_n_183;
  wire bank13_n_184;
  wire bank13_n_185;
  wire bank13_n_186;
  wire bank13_n_187;
  wire bank13_n_188;
  wire bank13_n_189;
  wire bank13_n_190;
  wire bank13_n_191;
  wire bank13_n_192;
  wire bank13_n_193;
  wire bank13_n_194;
  wire bank13_n_195;
  wire bank13_n_196;
  wire bank13_n_197;
  wire bank13_n_198;
  wire bank13_n_199;
  wire bank13_n_200;
  wire bank13_n_201;
  wire bank13_n_202;
  wire bank13_n_203;
  wire bank13_n_204;
  wire bank13_n_205;
  wire bank13_n_206;
  wire bank13_n_207;
  wire bank13_n_208;
  wire bank13_n_209;
  wire bank13_n_210;
  wire bank13_n_211;
  wire bank13_n_212;
  wire bank13_n_213;
  wire bank13_n_214;
  wire bank13_n_215;
  wire bank13_n_216;
  wire bank13_n_217;
  wire bank13_n_218;
  wire bank13_n_219;
  wire bank13_n_220;
  wire bank13_n_221;
  wire bank13_n_222;
  wire bank13_n_223;
  wire bank13_n_224;
  wire bank13_n_225;
  wire bank13_n_226;
  wire bank13_n_227;
  wire bank13_n_228;
  wire bank13_n_229;
  wire bank13_n_230;
  wire bank13_n_231;
  wire bank13_n_232;
  wire bank13_n_233;
  wire bank13_n_234;
  wire bank13_n_235;
  wire bank13_n_236;
  wire bank13_n_237;
  wire bank13_n_238;
  wire bank13_n_239;
  wire bank13_n_240;
  wire bank13_n_241;
  wire bank13_n_242;
  wire bank13_n_243;
  wire bank13_n_244;
  wire bank13_n_245;
  wire bank13_n_246;
  wire bank13_n_247;
  wire bank13_n_248;
  wire bank13_n_250;
  wire bank13_n_251;
  wire bank13_n_252;
  wire bank13_n_253;
  wire bank13_n_254;
  wire bank13_n_255;
  wire bank13_n_256;
  wire bank13_n_257;
  wire bank13_n_258;
  wire bank13_n_259;
  wire bank13_n_26;
  wire bank13_n_260;
  wire bank13_n_261;
  wire bank13_n_262;
  wire bank13_n_263;
  wire bank13_n_264;
  wire bank13_n_265;
  wire bank13_n_266;
  wire bank13_n_267;
  wire bank13_n_268;
  wire bank13_n_269;
  wire bank13_n_27;
  wire bank13_n_270;
  wire bank13_n_271;
  wire bank13_n_272;
  wire bank13_n_273;
  wire bank13_n_274;
  wire bank13_n_275;
  wire bank13_n_276;
  wire bank13_n_277;
  wire bank13_n_278;
  wire bank13_n_279;
  wire bank13_n_28;
  wire bank13_n_280;
  wire bank13_n_281;
  wire bank13_n_282;
  wire bank13_n_283;
  wire bank13_n_284;
  wire bank13_n_285;
  wire bank13_n_286;
  wire bank13_n_287;
  wire bank13_n_288;
  wire bank13_n_289;
  wire bank13_n_29;
  wire bank13_n_290;
  wire bank13_n_291;
  wire bank13_n_292;
  wire bank13_n_293;
  wire bank13_n_294;
  wire bank13_n_295;
  wire bank13_n_296;
  wire bank13_n_297;
  wire bank13_n_298;
  wire bank13_n_299;
  wire bank13_n_30;
  wire bank13_n_300;
  wire bank13_n_301;
  wire bank13_n_302;
  wire bank13_n_31;
  wire bank13_n_319;
  wire bank13_n_32;
  wire bank13_n_320;
  wire bank13_n_321;
  wire bank13_n_322;
  wire bank13_n_323;
  wire bank13_n_324;
  wire bank13_n_325;
  wire bank13_n_326;
  wire bank13_n_327;
  wire bank13_n_328;
  wire bank13_n_329;
  wire bank13_n_33;
  wire bank13_n_330;
  wire bank13_n_331;
  wire bank13_n_332;
  wire bank13_n_333;
  wire bank13_n_334;
  wire bank13_n_335;
  wire bank13_n_336;
  wire bank13_n_337;
  wire bank13_n_338;
  wire bank13_n_339;
  wire bank13_n_34;
  wire bank13_n_340;
  wire bank13_n_341;
  wire bank13_n_342;
  wire bank13_n_343;
  wire bank13_n_344;
  wire bank13_n_345;
  wire bank13_n_346;
  wire bank13_n_347;
  wire bank13_n_348;
  wire bank13_n_349;
  wire bank13_n_35;
  wire bank13_n_350;
  wire bank13_n_351;
  wire bank13_n_352;
  wire bank13_n_353;
  wire bank13_n_354;
  wire bank13_n_355;
  wire bank13_n_356;
  wire bank13_n_357;
  wire bank13_n_358;
  wire bank13_n_359;
  wire bank13_n_36;
  wire bank13_n_360;
  wire bank13_n_361;
  wire bank13_n_362;
  wire bank13_n_363;
  wire bank13_n_364;
  wire bank13_n_365;
  wire bank13_n_366;
  wire bank13_n_367;
  wire bank13_n_368;
  wire bank13_n_369;
  wire bank13_n_370;
  wire bank13_n_371;
  wire bank13_n_372;
  wire bank13_n_373;
  wire bank13_n_374;
  wire bank13_n_375;
  wire bank13_n_376;
  wire bank13_n_377;
  wire bank13_n_378;
  wire bank13_n_379;
  wire bank13_n_380;
  wire bank13_n_381;
  wire bank13_n_382;
  wire bank13_n_383;
  wire bank13_n_385;
  wire bank13_n_386;
  wire bank13_n_387;
  wire bank13_n_388;
  wire bank13_n_389;
  wire bank13_n_390;
  wire bank13_n_391;
  wire bank13_n_392;
  wire bank13_n_393;
  wire bank13_n_394;
  wire bank13_n_395;
  wire bank13_n_396;
  wire bank13_n_397;
  wire bank13_n_398;
  wire bank13_n_399;
  wire bank13_n_400;
  wire bank13_n_401;
  wire bank13_n_402;
  wire bank13_n_403;
  wire bank13_n_404;
  wire bank13_n_405;
  wire bank13_n_406;
  wire bank13_n_407;
  wire bank13_n_408;
  wire bank13_n_409;
  wire bank13_n_410;
  wire bank13_n_411;
  wire bank13_n_412;
  wire bank13_n_413;
  wire bank13_n_414;
  wire bank13_n_415;
  wire bank13_n_416;
  wire bank13_n_417;
  wire bank13_n_418;
  wire bank13_n_419;
  wire bank13_n_42;
  wire bank13_n_420;
  wire bank13_n_421;
  wire bank13_n_422;
  wire bank13_n_423;
  wire bank13_n_424;
  wire bank13_n_425;
  wire bank13_n_426;
  wire bank13_n_427;
  wire bank13_n_428;
  wire bank13_n_429;
  wire bank13_n_43;
  wire bank13_n_430;
  wire bank13_n_431;
  wire bank13_n_432;
  wire bank13_n_433;
  wire bank13_n_434;
  wire bank13_n_435;
  wire bank13_n_436;
  wire bank13_n_437;
  wire bank13_n_438;
  wire bank13_n_439;
  wire bank13_n_44;
  wire bank13_n_440;
  wire bank13_n_441;
  wire bank13_n_442;
  wire bank13_n_443;
  wire bank13_n_444;
  wire bank13_n_445;
  wire bank13_n_446;
  wire bank13_n_45;
  wire bank13_n_46;
  wire bank13_n_47;
  wire bank13_n_48;
  wire bank13_n_49;
  wire bank13_n_50;
  wire bank13_n_51;
  wire bank13_n_52;
  wire bank13_n_89;
  wire bank13_n_90;
  wire bank13_n_91;
  wire bank13_n_92;
  wire bank13_n_93;
  wire bank13_n_94;
  wire bank13_n_95;
  wire bank13_n_96;
  wire bank13_n_97;
  wire bank13_n_98;
  wire bank13_n_99;
  wire [0:0]bank_sel;
  wire [0:0]bbus_o;
  wire \bbus_o[0]_INST_0_i_7 ;
  wire \bbus_o[0]_INST_0_i_7_0 ;
  wire \bbus_o[0]_INST_0_i_7_1 ;
  wire \bbus_o[0]_INST_0_i_7_2 ;
  wire \bbus_o[0]_INST_0_i_7_3 ;
  wire \bbus_o[0]_INST_0_i_7_4 ;
  wire \bbus_o[0]_INST_0_i_7_5 ;
  wire \bbus_o[0]_INST_0_i_7_6 ;
  wire \bbus_o[1]_INST_0_i_7 ;
  wire \bbus_o[1]_INST_0_i_7_0 ;
  wire \bbus_o[1]_INST_0_i_7_1 ;
  wire \bbus_o[1]_INST_0_i_7_2 ;
  wire \bbus_o[1]_INST_0_i_7_3 ;
  wire \bbus_o[1]_INST_0_i_7_4 ;
  wire \bbus_o[1]_INST_0_i_7_5 ;
  wire \bbus_o[1]_INST_0_i_7_6 ;
  wire \bbus_o[2]_INST_0_i_7 ;
  wire \bbus_o[2]_INST_0_i_7_0 ;
  wire \bbus_o[2]_INST_0_i_7_1 ;
  wire \bbus_o[2]_INST_0_i_7_2 ;
  wire \bbus_o[2]_INST_0_i_7_3 ;
  wire \bbus_o[2]_INST_0_i_7_4 ;
  wire \bbus_o[2]_INST_0_i_7_5 ;
  wire \bbus_o[2]_INST_0_i_7_6 ;
  wire \bbus_o[3]_INST_0_i_7 ;
  wire \bbus_o[3]_INST_0_i_7_0 ;
  wire \bbus_o[3]_INST_0_i_7_1 ;
  wire \bbus_o[3]_INST_0_i_7_2 ;
  wire \bbus_o[3]_INST_0_i_7_3 ;
  wire \bbus_o[3]_INST_0_i_7_4 ;
  wire \bbus_o[3]_INST_0_i_7_5 ;
  wire \bbus_o[3]_INST_0_i_7_6 ;
  wire \bbus_o[4]_INST_0_i_7 ;
  wire \bbus_o[4]_INST_0_i_7_0 ;
  wire \bbus_o[4]_INST_0_i_7_1 ;
  wire \bbus_o[4]_INST_0_i_7_2 ;
  wire \bbus_o[4]_INST_0_i_7_3 ;
  wire \bbus_o[4]_INST_0_i_7_4 ;
  wire \bbus_o[4]_INST_0_i_7_5 ;
  wire \bbus_o[4]_INST_0_i_7_6 ;
  wire \bbus_o[5] ;
  wire \bbus_o[5]_0 ;
  wire \bbus_o[5]_1 ;
  wire \bbus_o[6] ;
  wire \bbus_o[6]_0 ;
  wire \bbus_o[7] ;
  wire \bbus_o[7]_0 ;
  wire [1:0]bdatw;
  wire \bdatw[10] ;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_1 ;
  wire \bdatw[10]_2 ;
  wire \bdatw[10]_INST_0_i_43 ;
  wire \bdatw[10]_INST_0_i_43_0 ;
  wire \bdatw[11] ;
  wire \bdatw[11]_0 ;
  wire \bdatw[11]_1 ;
  wire \bdatw[11]_2 ;
  wire \bdatw[11]_INST_0_i_44 ;
  wire \bdatw[11]_INST_0_i_44_0 ;
  wire \bdatw[12] ;
  wire \bdatw[12]_0 ;
  wire \bdatw[12]_1 ;
  wire \bdatw[12]_2 ;
  wire \bdatw[12]_INST_0_i_42 ;
  wire \bdatw[12]_INST_0_i_42_0 ;
  wire \bdatw[13] ;
  wire \bdatw[13]_0 ;
  wire \bdatw[13]_1 ;
  wire \bdatw[13]_2 ;
  wire \bdatw[13]_3 ;
  wire \bdatw[13]_4 ;
  wire \bdatw[13]_5 ;
  wire \bdatw[14] ;
  wire \bdatw[14]_0 ;
  wire \bdatw[14]_1 ;
  wire \bdatw[14]_2 ;
  wire \bdatw[15] ;
  wire \bdatw[15]_0 ;
  wire \bdatw[8] ;
  wire \bdatw[8]_0 ;
  wire \bdatw[8]_1 ;
  wire \bdatw[8]_2 ;
  wire \bdatw[8]_INST_0_i_43 ;
  wire \bdatw[8]_INST_0_i_43_0 ;
  wire \bdatw[9] ;
  wire \bdatw[9]_0 ;
  wire \bdatw[9]_1 ;
  wire \bdatw[9]_2 ;
  wire \bdatw[9]_INST_0_i_42 ;
  wire \bdatw[9]_INST_0_i_42_0 ;
  wire clk;
  wire ctl_fetch1_fl_i_15;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [15:1]data3;
  wire [2:0]fadr;
  wire \fadr[15] ;
  wire \fadr[15]_0 ;
  wire fch_irq_req;
  wire [13:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_12_sn_1;
  wire [13:0]fdatx;
  wire \fdatx[15] ;
  wire [0:0]\grn_reg[0] ;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15] ;
  wire [15:0]\grn_reg[15]_0 ;
  wire [0:0]\grn_reg[15]_1 ;
  wire [0:0]\grn_reg[15]_10 ;
  wire [15:0]\grn_reg[15]_11 ;
  wire [0:0]\grn_reg[15]_12 ;
  wire [15:0]\grn_reg[15]_13 ;
  wire [0:0]\grn_reg[15]_14 ;
  wire [15:0]\grn_reg[15]_15 ;
  wire [0:0]\grn_reg[15]_16 ;
  wire [15:0]\grn_reg[15]_17 ;
  wire [0:0]\grn_reg[15]_18 ;
  wire [15:0]\grn_reg[15]_19 ;
  wire [0:0]\grn_reg[15]_2 ;
  wire [0:0]\grn_reg[15]_20 ;
  wire [15:0]\grn_reg[15]_21 ;
  wire [0:0]\grn_reg[15]_22 ;
  wire [15:0]\grn_reg[15]_23 ;
  wire [0:0]\grn_reg[15]_24 ;
  wire [15:0]\grn_reg[15]_25 ;
  wire [0:0]\grn_reg[15]_26 ;
  wire [15:0]\grn_reg[15]_27 ;
  wire [0:0]\grn_reg[15]_28 ;
  wire [15:0]\grn_reg[15]_29 ;
  wire [15:0]\grn_reg[15]_3 ;
  wire [0:0]\grn_reg[15]_30 ;
  wire [15:0]\grn_reg[15]_31 ;
  wire [0:0]\grn_reg[15]_32 ;
  wire [15:0]\grn_reg[15]_33 ;
  wire [0:0]\grn_reg[15]_34 ;
  wire [15:0]\grn_reg[15]_35 ;
  wire [0:0]\grn_reg[15]_36 ;
  wire [15:0]\grn_reg[15]_37 ;
  wire [0:0]\grn_reg[15]_38 ;
  wire [15:0]\grn_reg[15]_39 ;
  wire [0:0]\grn_reg[15]_4 ;
  wire [0:0]\grn_reg[15]_40 ;
  wire [15:0]\grn_reg[15]_41 ;
  wire [0:0]\grn_reg[15]_42 ;
  wire [15:0]\grn_reg[15]_43 ;
  wire [0:0]\grn_reg[15]_44 ;
  wire [15:0]\grn_reg[15]_45 ;
  wire [0:0]\grn_reg[15]_46 ;
  wire [15:0]\grn_reg[15]_47 ;
  wire [0:0]\grn_reg[15]_48 ;
  wire [15:0]\grn_reg[15]_49 ;
  wire [15:0]\grn_reg[15]_5 ;
  wire [0:0]\grn_reg[15]_50 ;
  wire [15:0]\grn_reg[15]_51 ;
  wire [0:0]\grn_reg[15]_52 ;
  wire [15:0]\grn_reg[15]_53 ;
  wire [0:0]\grn_reg[15]_54 ;
  wire [15:0]\grn_reg[15]_55 ;
  wire [0:0]\grn_reg[15]_56 ;
  wire [15:0]\grn_reg[15]_57 ;
  wire [0:0]\grn_reg[15]_58 ;
  wire [15:0]\grn_reg[15]_59 ;
  wire [0:0]\grn_reg[15]_6 ;
  wire [0:0]\grn_reg[15]_60 ;
  wire [15:0]\grn_reg[15]_61 ;
  wire [0:0]\grn_reg[15]_62 ;
  wire [15:0]\grn_reg[15]_63 ;
  wire [0:0]\grn_reg[15]_64 ;
  wire [15:0]\grn_reg[15]_65 ;
  wire [15:0]\grn_reg[15]_7 ;
  wire [0:0]\grn_reg[15]_8 ;
  wire [15:0]\grn_reg[15]_9 ;
  wire [4:0]\grn_reg[4] ;
  wire [4:0]\grn_reg[4]_0 ;
  wire [4:0]\grn_reg[4]_1 ;
  wire [4:0]\grn_reg[4]_2 ;
  wire [4:0]\grn_reg[4]_3 ;
  wire [4:0]\grn_reg[4]_4 ;
  wire [4:0]\grn_reg[4]_5 ;
  wire [4:0]\grn_reg[4]_6 ;
  wire [4:0]\grn_reg[4]_7 ;
  wire [4:0]\grn_reg[4]_8 ;
  wire [4:0]\grn_reg[4]_9 ;
  wire \i_/badr[15]_INST_0_i_19 ;
  wire \i_/badr[15]_INST_0_i_19_0 ;
  wire \i_/badr[15]_INST_0_i_19_1 ;
  wire \i_/badr[15]_INST_0_i_43 ;
  wire \i_/badr[15]_INST_0_i_43_0 ;
  wire \i_/bbus_o[4]_INST_0_i_20 ;
  wire \i_/bbus_o[4]_INST_0_i_20_0 ;
  wire \i_/bdatw[15]_INST_0_i_112 ;
  wire \i_/bdatw[15]_INST_0_i_112_0 ;
  wire \i_/bdatw[15]_INST_0_i_112_1 ;
  wire \i_/bdatw[15]_INST_0_i_113 ;
  wire \i_/bdatw[15]_INST_0_i_24 ;
  wire \i_/bdatw[15]_INST_0_i_24_0 ;
  wire \i_/bdatw[15]_INST_0_i_44 ;
  wire \i_/bdatw[15]_INST_0_i_77 ;
  wire \i_/bdatw[15]_INST_0_i_9 ;
  wire \i_/bdatw[15]_INST_0_i_9_0 ;
  wire \i_/bdatw[15]_INST_0_i_9_1 ;
  wire \i_/bdatw[15]_INST_0_i_9_2 ;
  wire \i_/bdatw[15]_INST_0_i_9_3 ;
  wire \ir0_id_fl[20]_i_4 ;
  wire irq;
  wire irq_0;
  wire [1:0]irq_lev;
  wire [15:0]\iv_reg[15] ;
  wire \iv_reg[15]_0 ;
  wire [15:0]\iv_reg[15]_1 ;
  wire \nir_id_reg[20] ;
  wire [14:0]out;
  wire [15:1]p_0_in;
  wire [15:0]p_0_in0_in;
  wire [15:0]p_0_in_1;
  wire [15:1]p_0_in_2;
  wire [15:1]p_1_in;
  wire [15:0]p_1_in1_in;
  wire p_2_in;
  wire [2:0]\pc0_reg[15] ;
  wire \pc0_reg[15]_0 ;
  wire \pc0_reg[15]_1 ;
  wire \pc_reg[13] ;
  wire \pc_reg[13]_0 ;
  wire \pc_reg[14] ;
  wire [15:0]\pc_reg[15] ;
  wire \pc_reg[15]_0 ;
  wire [2:0]\pc_reg[15]_1 ;
  wire [15:0]\pc_reg[15]_2 ;
  wire [0:0]\pc_reg[1] ;
  wire \rgf_c0bus_wb[0]_i_14 ;
  wire \rgf_c0bus_wb[10]_i_4 ;
  wire \rgf_c0bus_wb[10]_i_8 ;
  wire \rgf_c0bus_wb[11]_i_11 ;
  wire \rgf_c0bus_wb[11]_i_11_0 ;
  wire \rgf_c0bus_wb[11]_i_11_1 ;
  wire \rgf_c0bus_wb[11]_i_11_2 ;
  wire \rgf_c0bus_wb[11]_i_22 ;
  wire \rgf_c0bus_wb[11]_i_22_0 ;
  wire \rgf_c0bus_wb[11]_i_3 ;
  wire \rgf_c0bus_wb[11]_i_3_0 ;
  wire \rgf_c0bus_wb[11]_i_3_1 ;
  wire \rgf_c0bus_wb[11]_i_3_2 ;
  wire \rgf_c0bus_wb[11]_i_3_3 ;
  wire \rgf_c0bus_wb[11]_i_8 ;
  wire \rgf_c0bus_wb[11]_i_9 ;
  wire \rgf_c0bus_wb[11]_i_9_0 ;
  wire \rgf_c0bus_wb[11]_i_9_1 ;
  wire \rgf_c0bus_wb[11]_i_9_2 ;
  wire \rgf_c0bus_wb[11]_i_9_3 ;
  wire \rgf_c0bus_wb[11]_i_9_4 ;
  wire \rgf_c0bus_wb[12]_i_2 ;
  wire \rgf_c0bus_wb[12]_i_24 ;
  wire \rgf_c0bus_wb[12]_i_25 ;
  wire \rgf_c0bus_wb[13]_i_27 ;
  wire \rgf_c0bus_wb[13]_i_28 ;
  wire \rgf_c0bus_wb[13]_i_29 ;
  wire \rgf_c0bus_wb[13]_i_30 ;
  wire \rgf_c0bus_wb[13]_i_4 ;
  wire \rgf_c0bus_wb[14]_i_2 ;
  wire \rgf_c0bus_wb[15]_i_14 ;
  wire \rgf_c0bus_wb[15]_i_18 ;
  wire \rgf_c0bus_wb[15]_i_25 ;
  wire \rgf_c0bus_wb[15]_i_26 ;
  wire \rgf_c0bus_wb[15]_i_6 ;
  wire \rgf_c0bus_wb[15]_i_6_0 ;
  wire \rgf_c0bus_wb[15]_i_6_1 ;
  wire \rgf_c0bus_wb[3]_i_7 ;
  wire \rgf_c0bus_wb[3]_i_7_0 ;
  wire [15:0]\rgf_c0bus_wb[4]_i_21 ;
  wire \rgf_c0bus_wb[4]_i_26 ;
  wire \rgf_c0bus_wb[4]_i_29 ;
  wire \rgf_c0bus_wb[4]_i_31 ;
  wire \rgf_c0bus_wb[4]_i_32 ;
  wire \rgf_c0bus_wb[4]_i_33 ;
  wire \rgf_c0bus_wb[6]_i_11 ;
  wire \rgf_c0bus_wb[7]_i_7 ;
  wire \rgf_c0bus_wb[7]_i_7_0 ;
  wire \rgf_c0bus_wb[8]_i_6 ;
  wire \rgf_c0bus_wb_reg[10] ;
  wire \rgf_c0bus_wb_reg[10]_0 ;
  wire \rgf_c0bus_wb_reg[10]_1 ;
  wire [15:0]\rgf_c0bus_wb_reg[15] ;
  wire [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire \rgf_c0bus_wb_reg[7]_i_11 ;
  wire \rgf_c1bus_wb[11]_i_10 ;
  wire \rgf_c1bus_wb[11]_i_10_0 ;
  wire \rgf_c1bus_wb[11]_i_10_1 ;
  wire \rgf_c1bus_wb[11]_i_10_2 ;
  wire \rgf_c1bus_wb[11]_i_10_3 ;
  wire \rgf_c1bus_wb[11]_i_10_4 ;
  wire \rgf_c1bus_wb[11]_i_10_5 ;
  wire \rgf_c1bus_wb[11]_i_13 ;
  wire \rgf_c1bus_wb[12]_i_2 ;
  wire \rgf_c1bus_wb[12]_i_20 ;
  wire \rgf_c1bus_wb[13]_i_16 ;
  wire \rgf_c1bus_wb[13]_i_9 ;
  wire \rgf_c1bus_wb[14]_i_11 ;
  wire \rgf_c1bus_wb[14]_i_11_0 ;
  wire \rgf_c1bus_wb[14]_i_28 ;
  wire \rgf_c1bus_wb[14]_i_28_0 ;
  wire \rgf_c1bus_wb[14]_i_28_1 ;
  wire \rgf_c1bus_wb[14]_i_28_2 ;
  wire \rgf_c1bus_wb[14]_i_28_3 ;
  wire \rgf_c1bus_wb[14]_i_28_4 ;
  wire \rgf_c1bus_wb[14]_i_28_5 ;
  wire \rgf_c1bus_wb[14]_i_28_6 ;
  wire \rgf_c1bus_wb[14]_i_28_7 ;
  wire \rgf_c1bus_wb[14]_i_30 ;
  wire \rgf_c1bus_wb[14]_i_32 ;
  wire \rgf_c1bus_wb[14]_i_32_0 ;
  wire \rgf_c1bus_wb[15]_i_14 ;
  wire \rgf_c1bus_wb[15]_i_14_0 ;
  wire \rgf_c1bus_wb[15]_i_14_1 ;
  wire \rgf_c1bus_wb[15]_i_14_2 ;
  wire \rgf_c1bus_wb[15]_i_14_3 ;
  wire \rgf_c1bus_wb[15]_i_19 ;
  wire \rgf_c1bus_wb[15]_i_19_0 ;
  wire \rgf_c1bus_wb[15]_i_27 ;
  wire \rgf_c1bus_wb[1]_i_14 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_22 ;
  wire \rgf_c1bus_wb[4]_i_28 ;
  wire \rgf_c1bus_wb[4]_i_32 ;
  wire \rgf_c1bus_wb[4]_i_32_0 ;
  wire \rgf_c1bus_wb[4]_i_33 ;
  wire \rgf_c1bus_wb[4]_i_34 ;
  wire \rgf_c1bus_wb[4]_i_34_0 ;
  wire \rgf_c1bus_wb[4]_i_36 ;
  wire \rgf_c1bus_wb[4]_i_36_0 ;
  wire \rgf_c1bus_wb[4]_i_37 ;
  wire \rgf_c1bus_wb[4]_i_38 ;
  wire \rgf_c1bus_wb[4]_i_38_0 ;
  wire \rgf_c1bus_wb[4]_i_40 ;
  wire \rgf_c1bus_wb[4]_i_41 ;
  wire \rgf_c1bus_wb[4]_i_42 ;
  wire \rgf_c1bus_wb[4]_i_42_0 ;
  wire \rgf_c1bus_wb[4]_i_44 ;
  wire \rgf_c1bus_wb[4]_i_45 ;
  wire \rgf_c1bus_wb[4]_i_47 ;
  wire \rgf_c1bus_wb[4]_i_48 ;
  wire \rgf_c1bus_wb[4]_i_48_0 ;
  wire \rgf_c1bus_wb[4]_i_50 ;
  wire \rgf_c1bus_wb[4]_i_50_0 ;
  wire \rgf_c1bus_wb[4]_i_51 ;
  wire \rgf_c1bus_wb[4]_i_52 ;
  wire \rgf_c1bus_wb[4]_i_52_0 ;
  wire \rgf_c1bus_wb[4]_i_53 ;
  wire \rgf_c1bus_wb[4]_i_54 ;
  wire \rgf_c1bus_wb[4]_i_54_0 ;
  wire \rgf_c1bus_wb[4]_i_56 ;
  wire \rgf_c1bus_wb[4]_i_56_0 ;
  wire \rgf_c1bus_wb[4]_i_57 ;
  wire \rgf_c1bus_wb[4]_i_58 ;
  wire \rgf_c1bus_wb[4]_i_58_0 ;
  wire \rgf_c1bus_wb[4]_i_60 ;
  wire \rgf_c1bus_wb[4]_i_60_0 ;
  wire \rgf_c1bus_wb[4]_i_61 ;
  wire \rgf_c1bus_wb[4]_i_62 ;
  wire \rgf_c1bus_wb[4]_i_62_0 ;
  wire \rgf_c1bus_wb[4]_i_64 ;
  wire \rgf_c1bus_wb[4]_i_64_0 ;
  wire \rgf_c1bus_wb[4]_i_65 ;
  wire \rgf_c1bus_wb[4]_i_67 ;
  wire \rgf_c1bus_wb[4]_i_9 ;
  wire \rgf_c1bus_wb[4]_i_9_0 ;
  wire \rgf_c1bus_wb[5]_i_10 ;
  wire \rgf_c1bus_wb[7]_i_4 ;
  wire \rgf_c1bus_wb[7]_i_4_0 ;
  wire \rgf_c1bus_wb[9]_i_17 ;
  wire \rgf_c1bus_wb_reg[0] ;
  wire \rgf_c1bus_wb_reg[10] ;
  wire [15:0]\rgf_c1bus_wb_reg[15] ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire \rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[5]_0 ;
  wire \rgf_c1bus_wb_reg[5]_1 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2] ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  wire rgf_selc0_stat;
  wire [1:0]\rgf_selc0_wb_reg[1] ;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2] ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg;
  wire [3:0]\rgf_selc1_wb[1]_i_16 ;
  wire [0:0]\rgf_selc1_wb_reg[0] ;
  wire [1:0]\rgf_selc1_wb_reg[1] ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire rst_n;
  wire [0:0]\sp_reg[0] ;
  wire \sp_reg[0]_0 ;
  wire \sp_reg[0]_1 ;
  wire \sp_reg[0]_2 ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[11]_0 ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[13]_0 ;
  wire \sp_reg[14] ;
  wire \sp_reg[14]_0 ;
  wire \sp_reg[14]_1 ;
  wire \sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire [15:0]\sp_reg[15]_1 ;
  wire [0:0]\sp_reg[1] ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[1]_1 ;
  wire \sp_reg[1]_2 ;
  wire \sp_reg[1]_3 ;
  wire \sp_reg[2] ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[2]_1 ;
  wire \sp_reg[2]_2 ;
  wire \sp_reg[3] ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[3]_1 ;
  wire \sp_reg[4] ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[4]_1 ;
  wire \sp_reg[4]_2 ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[4]_i_129 ;
  wire \sr[4]_i_133 ;
  wire \sr[4]_i_15 ;
  wire \sr[4]_i_156 ;
  wire \sr[4]_i_15_0 ;
  wire \sr[4]_i_15_1 ;
  wire \sr[4]_i_195 ;
  wire \sr[4]_i_200 ;
  wire \sr[4]_i_219 ;
  wire \sr[4]_i_220 ;
  wire \sr[4]_i_232 ;
  wire \sr[4]_i_235 ;
  wire \sr[4]_i_237 ;
  wire \sr[4]_i_239 ;
  wire \sr[4]_i_240 ;
  wire \sr[4]_i_243 ;
  wire \sr[4]_i_245 ;
  wire \sr[4]_i_27 ;
  wire \sr[4]_i_30 ;
  wire \sr[4]_i_38 ;
  wire \sr[4]_i_44 ;
  wire \sr[4]_i_55 ;
  wire \sr[4]_i_66 ;
  wire \sr[4]_i_67 ;
  wire \sr[4]_i_84 ;
  wire \sr[6]_i_11 ;
  wire \sr[6]_i_11_0 ;
  wire \sr[6]_i_11_1 ;
  wire \sr[6]_i_15 ;
  wire \sr_reg[0] ;
  wire \sr_reg[0]_0 ;
  wire [0:0]\sr_reg[0]_1 ;
  wire \sr_reg[0]_2 ;
  wire \sr_reg[10] ;
  wire \sr_reg[14] ;
  wire [15:0]\sr_reg[15] ;
  wire \sr_reg[15]_0 ;
  wire \sr_reg[15]_1 ;
  wire [15:0]\sr_reg[15]_2 ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[5]_3 ;
  wire \sr_reg[5]_4 ;
  wire \sr_reg[5]_5 ;
  wire \sr_reg[5]_6 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_11 ;
  wire \sr_reg[6]_12 ;
  wire \sr_reg[6]_13 ;
  wire \sr_reg[6]_14 ;
  wire \sr_reg[6]_15 ;
  wire \sr_reg[6]_16 ;
  wire \sr_reg[6]_17 ;
  wire \sr_reg[6]_18 ;
  wire \sr_reg[6]_19 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_20 ;
  wire \sr_reg[6]_21 ;
  wire \sr_reg[6]_22 ;
  wire \sr_reg[6]_23 ;
  wire \sr_reg[6]_24 ;
  wire \sr_reg[6]_25 ;
  wire \sr_reg[6]_26 ;
  wire \sr_reg[6]_27 ;
  wire \sr_reg[6]_28 ;
  wire \sr_reg[6]_29 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_30 ;
  wire \sr_reg[6]_31 ;
  wire \sr_reg[6]_32 ;
  wire \sr_reg[6]_33 ;
  wire \sr_reg[6]_34 ;
  wire \sr_reg[6]_35 ;
  wire \sr_reg[6]_36 ;
  wire \sr_reg[6]_37 ;
  wire \sr_reg[6]_38 ;
  wire \sr_reg[6]_39 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_40 ;
  wire \sr_reg[6]_41 ;
  wire \sr_reg[6]_42 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_7 ;
  wire \sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;
  wire \sr_reg[7] ;
  wire sreg_n_100;
  wire sreg_n_101;
  wire sreg_n_102;
  wire sreg_n_103;
  wire sreg_n_104;
  wire sreg_n_105;
  wire sreg_n_106;
  wire sreg_n_107;
  wire sreg_n_108;
  wire sreg_n_109;
  wire sreg_n_110;
  wire sreg_n_111;
  wire sreg_n_112;
  wire sreg_n_113;
  wire sreg_n_114;
  wire sreg_n_115;
  wire sreg_n_116;
  wire sreg_n_117;
  wire sreg_n_118;
  wire sreg_n_119;
  wire sreg_n_120;
  wire sreg_n_121;
  wire sreg_n_122;
  wire sreg_n_123;
  wire sreg_n_124;
  wire sreg_n_125;
  wire sreg_n_126;
  wire sreg_n_127;
  wire sreg_n_128;
  wire sreg_n_129;
  wire sreg_n_130;
  wire sreg_n_131;
  wire sreg_n_132;
  wire sreg_n_133;
  wire sreg_n_134;
  wire sreg_n_135;
  wire sreg_n_136;
  wire sreg_n_137;
  wire sreg_n_138;
  wire sreg_n_139;
  wire sreg_n_140;
  wire sreg_n_141;
  wire sreg_n_142;
  wire sreg_n_143;
  wire sreg_n_144;
  wire sreg_n_145;
  wire sreg_n_146;
  wire sreg_n_147;
  wire sreg_n_148;
  wire sreg_n_149;
  wire sreg_n_150;
  wire sreg_n_151;
  wire sreg_n_152;
  wire sreg_n_153;
  wire sreg_n_154;
  wire sreg_n_155;
  wire sreg_n_156;
  wire sreg_n_157;
  wire sreg_n_158;
  wire sreg_n_159;
  wire sreg_n_18;
  wire sreg_n_34;
  wire sreg_n_35;
  wire sreg_n_36;
  wire sreg_n_37;
  wire sreg_n_38;
  wire sreg_n_39;
  wire sreg_n_40;
  wire sreg_n_41;
  wire sreg_n_42;
  wire sreg_n_43;
  wire sreg_n_44;
  wire sreg_n_45;
  wire sreg_n_46;
  wire sreg_n_47;
  wire sreg_n_48;
  wire sreg_n_49;
  wire sreg_n_50;
  wire sreg_n_51;
  wire sreg_n_52;
  wire sreg_n_53;
  wire sreg_n_54;
  wire sreg_n_55;
  wire sreg_n_56;
  wire sreg_n_57;
  wire sreg_n_58;
  wire sreg_n_59;
  wire sreg_n_60;
  wire sreg_n_61;
  wire sreg_n_62;
  wire sreg_n_63;
  wire sreg_n_64;
  wire sreg_n_65;
  wire sreg_n_66;
  wire sreg_n_67;
  wire sreg_n_68;
  wire sreg_n_69;
  wire sreg_n_70;
  wire sreg_n_71;
  wire sreg_n_72;
  wire sreg_n_73;
  wire sreg_n_74;
  wire sreg_n_75;
  wire sreg_n_76;
  wire sreg_n_77;
  wire sreg_n_78;
  wire sreg_n_79;
  wire sreg_n_80;
  wire sreg_n_81;
  wire sreg_n_82;
  wire sreg_n_83;
  wire sreg_n_84;
  wire sreg_n_85;
  wire sreg_n_86;
  wire sreg_n_87;
  wire sreg_n_88;
  wire sreg_n_89;
  wire sreg_n_90;
  wire sreg_n_95;
  wire sreg_n_96;
  wire sreg_n_97;
  wire sreg_n_98;
  wire sreg_n_99;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[2] ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire [1:0]tout__1_carry__0_i_1__0;
  wire tout__1_carry__0_i_7__0;
  wire tout__1_carry__0_i_7__0_0;
  wire [3:0]tout__1_carry__1_i_1__0;
  wire tout__1_carry__2;
  wire tout__1_carry__2_0;
  wire tout__1_carry__2_1;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[10] ;
  wire \tr_reg[10]_0 ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[11]_1 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[12]_1 ;
  wire \tr_reg[12]_2 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[13]_1 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire \tr_reg[14]_1 ;
  wire \tr_reg[14]_2 ;
  wire [15:0]\tr_reg[15] ;
  wire \tr_reg[15]_0 ;
  wire \tr_reg[15]_1 ;
  wire [15:0]\tr_reg[15]_2 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[1]_1 ;
  wire \tr_reg[1]_2 ;
  wire \tr_reg[2] ;
  wire \tr_reg[2]_0 ;
  wire \tr_reg[3] ;
  wire \tr_reg[3]_0 ;
  wire \tr_reg[3]_1 ;
  wire \tr_reg[4] ;
  wire \tr_reg[4]_0 ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[8] ;
  wire \tr_reg[8]_0 ;
  wire \tr_reg[9] ;
  wire \tr_reg[9]_0 ;

  mcss_rgf_bus a0bus_out
       (.O(\sp_reg[1] ),
        .a0bus_sel_cr(a0bus_sel_cr),
        .\abus_o[0] (\abus_o[0] ),
        .\abus_o[0]_0 (\grn_reg[0] ),
        .\abus_o[0]_1 (\grn_reg[0]_0 ),
        .\abus_o[10] (\abus_o[10] ),
        .\abus_o[11] (\abus_o[11] ),
        .\abus_o[12] (\abus_o[12] ),
        .\abus_o[13] (\abus_o[13] ),
        .\abus_o[14] (\abus_o[14] ),
        .\abus_o[15] (\abus_o[15] ),
        .\abus_o[1] (\abus_o[1] ),
        .\abus_o[2] (\abus_o[2] ),
        .\abus_o[3] (\abus_o[3] ),
        .\abus_o[4] (\abus_o[4] ),
        .\abus_o[5] (\abus_o[5] ),
        .\abus_o[6] (\abus_o[6] ),
        .\abus_o[7] (\abus_o[7] ),
        .\abus_o[8] (\abus_o[8] ),
        .\abus_o[9] (\abus_o[9] ),
        .data3(data3),
        .\grn_reg[0] (a0bus_out_n_63),
        .\grn_reg[10] (a0bus_out_n_23),
        .\grn_reg[11] (a0bus_out_n_19),
        .\grn_reg[12] (a0bus_out_n_15),
        .\grn_reg[13] (a0bus_out_n_11),
        .\grn_reg[14] (a0bus_out_n_7),
        .\grn_reg[15] (a0bus_out_n_3),
        .\grn_reg[1] (a0bus_out_n_59),
        .\grn_reg[2] (a0bus_out_n_55),
        .\grn_reg[3] (a0bus_out_n_51),
        .\grn_reg[4] (a0bus_out_n_47),
        .\grn_reg[5] (a0bus_out_n_43),
        .\grn_reg[6] (a0bus_out_n_39),
        .\grn_reg[7] (a0bus_out_n_35),
        .\grn_reg[8] (a0bus_out_n_31),
        .\grn_reg[9] (a0bus_out_n_27),
        .out(\sr_reg[15] ),
        .p_0_in(p_0_in),
        .p_0_in_0(p_0_in_1),
        .p_1_in(p_1_in),
        .\rgf_c0bus_wb[12]_i_22 (bank02_n_452),
        .\rgf_c0bus_wb[12]_i_22_0 (bank02_n_435),
        .\rgf_c0bus_wb[12]_i_22_1 (bank02_n_341),
        .\rgf_c0bus_wb[12]_i_22_10 (bank13_n_340),
        .\rgf_c0bus_wb[12]_i_22_2 (bank02_n_340),
        .\rgf_c0bus_wb[12]_i_22_3 (bank02_n_453),
        .\rgf_c0bus_wb[12]_i_22_4 (bank02_n_436),
        .\rgf_c0bus_wb[12]_i_22_5 (bank02_n_343),
        .\rgf_c0bus_wb[12]_i_22_6 (bank02_n_342),
        .\rgf_c0bus_wb[12]_i_22_7 (bank13_n_173),
        .\rgf_c0bus_wb[12]_i_22_8 (bank13_n_189),
        .\rgf_c0bus_wb[12]_i_22_9 (bank13_n_324),
        .\rgf_c0bus_wb[12]_i_23 (bank02_n_450),
        .\rgf_c0bus_wb[12]_i_23_0 (bank02_n_433),
        .\rgf_c0bus_wb[12]_i_23_1 (bank02_n_337),
        .\rgf_c0bus_wb[12]_i_23_10 (bank13_n_338),
        .\rgf_c0bus_wb[12]_i_23_2 (bank02_n_336),
        .\rgf_c0bus_wb[12]_i_23_3 (bank02_n_451),
        .\rgf_c0bus_wb[12]_i_23_4 (bank02_n_434),
        .\rgf_c0bus_wb[12]_i_23_5 (bank02_n_339),
        .\rgf_c0bus_wb[12]_i_23_6 (bank02_n_338),
        .\rgf_c0bus_wb[12]_i_23_7 (bank13_n_171),
        .\rgf_c0bus_wb[12]_i_23_8 (bank13_n_187),
        .\rgf_c0bus_wb[12]_i_23_9 (bank13_n_322),
        .\rgf_c0bus_wb[12]_i_25 (bank02_n_454),
        .\rgf_c0bus_wb[12]_i_25_0 (bank02_n_437),
        .\rgf_c0bus_wb[12]_i_25_1 (bank02_n_345),
        .\rgf_c0bus_wb[12]_i_25_10 (bank13_n_342),
        .\rgf_c0bus_wb[12]_i_25_2 (bank02_n_344),
        .\rgf_c0bus_wb[12]_i_25_3 (bank02_n_455),
        .\rgf_c0bus_wb[12]_i_25_4 (bank02_n_438),
        .\rgf_c0bus_wb[12]_i_25_5 (bank02_n_347),
        .\rgf_c0bus_wb[12]_i_25_6 (bank02_n_346),
        .\rgf_c0bus_wb[12]_i_25_7 (bank13_n_175),
        .\rgf_c0bus_wb[12]_i_25_8 (bank13_n_191),
        .\rgf_c0bus_wb[12]_i_25_9 (bank13_n_326),
        .\rgf_c0bus_wb[13]_i_30 (bank02_n_459),
        .\rgf_c0bus_wb[13]_i_30_0 (bank02_n_442),
        .\rgf_c0bus_wb[13]_i_30_1 (bank02_n_355),
        .\rgf_c0bus_wb[13]_i_30_10 (bank13_n_347),
        .\rgf_c0bus_wb[13]_i_30_2 (bank02_n_354),
        .\rgf_c0bus_wb[13]_i_30_3 (bank02_n_460),
        .\rgf_c0bus_wb[13]_i_30_4 (bank02_n_443),
        .\rgf_c0bus_wb[13]_i_30_5 (bank02_n_357),
        .\rgf_c0bus_wb[13]_i_30_6 (bank02_n_356),
        .\rgf_c0bus_wb[13]_i_30_7 (bank13_n_180),
        .\rgf_c0bus_wb[13]_i_30_8 (bank13_n_196),
        .\rgf_c0bus_wb[13]_i_30_9 (bank13_n_331),
        .\rgf_c0bus_wb[13]_i_31 (bank02_n_457),
        .\rgf_c0bus_wb[13]_i_31_0 (bank02_n_440),
        .\rgf_c0bus_wb[13]_i_31_1 (bank02_n_351),
        .\rgf_c0bus_wb[13]_i_31_10 (bank13_n_345),
        .\rgf_c0bus_wb[13]_i_31_2 (bank02_n_350),
        .\rgf_c0bus_wb[13]_i_31_3 (bank02_n_458),
        .\rgf_c0bus_wb[13]_i_31_4 (bank02_n_441),
        .\rgf_c0bus_wb[13]_i_31_5 (bank02_n_353),
        .\rgf_c0bus_wb[13]_i_31_6 (bank02_n_352),
        .\rgf_c0bus_wb[13]_i_31_7 (bank13_n_178),
        .\rgf_c0bus_wb[13]_i_31_8 (bank13_n_194),
        .\rgf_c0bus_wb[13]_i_31_9 (bank13_n_329),
        .\rgf_c0bus_wb[13]_i_32 (bank02_n_461),
        .\rgf_c0bus_wb[13]_i_32_0 (bank02_n_444),
        .\rgf_c0bus_wb[13]_i_32_1 (bank02_n_359),
        .\rgf_c0bus_wb[13]_i_32_10 (bank13_n_349),
        .\rgf_c0bus_wb[13]_i_32_2 (bank02_n_358),
        .\rgf_c0bus_wb[13]_i_32_3 (bank02_n_462),
        .\rgf_c0bus_wb[13]_i_32_4 (bank02_n_446),
        .\rgf_c0bus_wb[13]_i_32_5 (bank02_n_362),
        .\rgf_c0bus_wb[13]_i_32_6 (bank02_n_361),
        .\rgf_c0bus_wb[13]_i_32_7 (bank13_n_182),
        .\rgf_c0bus_wb[13]_i_32_8 (bank13_n_198),
        .\rgf_c0bus_wb[13]_i_32_9 (bank13_n_333),
        .\rgf_c0bus_wb[15]_i_30 (bank13_n_181),
        .\rgf_c0bus_wb[15]_i_30_0 (bank13_n_197),
        .\rgf_c0bus_wb[15]_i_30_1 (bank13_n_332),
        .\rgf_c0bus_wb[15]_i_30_2 (bank13_n_348),
        .\rgf_c0bus_wb[4]_i_20 (bank13_n_183),
        .\rgf_c0bus_wb[4]_i_20_0 (bank13_n_199),
        .\rgf_c0bus_wb[4]_i_20_1 (bank13_n_334),
        .\rgf_c0bus_wb[4]_i_20_2 (bank13_n_350),
        .\rgf_c0bus_wb[4]_i_21 (bank02_n_447),
        .\rgf_c0bus_wb[4]_i_21_0 (bank02_n_430),
        .\rgf_c0bus_wb[4]_i_21_1 (bank02_n_331),
        .\rgf_c0bus_wb[4]_i_21_10 (bank13_n_335),
        .\rgf_c0bus_wb[4]_i_21_11 ({p_0_in_2,\sp_reg[0] }),
        .\rgf_c0bus_wb[4]_i_21_12 (\rgf_c0bus_wb[4]_i_21 ),
        .\rgf_c0bus_wb[4]_i_21_2 (bank02_n_330),
        .\rgf_c0bus_wb[4]_i_21_3 (bank02_n_448),
        .\rgf_c0bus_wb[4]_i_21_4 (bank02_n_431),
        .\rgf_c0bus_wb[4]_i_21_5 (bank02_n_333),
        .\rgf_c0bus_wb[4]_i_21_6 (bank02_n_332),
        .\rgf_c0bus_wb[4]_i_21_7 (bank13_n_168),
        .\rgf_c0bus_wb[4]_i_21_8 (bank13_n_184),
        .\rgf_c0bus_wb[4]_i_21_9 (bank13_n_319),
        .\rgf_c0bus_wb[4]_i_23 (bank13_n_172),
        .\rgf_c0bus_wb[4]_i_23_0 (bank13_n_188),
        .\rgf_c0bus_wb[4]_i_23_1 (bank13_n_323),
        .\rgf_c0bus_wb[4]_i_23_2 (bank13_n_339),
        .\rgf_c0bus_wb[4]_i_24 (bank13_n_170),
        .\rgf_c0bus_wb[4]_i_24_0 (bank13_n_186),
        .\rgf_c0bus_wb[4]_i_24_1 (bank13_n_321),
        .\rgf_c0bus_wb[4]_i_24_2 (bank13_n_337),
        .\rgf_c0bus_wb[4]_i_25 (bank02_n_456),
        .\rgf_c0bus_wb[4]_i_25_0 (bank02_n_439),
        .\rgf_c0bus_wb[4]_i_25_1 (bank02_n_349),
        .\rgf_c0bus_wb[4]_i_25_2 (bank02_n_348),
        .\rgf_c0bus_wb[4]_i_25_3 (bank13_n_176),
        .\rgf_c0bus_wb[4]_i_25_4 (bank13_n_192),
        .\rgf_c0bus_wb[4]_i_25_5 (bank13_n_327),
        .\rgf_c0bus_wb[4]_i_25_6 (bank13_n_343),
        .\rgf_c0bus_wb[4]_i_26 (bank13_n_174),
        .\rgf_c0bus_wb[4]_i_26_0 (bank13_n_190),
        .\rgf_c0bus_wb[4]_i_26_1 (bank13_n_325),
        .\rgf_c0bus_wb[4]_i_26_2 (bank13_n_341),
        .\rgf_c0bus_wb[4]_i_29 (bank13_n_177),
        .\rgf_c0bus_wb[4]_i_29_0 (bank13_n_193),
        .\rgf_c0bus_wb[4]_i_29_1 (bank13_n_328),
        .\rgf_c0bus_wb[4]_i_29_2 (bank13_n_344),
        .\rgf_c0bus_wb[4]_i_30 (bank13_n_179),
        .\rgf_c0bus_wb[4]_i_30_0 (bank13_n_195),
        .\rgf_c0bus_wb[4]_i_30_1 (bank13_n_330),
        .\rgf_c0bus_wb[4]_i_30_2 (bank13_n_346),
        .\sp_reg[0] (\sp_reg[0]_0 ),
        .\sp_reg[10] (a0bus_out_n_22),
        .\sp_reg[11] (a0bus_out_n_18),
        .\sp_reg[12] (a0bus_out_n_14),
        .\sp_reg[13] (a0bus_out_n_10),
        .\sp_reg[14] (a0bus_out_n_6),
        .\sp_reg[15] (a0bus_out_n_2),
        .\sp_reg[1] (a0bus_out_n_58),
        .\sp_reg[2] (a0bus_out_n_54),
        .\sp_reg[3] (a0bus_out_n_50),
        .\sp_reg[4] (a0bus_out_n_46),
        .\sp_reg[5] (a0bus_out_n_42),
        .\sp_reg[6] (a0bus_out_n_38),
        .\sp_reg[7] (a0bus_out_n_34),
        .\sp_reg[8] (a0bus_out_n_30),
        .\sp_reg[9] (a0bus_out_n_26),
        .\sr[4]_i_226 (bank02_n_449),
        .\sr[4]_i_226_0 (bank02_n_432),
        .\sr[4]_i_226_1 (bank02_n_335),
        .\sr[4]_i_226_2 (bank02_n_334),
        .\sr[4]_i_226_3 (bank13_n_169),
        .\sr[4]_i_226_4 (bank13_n_185),
        .\sr[4]_i_226_5 (bank13_n_320),
        .\sr[4]_i_226_6 (bank13_n_336),
        .\sr_reg[0] (\sr_reg[0] ),
        .\sr_reg[0]_0 (a0bus_out_n_79),
        .\sr_reg[10] (a0bus_out_n_21),
        .\sr_reg[10]_0 (a0bus_out_n_69),
        .\sr_reg[11] (a0bus_out_n_17),
        .\sr_reg[11]_0 (a0bus_out_n_68),
        .\sr_reg[12] (a0bus_out_n_13),
        .\sr_reg[12]_0 (a0bus_out_n_67),
        .\sr_reg[13] (a0bus_out_n_9),
        .\sr_reg[13]_0 (a0bus_out_n_66),
        .\sr_reg[14] (a0bus_out_n_5),
        .\sr_reg[14]_0 (a0bus_out_n_65),
        .\sr_reg[15] (a0bus_out_n_1),
        .\sr_reg[15]_0 (a0bus_out_n_64),
        .\sr_reg[1] (a0bus_out_n_57),
        .\sr_reg[1]_0 (a0bus_out_n_78),
        .\sr_reg[2] (a0bus_out_n_53),
        .\sr_reg[2]_0 (a0bus_out_n_77),
        .\sr_reg[3] (a0bus_out_n_49),
        .\sr_reg[3]_0 (a0bus_out_n_76),
        .\sr_reg[4] (a0bus_out_n_45),
        .\sr_reg[4]_0 (a0bus_out_n_75),
        .\sr_reg[5] (a0bus_out_n_41),
        .\sr_reg[5]_0 (a0bus_out_n_74),
        .\sr_reg[6] (a0bus_out_n_37),
        .\sr_reg[6]_0 (a0bus_out_n_73),
        .\sr_reg[7] (a0bus_out_n_33),
        .\sr_reg[7]_0 (a0bus_out_n_72),
        .\sr_reg[8] (a0bus_out_n_29),
        .\sr_reg[8]_0 (a0bus_out_n_71),
        .\sr_reg[9] (a0bus_out_n_25),
        .\sr_reg[9]_0 (a0bus_out_n_70),
        .\tr_reg[0] (a0bus_0[0]),
        .\tr_reg[10] (a0bus_0[10]),
        .\tr_reg[11] (a0bus_0[11]),
        .\tr_reg[12] (a0bus_0[12]),
        .\tr_reg[13] (a0bus_0[13]),
        .\tr_reg[14] (a0bus_0[14]),
        .\tr_reg[15] (a0bus_0[15]),
        .\tr_reg[1] (a0bus_0[1]),
        .\tr_reg[2] (a0bus_0[2]),
        .\tr_reg[3] (a0bus_0[3]),
        .\tr_reg[4] (a0bus_0[4]),
        .\tr_reg[5] (a0bus_0[5]),
        .\tr_reg[6] (a0bus_0[6]),
        .\tr_reg[7] (a0bus_0[7]),
        .\tr_reg[8] (a0bus_0[8]),
        .\tr_reg[9] (a0bus_0[9]));
  mcss_rgf_bus_2 a1bus_out
       (.O(\sp_reg[1] ),
        .a1bus_b13(a1bus_b13),
        .a1bus_sel_cr(a1bus_sel_cr),
        .a1bus_sr(a1bus_sr),
        .data3(data3),
        .\grn_reg[0] (a1bus_out_n_48),
        .\grn_reg[10] (a1bus_out_n_18),
        .\grn_reg[11] (a1bus_out_n_15),
        .\grn_reg[12] (a1bus_out_n_12),
        .\grn_reg[13] (a1bus_out_n_9),
        .\grn_reg[14] (a1bus_out_n_6),
        .\grn_reg[15] (a1bus_out_n_3),
        .\grn_reg[1] (a1bus_out_n_44),
        .\grn_reg[2] (a1bus_out_n_41),
        .\grn_reg[3] (a1bus_out_n_38),
        .\grn_reg[4] (a1bus_out_n_35),
        .\grn_reg[5] (a1bus_out_n_32),
        .\grn_reg[6] (a1bus_out_n_29),
        .\grn_reg[7] (a1bus_out_n_26),
        .\grn_reg[9] (a1bus_out_n_21),
        .out(\tr_reg[15] ),
        .p_0_in0_in(p_0_in0_in),
        .p_1_in1_in(p_1_in1_in),
        .\rgf_c1bus_wb[4]_i_18 (bank02_n_511),
        .\rgf_c1bus_wb[4]_i_18_0 (bank02_n_495),
        .\rgf_c1bus_wb[4]_i_18_1 (sreg_n_108),
        .\rgf_c1bus_wb[4]_i_18_2 (bank02_n_407),
        .\rgf_c1bus_wb[4]_i_18_3 (bank02_n_406),
        .\rgf_c1bus_wb[4]_i_18_4 (bank13_n_244),
        .\rgf_c1bus_wb[4]_i_18_5 (bank13_n_262),
        .\rgf_c1bus_wb[4]_i_18_6 (bank13_n_412),
        .\rgf_c1bus_wb[4]_i_18_7 (bank13_n_396),
        .\rgf_c1bus_wb[4]_i_19 (bank02_n_513),
        .\rgf_c1bus_wb[4]_i_19_0 (bank02_n_497),
        .\rgf_c1bus_wb[4]_i_19_1 (sreg_n_110),
        .\rgf_c1bus_wb[4]_i_19_10 (bank13_n_414),
        .\rgf_c1bus_wb[4]_i_19_11 (bank13_n_398),
        .\rgf_c1bus_wb[4]_i_19_2 (bank02_n_411),
        .\rgf_c1bus_wb[4]_i_19_3 (bank02_n_410),
        .\rgf_c1bus_wb[4]_i_19_4 (bank13_n_245),
        .\rgf_c1bus_wb[4]_i_19_5 (bank13_n_263),
        .\rgf_c1bus_wb[4]_i_19_6 (bank13_n_413),
        .\rgf_c1bus_wb[4]_i_19_7 (bank13_n_397),
        .\rgf_c1bus_wb[4]_i_19_8 (bank13_n_246),
        .\rgf_c1bus_wb[4]_i_19_9 (bank13_n_264),
        .\rgf_c1bus_wb[4]_i_20 (bank02_n_501),
        .\rgf_c1bus_wb[4]_i_20_0 (bank02_n_485),
        .\rgf_c1bus_wb[4]_i_20_1 (sreg_n_97),
        .\rgf_c1bus_wb[4]_i_20_2 (bank02_n_387),
        .\rgf_c1bus_wb[4]_i_20_3 (bank02_n_386),
        .\rgf_c1bus_wb[4]_i_20_4 (bank13_n_248),
        .\rgf_c1bus_wb[4]_i_21 (bank13_n_247),
        .\rgf_c1bus_wb[4]_i_21_0 (bank13_n_415),
        .\rgf_c1bus_wb[4]_i_21_1 (bank13_n_399),
        .\rgf_c1bus_wb[4]_i_21_2 (sreg_n_128),
        .\rgf_c1bus_wb[4]_i_21_3 (bank13_n_266),
        .\rgf_c1bus_wb[4]_i_22 (bank13_n_232),
        .\rgf_c1bus_wb[4]_i_22_0 (bank13_n_400),
        .\rgf_c1bus_wb[4]_i_22_1 (bank13_n_383),
        .\rgf_c1bus_wb[4]_i_22_2 (sreg_n_143),
        .\rgf_c1bus_wb[4]_i_22_3 (bank13_n_250),
        .\rgf_c1bus_wb[4]_i_22_4 (\iv_reg[15] ),
        .\rgf_c1bus_wb[4]_i_22_5 ({p_0_in_2,\sp_reg[0] }),
        .\rgf_c1bus_wb[4]_i_22_6 (\rgf_c1bus_wb[4]_i_22 ),
        .\rgf_c1bus_wb[4]_i_23 (bank02_n_499),
        .\rgf_c1bus_wb[4]_i_23_0 (bank02_n_484),
        .\rgf_c1bus_wb[4]_i_23_1 (sreg_n_96),
        .\rgf_c1bus_wb[4]_i_23_2 (bank02_n_385),
        .\rgf_c1bus_wb[4]_i_23_3 (bank02_n_384),
        .\sp_reg[0] (a1bus_out_n_47),
        .\sp_reg[0]_0 (a1bus_out_n_65),
        .\sp_reg[10] (a1bus_out_n_55),
        .\sp_reg[11] (a1bus_out_n_54),
        .\sp_reg[12] (a1bus_out_n_53),
        .\sp_reg[13] (a1bus_out_n_52),
        .\sp_reg[14] (a1bus_out_n_51),
        .\sp_reg[15] (\sp_reg[15]_0 ),
        .\sp_reg[15]_0 (a1bus_out_n_49),
        .\sp_reg[1] (a1bus_out_n_64),
        .\sp_reg[2] (a1bus_out_n_63),
        .\sp_reg[3] (a1bus_out_n_62),
        .\sp_reg[4] (a1bus_out_n_61),
        .\sp_reg[5] (a1bus_out_n_60),
        .\sp_reg[6] (a1bus_out_n_59),
        .\sp_reg[7] (a1bus_out_n_58),
        .\sp_reg[8] (a1bus_out_n_57),
        .\sp_reg[9] (a1bus_out_n_56),
        .\sr[4]_i_207 (bank02_n_503),
        .\sr[4]_i_207_0 (bank02_n_487),
        .\sr[4]_i_207_1 (sreg_n_99),
        .\sr[4]_i_207_2 (bank02_n_391),
        .\sr[4]_i_207_3 (bank02_n_390),
        .\sr[4]_i_208 (bank02_n_505),
        .\sr[4]_i_208_0 (bank02_n_489),
        .\sr[4]_i_208_1 (sreg_n_101),
        .\sr[4]_i_208_2 (bank02_n_395),
        .\sr[4]_i_208_3 (bank02_n_394),
        .\sr[4]_i_210 (bank13_n_265),
        .\sr[4]_i_213 (bank02_n_514),
        .\sr[4]_i_213_0 (bank02_n_498),
        .\sr[4]_i_213_1 (sreg_n_111),
        .\sr[4]_i_213_2 (bank02_n_413),
        .\sr[4]_i_213_3 (bank02_n_412),
        .\sr[4]_i_215 (bank02_n_504),
        .\sr[4]_i_215_0 (bank02_n_488),
        .\sr[4]_i_215_1 (sreg_n_100),
        .\sr[4]_i_215_10 (bank13_n_404),
        .\sr[4]_i_215_11 (bank13_n_388),
        .\sr[4]_i_215_2 (bank02_n_393),
        .\sr[4]_i_215_3 (bank02_n_392),
        .\sr[4]_i_215_4 (bank13_n_235),
        .\sr[4]_i_215_5 (bank13_n_253),
        .\sr[4]_i_215_6 (bank13_n_403),
        .\sr[4]_i_215_7 (bank13_n_387),
        .\sr[4]_i_215_8 (bank13_n_236),
        .\sr[4]_i_215_9 (bank13_n_254),
        .\sr[4]_i_216 (bank02_n_502),
        .\sr[4]_i_216_0 (bank02_n_486),
        .\sr[4]_i_216_1 (sreg_n_98),
        .\sr[4]_i_216_10 (bank13_n_402),
        .\sr[4]_i_216_11 (bank13_n_386),
        .\sr[4]_i_216_2 (bank02_n_389),
        .\sr[4]_i_216_3 (bank02_n_388),
        .\sr[4]_i_216_4 (bank13_n_233),
        .\sr[4]_i_216_5 (bank13_n_251),
        .\sr[4]_i_216_6 (bank13_n_401),
        .\sr[4]_i_216_7 (bank13_n_385),
        .\sr[4]_i_216_8 (bank13_n_234),
        .\sr[4]_i_216_9 (bank13_n_252),
        .\sr[4]_i_217 (bank02_n_507),
        .\sr[4]_i_217_0 (bank02_n_491),
        .\sr[4]_i_217_1 (sreg_n_104),
        .\sr[4]_i_217_2 (bank02_n_399),
        .\sr[4]_i_217_3 (bank02_n_398),
        .\sr[4]_i_217_4 (bank13_n_239),
        .\sr[4]_i_217_5 (bank13_n_257),
        .\sr[4]_i_217_6 (bank13_n_407),
        .\sr[4]_i_217_7 (bank13_n_391),
        .\sr[4]_i_218 (bank02_n_506),
        .\sr[4]_i_218_0 (bank02_n_490),
        .\sr[4]_i_218_1 (sreg_n_102),
        .\sr[4]_i_218_10 (bank13_n_406),
        .\sr[4]_i_218_11 (bank13_n_390),
        .\sr[4]_i_218_2 (bank02_n_397),
        .\sr[4]_i_218_3 (bank02_n_396),
        .\sr[4]_i_218_4 (bank13_n_237),
        .\sr[4]_i_218_5 (bank13_n_255),
        .\sr[4]_i_218_6 (bank13_n_405),
        .\sr[4]_i_218_7 (bank13_n_389),
        .\sr[4]_i_218_8 (bank13_n_238),
        .\sr[4]_i_218_9 (bank13_n_256),
        .\sr[4]_i_219 (bank02_n_509),
        .\sr[4]_i_219_0 (bank02_n_493),
        .\sr[4]_i_219_1 (sreg_n_106),
        .\sr[4]_i_219_2 (bank02_n_403),
        .\sr[4]_i_219_3 (bank02_n_402),
        .\sr[4]_i_220 (bank02_n_512),
        .\sr[4]_i_220_0 (bank02_n_496),
        .\sr[4]_i_220_1 (sreg_n_109),
        .\sr[4]_i_220_2 (bank02_n_409),
        .\sr[4]_i_220_3 (bank02_n_408),
        .\sr[4]_i_224 (bank02_n_510),
        .\sr[4]_i_224_0 (bank02_n_494),
        .\sr[4]_i_224_1 (sreg_n_107),
        .\sr[4]_i_224_10 (bank13_n_411),
        .\sr[4]_i_224_11 (bank13_n_395),
        .\sr[4]_i_224_2 (bank02_n_405),
        .\sr[4]_i_224_3 (bank02_n_404),
        .\sr[4]_i_224_4 (bank13_n_242),
        .\sr[4]_i_224_5 (bank13_n_260),
        .\sr[4]_i_224_6 (bank13_n_410),
        .\sr[4]_i_224_7 (bank13_n_394),
        .\sr[4]_i_224_8 (bank13_n_243),
        .\sr[4]_i_224_9 (bank13_n_261),
        .\sr[4]_i_225 (bank02_n_508),
        .\sr[4]_i_225_0 (bank02_n_492),
        .\sr[4]_i_225_1 (sreg_n_105),
        .\sr[4]_i_225_10 (bank13_n_409),
        .\sr[4]_i_225_11 (bank13_n_393),
        .\sr[4]_i_225_2 (bank02_n_401),
        .\sr[4]_i_225_3 (bank02_n_400),
        .\sr[4]_i_225_4 (bank13_n_240),
        .\sr[4]_i_225_5 (bank13_n_258),
        .\sr[4]_i_225_6 (bank13_n_408),
        .\sr[4]_i_225_7 (bank13_n_392),
        .\sr[4]_i_225_8 (bank13_n_241),
        .\sr[4]_i_225_9 (bank13_n_259),
        .\sr_reg[0] (a1bus_out_n_66),
        .\sr_reg[15] (\sr_reg[15]_0 ),
        .\tr_reg[0] (a1bus_0[0]),
        .\tr_reg[0]_0 (a1bus_out_n_46),
        .\tr_reg[10] (a1bus_0[10]),
        .\tr_reg[10]_0 (a1bus_out_n_17),
        .\tr_reg[11] (a1bus_0[11]),
        .\tr_reg[11]_0 (a1bus_out_n_14),
        .\tr_reg[12] (a1bus_0[12]),
        .\tr_reg[12]_0 (a1bus_out_n_11),
        .\tr_reg[13] (a1bus_0[13]),
        .\tr_reg[13]_0 (a1bus_out_n_8),
        .\tr_reg[14] (a1bus_0[14]),
        .\tr_reg[14]_0 (a1bus_out_n_5),
        .\tr_reg[15] (a1bus_0[15]),
        .\tr_reg[15]_0 (\tr_reg[15]_0 ),
        .\tr_reg[1] (a1bus_0[1]),
        .\tr_reg[1]_0 (a1bus_out_n_43),
        .\tr_reg[2] (a1bus_0[2]),
        .\tr_reg[2]_0 (a1bus_out_n_40),
        .\tr_reg[3] (a1bus_0[3]),
        .\tr_reg[3]_0 (a1bus_out_n_37),
        .\tr_reg[4] (a1bus_0[4]),
        .\tr_reg[4]_0 (a1bus_out_n_34),
        .\tr_reg[5] (a1bus_0[5]),
        .\tr_reg[5]_0 (a1bus_out_n_31),
        .\tr_reg[6] (a1bus_0[6]),
        .\tr_reg[6]_0 (a1bus_out_n_28),
        .\tr_reg[7] (a1bus_0[7]),
        .\tr_reg[7]_0 (a1bus_out_n_25),
        .\tr_reg[8] (a1bus_0[8]),
        .\tr_reg[8]_0 (a1bus_out_n_23),
        .\tr_reg[9] (a1bus_0[9]),
        .\tr_reg[9]_0 (a1bus_out_n_20));
  mcss_rgf_bus_3 b0bus_out
       (.O(\sp_reg[1] ),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b0bus_sr(b0bus_sr),
        .\bbus_o[0]_INST_0_i_1 (bank13_n_215),
        .\bbus_o[0]_INST_0_i_1_0 (bank13_n_231),
        .\bbus_o[0]_INST_0_i_1_1 (bank13_n_382),
        .\bbus_o[0]_INST_0_i_1_2 (bank13_n_366),
        .\bbus_o[1]_INST_0_i_1 (bank13_n_214),
        .\bbus_o[1]_INST_0_i_1_0 (bank13_n_230),
        .\bbus_o[1]_INST_0_i_1_1 (bank13_n_381),
        .\bbus_o[1]_INST_0_i_1_2 (bank13_n_365),
        .\bbus_o[2]_INST_0_i_1 (bank13_n_213),
        .\bbus_o[2]_INST_0_i_1_0 (bank13_n_229),
        .\bbus_o[2]_INST_0_i_1_1 (bank13_n_380),
        .\bbus_o[2]_INST_0_i_1_2 (bank13_n_364),
        .\bbus_o[3]_INST_0_i_1 (bank13_n_212),
        .\bbus_o[3]_INST_0_i_1_0 (bank13_n_228),
        .\bbus_o[3]_INST_0_i_1_1 (bank13_n_379),
        .\bbus_o[3]_INST_0_i_1_2 (bank13_n_363),
        .\bbus_o[4]_INST_0_i_1 (bank13_n_211),
        .\bbus_o[4]_INST_0_i_1_0 (bank13_n_227),
        .\bbus_o[4]_INST_0_i_1_1 (bank13_n_378),
        .\bbus_o[4]_INST_0_i_1_2 (bank13_n_362),
        .\bbus_o[5]_INST_0_i_1 (bank13_n_210),
        .\bbus_o[5]_INST_0_i_1_0 (bank13_n_226),
        .\bbus_o[5]_INST_0_i_1_1 (bank13_n_377),
        .\bbus_o[5]_INST_0_i_1_2 (bank13_n_361),
        .\bbus_o[6]_INST_0_i_1 (bank13_n_209),
        .\bbus_o[6]_INST_0_i_1_0 (bank13_n_225),
        .\bbus_o[6]_INST_0_i_1_1 (bank13_n_376),
        .\bbus_o[6]_INST_0_i_1_2 (bank13_n_360),
        .\bbus_o[7]_INST_0_i_1 (bank13_n_208),
        .\bbus_o[7]_INST_0_i_1_0 (bank13_n_224),
        .\bbus_o[7]_INST_0_i_1_1 (bank13_n_375),
        .\bbus_o[7]_INST_0_i_1_2 (bank13_n_359),
        .\bdatw[10]_INST_0_i_1 (bank13_n_205),
        .\bdatw[10]_INST_0_i_1_0 (bank13_n_221),
        .\bdatw[10]_INST_0_i_1_1 (bank13_n_372),
        .\bdatw[10]_INST_0_i_1_2 (bank13_n_356),
        .\bdatw[11]_INST_0_i_1 (bank13_n_204),
        .\bdatw[11]_INST_0_i_1_0 (bank13_n_220),
        .\bdatw[11]_INST_0_i_1_1 (bank13_n_371),
        .\bdatw[11]_INST_0_i_1_2 (bank13_n_355),
        .\bdatw[12]_INST_0_i_1 (bank13_n_203),
        .\bdatw[12]_INST_0_i_1_0 (bank13_n_219),
        .\bdatw[12]_INST_0_i_1_1 (bank13_n_370),
        .\bdatw[12]_INST_0_i_1_2 (bank13_n_354),
        .\bdatw[13]_INST_0_i_1 (bank13_n_202),
        .\bdatw[13]_INST_0_i_1_0 (bank13_n_218),
        .\bdatw[13]_INST_0_i_1_1 (bank13_n_369),
        .\bdatw[13]_INST_0_i_1_2 (bank13_n_353),
        .\bdatw[14]_INST_0_i_1 (bank13_n_201),
        .\bdatw[14]_INST_0_i_1_0 (bank13_n_217),
        .\bdatw[14]_INST_0_i_1_1 (bank13_n_368),
        .\bdatw[14]_INST_0_i_1_2 (bank13_n_352),
        .\bdatw[15]_INST_0_i_1 (bank13_n_200),
        .\bdatw[15]_INST_0_i_11_0 ({p_0_in_2,\sp_reg[0] }),
        .\bdatw[15]_INST_0_i_11_1 (\rgf_c0bus_wb[4]_i_21 ),
        .\bdatw[15]_INST_0_i_1_0 (bank13_n_216),
        .\bdatw[15]_INST_0_i_1_1 (bank13_n_367),
        .\bdatw[15]_INST_0_i_1_2 (bank13_n_351),
        .\bdatw[15]_INST_0_i_1_3 (\iv_reg[15] ),
        .\bdatw[8]_INST_0_i_1 (bank13_n_207),
        .\bdatw[8]_INST_0_i_1_0 (bank13_n_223),
        .\bdatw[8]_INST_0_i_1_1 (bank13_n_374),
        .\bdatw[8]_INST_0_i_1_2 (bank13_n_358),
        .\bdatw[9]_INST_0_i_1 (bank13_n_206),
        .\bdatw[9]_INST_0_i_1_0 (bank13_n_222),
        .\bdatw[9]_INST_0_i_1_1 (bank13_n_373),
        .\bdatw[9]_INST_0_i_1_2 (bank13_n_357),
        .data3(data3),
        .out(\tr_reg[15] ),
        .\sp_reg[0] (\sp_reg[0]_1 ),
        .\sp_reg[10] (b0bus_out_n_5),
        .\sp_reg[11] (b0bus_out_n_4),
        .\sp_reg[12] (b0bus_out_n_3),
        .\sp_reg[13] (b0bus_out_n_2),
        .\sp_reg[14] (b0bus_out_n_1),
        .\sp_reg[15] (b0bus_out_n_0),
        .\sp_reg[1] (\sp_reg[1]_2 ),
        .\sp_reg[2] (\sp_reg[2]_1 ),
        .\sp_reg[3] (\sp_reg[3]_0 ),
        .\sp_reg[4] (\sp_reg[4]_1 ),
        .\sp_reg[5] (b0bus_out_n_10),
        .\sp_reg[6] (b0bus_out_n_9),
        .\sp_reg[7] (b0bus_out_n_8),
        .\sp_reg[8] (b0bus_out_n_7),
        .\sp_reg[9] (b0bus_out_n_6),
        .\tr_reg[0] (\tr_reg[0] ),
        .\tr_reg[10] (b0bus_out_n_26),
        .\tr_reg[11] (b0bus_out_n_27),
        .\tr_reg[12] (b0bus_out_n_28),
        .\tr_reg[13] (b0bus_out_n_29),
        .\tr_reg[14] (b0bus_out_n_30),
        .\tr_reg[15] (b0bus_out_n_31),
        .\tr_reg[1] (\tr_reg[1]_1 ),
        .\tr_reg[2] (\tr_reg[2] ),
        .\tr_reg[3] (\tr_reg[3]_0 ),
        .\tr_reg[4] (\tr_reg[4] ),
        .\tr_reg[5] (b0bus_out_n_21),
        .\tr_reg[6] (b0bus_out_n_22),
        .\tr_reg[7] (b0bus_out_n_23),
        .\tr_reg[8] (b0bus_out_n_24),
        .\tr_reg[9] (b0bus_out_n_25));
  mcss_rgf_bus_4 b1bus_out
       (.O(\sp_reg[1] ),
        .b1bus_sel_cr(b1bus_sel_cr),
        .b1bus_sr(b1bus_sr),
        .\bdatw[10]_INST_0_i_16 (bank13_n_429),
        .\bdatw[10]_INST_0_i_16_0 (bank13_n_444),
        .\bdatw[10]_INST_0_i_16_1 (bank13_n_300),
        .\bdatw[10]_INST_0_i_16_2 (bank13_n_295),
        .\bdatw[10]_INST_0_i_16_3 (bank13_n_280),
        .\bdatw[10]_INST_0_i_2 (bank13_n_272),
        .\bdatw[10]_INST_0_i_2_0 (bank13_n_287),
        .\bdatw[10]_INST_0_i_2_1 (bank13_n_436),
        .\bdatw[10]_INST_0_i_2_2 (bank13_n_421),
        .\bdatw[11]_INST_0_i_16 (bank13_n_428),
        .\bdatw[11]_INST_0_i_16_0 (bank13_n_443),
        .\bdatw[11]_INST_0_i_16_1 (bank13_n_299),
        .\bdatw[11]_INST_0_i_16_2 (bank13_n_294),
        .\bdatw[11]_INST_0_i_16_3 (bank13_n_279),
        .\bdatw[11]_INST_0_i_2 (bank13_n_271),
        .\bdatw[11]_INST_0_i_2_0 (bank13_n_286),
        .\bdatw[11]_INST_0_i_2_1 (bank13_n_435),
        .\bdatw[11]_INST_0_i_2_2 (bank13_n_420),
        .\bdatw[12]_INST_0_i_16 (bank13_n_427),
        .\bdatw[12]_INST_0_i_16_0 (bank13_n_442),
        .\bdatw[12]_INST_0_i_16_1 (bank13_n_298),
        .\bdatw[12]_INST_0_i_16_2 (bank13_n_293),
        .\bdatw[12]_INST_0_i_16_3 (bank13_n_278),
        .\bdatw[12]_INST_0_i_2 (bank13_n_270),
        .\bdatw[12]_INST_0_i_2_0 (bank13_n_285),
        .\bdatw[12]_INST_0_i_2_1 (bank13_n_434),
        .\bdatw[12]_INST_0_i_2_2 (bank13_n_419),
        .\bdatw[13]_INST_0_i_16 (bank13_n_277),
        .\bdatw[13]_INST_0_i_16_0 (bank13_n_292),
        .\bdatw[13]_INST_0_i_16_1 (bank13_n_441),
        .\bdatw[13]_INST_0_i_16_2 (bank13_n_426),
        .\bdatw[13]_INST_0_i_2 (bank13_n_269),
        .\bdatw[13]_INST_0_i_2_0 (bank13_n_284),
        .\bdatw[13]_INST_0_i_2_1 (bank13_n_433),
        .\bdatw[13]_INST_0_i_2_2 (bank13_n_418),
        .\bdatw[14]_INST_0_i_16 (bank13_n_276),
        .\bdatw[14]_INST_0_i_16_0 (bank13_n_291),
        .\bdatw[14]_INST_0_i_16_1 (bank13_n_440),
        .\bdatw[14]_INST_0_i_16_2 (bank13_n_425),
        .\bdatw[14]_INST_0_i_2 (bank13_n_268),
        .\bdatw[14]_INST_0_i_2_0 (bank13_n_283),
        .\bdatw[14]_INST_0_i_2_1 (bank13_n_432),
        .\bdatw[14]_INST_0_i_2_2 (bank13_n_417),
        .\bdatw[15]_INST_0_i_15_0 ({p_0_in_2,\sp_reg[0] }),
        .\bdatw[15]_INST_0_i_15_1 (\rgf_c1bus_wb[4]_i_22 ),
        .\bdatw[15]_INST_0_i_16 (bank13_n_275),
        .\bdatw[15]_INST_0_i_16_0 (bank13_n_290),
        .\bdatw[15]_INST_0_i_16_1 (bank13_n_439),
        .\bdatw[15]_INST_0_i_16_2 (bank13_n_424),
        .\bdatw[15]_INST_0_i_2 (bank02_n_515),
        .\bdatw[15]_INST_0_i_2_0 (bank02_n_414),
        .\bdatw[15]_INST_0_i_2_1 (\tr_reg[15] ),
        .\bdatw[15]_INST_0_i_2_2 (bank13_n_267),
        .\bdatw[15]_INST_0_i_2_3 (bank13_n_416),
        .\bdatw[15]_INST_0_i_2_4 (\sr_reg[15] [15]),
        .\bdatw[8]_INST_0_i_16 (bank13_n_431),
        .\bdatw[8]_INST_0_i_16_0 (bank13_n_446),
        .\bdatw[8]_INST_0_i_16_1 (bank13_n_302),
        .\bdatw[8]_INST_0_i_16_2 (bank13_n_297),
        .\bdatw[8]_INST_0_i_16_3 (bank13_n_282),
        .\bdatw[8]_INST_0_i_2 (bank13_n_274),
        .\bdatw[8]_INST_0_i_2_0 (bank13_n_289),
        .\bdatw[8]_INST_0_i_2_1 (bank13_n_438),
        .\bdatw[8]_INST_0_i_2_2 (bank13_n_423),
        .\bdatw[9]_INST_0_i_16 (bank13_n_430),
        .\bdatw[9]_INST_0_i_16_0 (bank13_n_445),
        .\bdatw[9]_INST_0_i_16_1 (bank13_n_301),
        .\bdatw[9]_INST_0_i_16_2 (bank13_n_296),
        .\bdatw[9]_INST_0_i_16_3 (bank13_n_281),
        .\bdatw[9]_INST_0_i_2 (bank13_n_273),
        .\bdatw[9]_INST_0_i_2_0 (bank13_n_288),
        .\bdatw[9]_INST_0_i_2_1 (bank13_n_437),
        .\bdatw[9]_INST_0_i_2_2 (bank13_n_422),
        .data3(data3),
        .\iv_reg[15] (\iv_reg[15]_0 ),
        .out(\iv_reg[15] ),
        .\sp_reg[0] (\sp_reg[0]_2 ),
        .\sp_reg[10] (b1bus_out_n_6),
        .\sp_reg[11] (b1bus_out_n_5),
        .\sp_reg[12] (b1bus_out_n_4),
        .\sp_reg[13] (b1bus_out_n_3),
        .\sp_reg[14] (b1bus_out_n_2),
        .\sp_reg[1] (\sp_reg[1]_3 ),
        .\sp_reg[2] (\sp_reg[2]_2 ),
        .\sp_reg[3] (\sp_reg[3]_1 ),
        .\sp_reg[4] (\sp_reg[4]_2 ),
        .\sp_reg[5] (b1bus_out_n_11),
        .\sp_reg[6] (b1bus_out_n_10),
        .\sp_reg[7] (b1bus_out_n_9),
        .\sp_reg[8] (b1bus_out_n_8),
        .\sp_reg[9] (b1bus_out_n_7),
        .\sr_reg[0] (\sr_reg[0]_2 ),
        .\sr_reg[15] (\sr_reg[15]_1 ),
        .\sr_reg[1] (\sr_reg[1] ),
        .\sr_reg[2] (\sr_reg[2] ),
        .\sr_reg[3] (\sr_reg[3] ),
        .\sr_reg[4] (\sr_reg[4]_2 ),
        .\tr_reg[0] (\tr_reg[0]_0 ),
        .\tr_reg[10] (b1bus_out_n_27),
        .\tr_reg[11] (b1bus_out_n_28),
        .\tr_reg[12] (b1bus_out_n_29),
        .\tr_reg[13] (b1bus_out_n_30),
        .\tr_reg[14] (b1bus_out_n_31),
        .\tr_reg[1] (\tr_reg[1]_2 ),
        .\tr_reg[2] (\tr_reg[2]_0 ),
        .\tr_reg[3] (\tr_reg[3]_1 ),
        .\tr_reg[4] (\tr_reg[4]_0 ),
        .\tr_reg[5] (b1bus_out_n_22),
        .\tr_reg[6] (b1bus_out_n_23),
        .\tr_reg[7] (b1bus_out_n_24),
        .\tr_reg[8] (b1bus_out_n_25),
        .\tr_reg[9] (b1bus_out_n_26));
  mcss_rgf_bank bank02
       (.SR(SR),
        .a0bus_sel_0(a0bus_sel_0),
        .a1bus_sel_0({a1bus_sel_0[3:2],a1bus_sel_0[0]}),
        .b0bus_sel_0(b0bus_sel_0),
        .b1bus_b02(b1bus_b02),
        .\badr[0]_INST_0_i_1 (\badr[0]_INST_0_i_1 ),
        .\badr[10]_INST_0_i_1 (\badr[10]_INST_0_i_1 ),
        .\badr[10]_INST_0_i_1_0 (\badr[10]_INST_0_i_1_0 ),
        .\badr[10]_INST_0_i_1_1 (\badr[10]_INST_0_i_1_1 ),
        .\badr[10]_INST_0_i_1_2 (\badr[10]_INST_0_i_1_2 ),
        .\badr[10]_INST_0_i_2 (\badr[10]_INST_0_i_2 ),
        .\badr[10]_INST_0_i_2_0 (\badr[10]_INST_0_i_2_0 ),
        .\badr[11]_INST_0_i_1 (\badr[11]_INST_0_i_1 ),
        .\badr[11]_INST_0_i_2 (\badr[11]_INST_0_i_2 ),
        .\badr[12]_INST_0_i_1 (\badr[12]_INST_0_i_1 ),
        .\badr[12]_INST_0_i_2 (\badr[12]_INST_0_i_2 ),
        .\badr[12]_INST_0_i_2_0 (\badr[12]_INST_0_i_2_0 ),
        .\badr[13]_INST_0_i_1 (\badr[13]_INST_0_i_1 ),
        .\badr[13]_INST_0_i_1_0 (\badr[13]_INST_0_i_1_0 ),
        .\badr[13]_INST_0_i_2 (\badr[13]_INST_0_i_2 ),
        .\badr[13]_INST_0_i_2_0 (\badr[13]_INST_0_i_2_0 ),
        .\badr[14]_INST_0_i_1 (\badr[14]_INST_0_i_1 ),
        .\badr[14]_INST_0_i_1_0 (\badr[14]_INST_0_i_1_0 ),
        .\badr[14]_INST_0_i_1_1 (\badr[14]_INST_0_i_1_1 ),
        .\badr[14]_INST_0_i_2 (\badr[14]_INST_0_i_2 ),
        .\badr[14]_INST_0_i_2_0 (\badr[14]_INST_0_i_2_0 ),
        .\badr[14]_INST_0_i_2_1 (\badr[14]_INST_0_i_2_1 ),
        .\badr[14]_INST_0_i_2_2 (\badr[14]_INST_0_i_2_2 ),
        .\badr[15]_INST_0_i_1 (\badr[15]_INST_0_i_1 ),
        .\badr[15]_INST_0_i_1_0 (\badr[15]_INST_0_i_1_0 ),
        .\badr[15]_INST_0_i_1_1 (\badr[15]_INST_0_i_1_2 ),
        .\badr[1]_INST_0_i_1 (\badr[1]_INST_0_i_1 ),
        .\badr[1]_INST_0_i_2 (\badr[1]_INST_0_i_2 ),
        .\badr[1]_INST_0_i_2_0 (\badr[1]_INST_0_i_2_0 ),
        .\badr[2]_INST_0_i_1 (\badr[2]_INST_0_i_1 ),
        .\badr[2]_INST_0_i_1_0 (\badr[2]_INST_0_i_1_0 ),
        .\badr[2]_INST_0_i_1_1 (\badr[2]_INST_0_i_1_1 ),
        .\badr[2]_INST_0_i_2 (\badr[2]_INST_0_i_2 ),
        .\badr[2]_INST_0_i_2_0 (\badr[2]_INST_0_i_2_0 ),
        .\badr[3]_INST_0_i_1 (\badr[3]_INST_0_i_1 ),
        .\badr[3]_INST_0_i_1_0 (\badr[3]_INST_0_i_1_0 ),
        .\badr[3]_INST_0_i_2 (\badr[3]_INST_0_i_2 ),
        .\badr[3]_INST_0_i_2_0 (\badr[3]_INST_0_i_2_0 ),
        .\badr[4]_INST_0_i_2 (\badr[4]_INST_0_i_2 ),
        .\badr[4]_INST_0_i_2_0 (\badr[4]_INST_0_i_2_0 ),
        .\badr[5]_INST_0_i_1 (\badr[5]_INST_0_i_1 ),
        .\badr[5]_INST_0_i_1_0 (\badr[5]_INST_0_i_1_0 ),
        .\badr[5]_INST_0_i_2 (\badr[5]_INST_0_i_2 ),
        .\badr[5]_INST_0_i_2_0 (\badr[5]_INST_0_i_2_0 ),
        .\badr[6]_INST_0_i_1 (\badr[6]_INST_0_i_1 ),
        .\badr[6]_INST_0_i_1_0 (\badr[6]_INST_0_i_1_0 ),
        .\badr[6]_INST_0_i_1_1 (\badr[6]_INST_0_i_1_1 ),
        .\badr[6]_INST_0_i_1_2 (\badr[6]_INST_0_i_1_2 ),
        .\badr[6]_INST_0_i_1_3 (\badr[6]_INST_0_i_1_3 ),
        .\badr[6]_INST_0_i_2 (\badr[6]_INST_0_i_2 ),
        .\badr[6]_INST_0_i_2_0 (\badr[6]_INST_0_i_2_0 ),
        .\badr[6]_INST_0_i_2_1 (\badr[6]_INST_0_i_2_1 ),
        .\badr[7]_INST_0_i_1 (\badr[7]_INST_0_i_1 ),
        .\badr[7]_INST_0_i_2 (\badr[7]_INST_0_i_2 ),
        .\badr[8]_INST_0_i_2 (\badr[8]_INST_0_i_2 ),
        .\badr[8]_INST_0_i_2_0 (\badr[8]_INST_0_i_2_0 ),
        .\badr[8]_INST_0_i_2_1 (\badr[8]_INST_0_i_2_1 ),
        .\badr[9]_INST_0_i_1 (\badr[9]_INST_0_i_1 ),
        .\badr[9]_INST_0_i_1_0 (\badr[9]_INST_0_i_1_0 ),
        .\badr[9]_INST_0_i_2 (\badr[9]_INST_0_i_2 ),
        .\badr[9]_INST_0_i_2_0 (\badr[9]_INST_0_i_2_0 ),
        .bank_sel(bank_sel),
        .bbus_o(bbus_o),
        .\bbus_o[0]_INST_0_i_1 (sreg_n_38),
        .\bbus_o[0]_INST_0_i_1_0 (sreg_n_59),
        .\bbus_o[1]_INST_0_i_1 (sreg_n_37),
        .\bbus_o[1]_INST_0_i_1_0 (sreg_n_58),
        .\bbus_o[2]_INST_0_i_1 (sreg_n_36),
        .\bbus_o[2]_INST_0_i_1_0 (sreg_n_57),
        .\bbus_o[3]_INST_0_i_1 (sreg_n_35),
        .\bbus_o[3]_INST_0_i_1_0 (sreg_n_56),
        .\bbus_o[4]_INST_0_i_1 (sreg_n_34),
        .\bbus_o[4]_INST_0_i_1_0 (sreg_n_55),
        .\bbus_o[5] (\bbus_o[5] ),
        .\bbus_o[5]_0 (\bbus_o[5]_0 ),
        .\bbus_o[5]_1 (b0bus_out_n_21),
        .\bbus_o[5]_2 (b0bus_out_n_10),
        .\bbus_o[5]_3 (\bbus_o[5]_1 ),
        .\bbus_o[6] (\bbus_o[6] ),
        .\bbus_o[6]_0 (\bbus_o[6]_0 ),
        .\bbus_o[6]_1 (b0bus_out_n_22),
        .\bbus_o[6]_2 (b0bus_out_n_9),
        .\bbus_o[7] (\bbus_o[7] ),
        .\bbus_o[7]_0 (\bbus_o[7]_0 ),
        .\bbus_o[7]_1 (b0bus_out_n_23),
        .\bbus_o[7]_2 (b0bus_out_n_8),
        .bdatw(bdatw),
        .\bdatw[10] (\bdatw[10] ),
        .\bdatw[10]_0 (\bdatw[10]_0 ),
        .\bdatw[10]_1 (b1bus_out_n_27),
        .\bdatw[10]_2 (b1bus_out_n_6),
        .\bdatw[10]_3 (\bdatw[10]_1 ),
        .\bdatw[10]_4 (\bdatw[10]_2 ),
        .\bdatw[10]_5 (b0bus_out_n_26),
        .\bdatw[10]_6 (b0bus_out_n_5),
        .\bdatw[11] (\bdatw[11] ),
        .\bdatw[11]_0 (\bdatw[11]_0 ),
        .\bdatw[11]_1 (b1bus_out_n_28),
        .\bdatw[11]_2 (b1bus_out_n_5),
        .\bdatw[11]_3 (\bdatw[11]_1 ),
        .\bdatw[11]_4 (\bdatw[11]_2 ),
        .\bdatw[11]_5 (b0bus_out_n_27),
        .\bdatw[11]_6 (b0bus_out_n_4),
        .\bdatw[12] (\bdatw[12] ),
        .\bdatw[12]_0 (\bdatw[12]_0 ),
        .\bdatw[12]_1 (b1bus_out_n_29),
        .\bdatw[12]_2 (b1bus_out_n_4),
        .\bdatw[12]_3 (\bdatw[12]_1 ),
        .\bdatw[12]_4 (\bdatw[12]_2 ),
        .\bdatw[12]_5 (b0bus_out_n_28),
        .\bdatw[12]_6 (b0bus_out_n_3),
        .\bdatw[13] (\bdatw[13] ),
        .\bdatw[13]_0 (\bdatw[13]_0 ),
        .\bdatw[13]_1 (\bdatw[13]_1 ),
        .\bdatw[13]_2 (\bdatw[13]_2 ),
        .\bdatw[13]_3 (\bdatw[13]_3 ),
        .\bdatw[13]_4 (b1bus_out_n_30),
        .\bdatw[13]_5 (b1bus_out_n_3),
        .\bdatw[13]_6 (\bdatw[13]_4 ),
        .\bdatw[13]_7 (\bdatw[13]_5 ),
        .\bdatw[13]_8 (b0bus_out_n_29),
        .\bdatw[13]_9 (b0bus_out_n_2),
        .\bdatw[14] (\bdatw[14] ),
        .\bdatw[14]_0 (\bdatw[14]_0 ),
        .\bdatw[14]_1 (b1bus_out_n_31),
        .\bdatw[14]_2 (b1bus_out_n_2),
        .\bdatw[14]_3 (\bdatw[14]_1 ),
        .\bdatw[14]_4 (\bdatw[14]_2 ),
        .\bdatw[14]_5 (b0bus_out_n_30),
        .\bdatw[14]_6 (b0bus_out_n_1),
        .\bdatw[15] (\bdatw[15] ),
        .\bdatw[15]_0 (\bdatw[15]_0 ),
        .\bdatw[15]_1 (b0bus_out_n_31),
        .\bdatw[15]_2 (b0bus_out_n_0),
        .\bdatw[8] (\bdatw[8] ),
        .\bdatw[8]_0 (\bdatw[8]_0 ),
        .\bdatw[8]_1 (b1bus_out_n_25),
        .\bdatw[8]_2 (b1bus_out_n_8),
        .\bdatw[8]_3 (\bdatw[8]_1 ),
        .\bdatw[8]_4 (\bdatw[8]_2 ),
        .\bdatw[8]_5 (b0bus_out_n_24),
        .\bdatw[8]_6 (b0bus_out_n_7),
        .\bdatw[9] (\bdatw[9] ),
        .\bdatw[9]_0 (\bdatw[9]_0 ),
        .\bdatw[9]_1 (b1bus_out_n_26),
        .\bdatw[9]_2 (b1bus_out_n_7),
        .\bdatw[9]_3 (\bdatw[9]_1 ),
        .\bdatw[9]_4 (\bdatw[9]_2 ),
        .\bdatw[9]_5 (b0bus_out_n_25),
        .\bdatw[9]_6 (b0bus_out_n_6),
        .clk(clk),
        .ctl_sela0(ctl_sela0),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .gr6_bus1(\a1buso2l/gr6_bus1 ),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (bank02_n_361),
        .\grn_reg[0]_1 (bank02_n_362),
        .\grn_reg[0]_2 (bank02_n_412),
        .\grn_reg[0]_3 (bank02_n_413),
        .\grn_reg[0]_4 (\grn_reg[0]_0 ),
        .\grn_reg[0]_5 (bank02_n_446),
        .\grn_reg[0]_6 (bank02_n_462),
        .\grn_reg[0]_7 (bank02_n_498),
        .\grn_reg[0]_8 (bank02_n_514),
        .\grn_reg[10] (bank02_n_340),
        .\grn_reg[10]_0 (bank02_n_341),
        .\grn_reg[10]_1 (bank02_n_394),
        .\grn_reg[10]_2 (bank02_n_395),
        .\grn_reg[10]_3 (bank02_n_435),
        .\grn_reg[10]_4 (bank02_n_452),
        .\grn_reg[10]_5 (bank02_n_489),
        .\grn_reg[10]_6 (bank02_n_505),
        .\grn_reg[11] (bank02_n_338),
        .\grn_reg[11]_0 (bank02_n_339),
        .\grn_reg[11]_1 (bank02_n_392),
        .\grn_reg[11]_2 (bank02_n_393),
        .\grn_reg[11]_3 (bank02_n_434),
        .\grn_reg[11]_4 (bank02_n_451),
        .\grn_reg[11]_5 (bank02_n_488),
        .\grn_reg[11]_6 (bank02_n_504),
        .\grn_reg[12] (bank02_n_336),
        .\grn_reg[12]_0 (bank02_n_337),
        .\grn_reg[12]_1 (bank02_n_390),
        .\grn_reg[12]_2 (bank02_n_391),
        .\grn_reg[12]_3 (bank02_n_433),
        .\grn_reg[12]_4 (bank02_n_450),
        .\grn_reg[12]_5 (bank02_n_487),
        .\grn_reg[12]_6 (bank02_n_503),
        .\grn_reg[13] (bank02_n_334),
        .\grn_reg[13]_0 (bank02_n_335),
        .\grn_reg[13]_1 (bank02_n_388),
        .\grn_reg[13]_2 (bank02_n_389),
        .\grn_reg[13]_3 (bank02_n_432),
        .\grn_reg[13]_4 (bank02_n_449),
        .\grn_reg[13]_5 (bank02_n_486),
        .\grn_reg[13]_6 (bank02_n_502),
        .\grn_reg[14] ({a1bus_b02[14:8],a1bus_b02[6],a1bus_b02[4:0]}),
        .\grn_reg[14]_0 (bank02_n_332),
        .\grn_reg[14]_1 (bank02_n_333),
        .\grn_reg[14]_2 (bank02_n_386),
        .\grn_reg[14]_3 (bank02_n_387),
        .\grn_reg[14]_4 (bank02_n_431),
        .\grn_reg[14]_5 (bank02_n_448),
        .\grn_reg[14]_6 (bank02_n_485),
        .\grn_reg[14]_7 (bank02_n_501),
        .\grn_reg[15] ({bank02_n_20,bank02_n_21,bank02_n_22,bank02_n_23,bank02_n_24,bank02_n_25,bank02_n_26,bank02_n_27,bank02_n_28,bank02_n_29,bank02_n_30,bank02_n_31,bank02_n_32,bank02_n_33,bank02_n_34,bank02_n_35}),
        .\grn_reg[15]_0 ({bank02_n_36,bank02_n_37,bank02_n_38,bank02_n_39,bank02_n_40,bank02_n_41,bank02_n_42,bank02_n_43,bank02_n_44,bank02_n_45,bank02_n_46,bank02_n_47,bank02_n_48,bank02_n_49,bank02_n_50,bank02_n_51}),
        .\grn_reg[15]_1 ({bank02_n_57,bank02_n_58,bank02_n_59,bank02_n_60,bank02_n_61,bank02_n_62,bank02_n_63,bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72}),
        .\grn_reg[15]_10 (bank02_n_447),
        .\grn_reg[15]_11 (bank02_n_484),
        .\grn_reg[15]_12 (bank02_n_499),
        .\grn_reg[15]_13 (bank02_n_515),
        .\grn_reg[15]_14 (\grn_reg[15]_2 ),
        .\grn_reg[15]_15 (\grn_reg[15]_3 ),
        .\grn_reg[15]_16 (\grn_reg[15]_4 ),
        .\grn_reg[15]_17 (\grn_reg[15]_5 ),
        .\grn_reg[15]_18 (\grn_reg[15]_6 ),
        .\grn_reg[15]_19 (\grn_reg[15]_7 ),
        .\grn_reg[15]_2 ({bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78,bank02_n_79,bank02_n_80,bank02_n_81,bank02_n_82,bank02_n_83,bank02_n_84,bank02_n_85,bank02_n_86,bank02_n_87,bank02_n_88}),
        .\grn_reg[15]_20 (\grn_reg[15]_8 ),
        .\grn_reg[15]_21 (\grn_reg[15]_9 ),
        .\grn_reg[15]_22 (\grn_reg[15]_10 ),
        .\grn_reg[15]_23 (\grn_reg[15]_11 ),
        .\grn_reg[15]_24 (\grn_reg[15]_12 ),
        .\grn_reg[15]_25 (\grn_reg[15]_13 ),
        .\grn_reg[15]_26 (\grn_reg[15]_14 ),
        .\grn_reg[15]_27 (\grn_reg[15]_15 ),
        .\grn_reg[15]_28 (\grn_reg[15]_16 ),
        .\grn_reg[15]_29 (\grn_reg[15]_17 ),
        .\grn_reg[15]_3 (\grn_reg[15]_1 ),
        .\grn_reg[15]_30 (\grn_reg[15]_18 ),
        .\grn_reg[15]_31 (\grn_reg[15]_19 ),
        .\grn_reg[15]_32 (\grn_reg[15]_20 ),
        .\grn_reg[15]_33 (\grn_reg[15]_21 ),
        .\grn_reg[15]_34 (\grn_reg[15]_22 ),
        .\grn_reg[15]_35 (\grn_reg[15]_23 ),
        .\grn_reg[15]_36 (\grn_reg[15]_24 ),
        .\grn_reg[15]_37 (\grn_reg[15]_25 ),
        .\grn_reg[15]_38 (\grn_reg[15]_26 ),
        .\grn_reg[15]_39 (\grn_reg[15]_27 ),
        .\grn_reg[15]_4 (bank02_n_330),
        .\grn_reg[15]_40 (\grn_reg[15]_28 ),
        .\grn_reg[15]_41 (\grn_reg[15]_29 ),
        .\grn_reg[15]_42 (\grn_reg[15]_30 ),
        .\grn_reg[15]_43 (\grn_reg[15]_31 ),
        .\grn_reg[15]_44 (\grn_reg[15]_32 ),
        .\grn_reg[15]_45 (\grn_reg[15]_33 ),
        .\grn_reg[15]_5 (bank02_n_331),
        .\grn_reg[15]_6 (bank02_n_384),
        .\grn_reg[15]_7 (bank02_n_385),
        .\grn_reg[15]_8 (bank02_n_414),
        .\grn_reg[15]_9 (bank02_n_430),
        .\grn_reg[1] (bank02_n_358),
        .\grn_reg[1]_0 (bank02_n_359),
        .\grn_reg[1]_1 (bank02_n_410),
        .\grn_reg[1]_2 (bank02_n_411),
        .\grn_reg[1]_3 (bank02_n_444),
        .\grn_reg[1]_4 (bank02_n_461),
        .\grn_reg[1]_5 (bank02_n_497),
        .\grn_reg[1]_6 (bank02_n_513),
        .\grn_reg[2] (bank02_n_356),
        .\grn_reg[2]_0 (bank02_n_357),
        .\grn_reg[2]_1 (bank02_n_408),
        .\grn_reg[2]_2 (bank02_n_409),
        .\grn_reg[2]_3 (bank02_n_443),
        .\grn_reg[2]_4 (bank02_n_460),
        .\grn_reg[2]_5 (bank02_n_496),
        .\grn_reg[2]_6 (bank02_n_512),
        .\grn_reg[3] (bank02_n_354),
        .\grn_reg[3]_0 (bank02_n_355),
        .\grn_reg[3]_1 (bank02_n_406),
        .\grn_reg[3]_2 (bank02_n_407),
        .\grn_reg[3]_3 (bank02_n_442),
        .\grn_reg[3]_4 (bank02_n_459),
        .\grn_reg[3]_5 (bank02_n_495),
        .\grn_reg[3]_6 (bank02_n_511),
        .\grn_reg[4] ({bank02_n_15,bank02_n_16,bank02_n_17,bank02_n_18,bank02_n_19}),
        .\grn_reg[4]_0 ({bank02_n_52,bank02_n_53,bank02_n_54,bank02_n_55,bank02_n_56}),
        .\grn_reg[4]_1 (bank02_n_352),
        .\grn_reg[4]_10 (bank02_n_510),
        .\grn_reg[4]_2 (bank02_n_353),
        .\grn_reg[4]_3 (\grn_reg[4]_8 ),
        .\grn_reg[4]_4 (bank02_n_404),
        .\grn_reg[4]_5 (bank02_n_405),
        .\grn_reg[4]_6 (bank02_n_441),
        .\grn_reg[4]_7 (bank02_n_458),
        .\grn_reg[4]_8 (\grn_reg[4]_9 ),
        .\grn_reg[4]_9 (bank02_n_494),
        .\grn_reg[5] (bank02_n_350),
        .\grn_reg[5]_0 (bank02_n_351),
        .\grn_reg[5]_1 (bank02_n_402),
        .\grn_reg[5]_2 (bank02_n_403),
        .\grn_reg[5]_3 (bank02_n_440),
        .\grn_reg[5]_4 (bank02_n_457),
        .\grn_reg[5]_5 (bank02_n_493),
        .\grn_reg[5]_6 (bank02_n_509),
        .\grn_reg[6] (bank02_n_348),
        .\grn_reg[6]_0 (bank02_n_349),
        .\grn_reg[6]_1 (bank02_n_400),
        .\grn_reg[6]_2 (bank02_n_401),
        .\grn_reg[6]_3 (bank02_n_439),
        .\grn_reg[6]_4 (bank02_n_456),
        .\grn_reg[6]_5 (bank02_n_492),
        .\grn_reg[6]_6 (bank02_n_508),
        .\grn_reg[7] (bank02_n_346),
        .\grn_reg[7]_0 (bank02_n_347),
        .\grn_reg[7]_1 (bank02_n_398),
        .\grn_reg[7]_2 (bank02_n_399),
        .\grn_reg[7]_3 (bank02_n_438),
        .\grn_reg[7]_4 (bank02_n_455),
        .\grn_reg[7]_5 (bank02_n_491),
        .\grn_reg[7]_6 (bank02_n_507),
        .\grn_reg[8] (bank02_n_344),
        .\grn_reg[8]_0 (bank02_n_345),
        .\grn_reg[8]_1 (bank02_n_437),
        .\grn_reg[8]_2 (bank02_n_454),
        .\grn_reg[9] (bank02_n_342),
        .\grn_reg[9]_0 (bank02_n_343),
        .\grn_reg[9]_1 (bank02_n_396),
        .\grn_reg[9]_2 (bank02_n_397),
        .\grn_reg[9]_3 (bank02_n_436),
        .\grn_reg[9]_4 (bank02_n_453),
        .\grn_reg[9]_5 (bank02_n_490),
        .\grn_reg[9]_6 (bank02_n_506),
        .\i_/badr[15]_INST_0_i_19 (\i_/badr[15]_INST_0_i_19 ),
        .\i_/badr[15]_INST_0_i_19_0 (\i_/badr[15]_INST_0_i_19_0 ),
        .\i_/badr[15]_INST_0_i_19_1 (\i_/badr[15]_INST_0_i_19_1 ),
        .\i_/badr[15]_INST_0_i_43 (\i_/badr[15]_INST_0_i_43 ),
        .\i_/badr[15]_INST_0_i_43_0 (\i_/badr[15]_INST_0_i_43_0 ),
        .\i_/badr[15]_INST_0_i_47 (sreg_n_95),
        .\i_/bdatw[15]_INST_0_i_112 (\i_/bdatw[15]_INST_0_i_112 ),
        .\i_/bdatw[15]_INST_0_i_112_0 (\i_/bdatw[15]_INST_0_i_112_0 ),
        .\i_/bdatw[15]_INST_0_i_112_1 (\i_/bdatw[15]_INST_0_i_112_1 ),
        .\i_/bdatw[15]_INST_0_i_113 (\i_/bdatw[15]_INST_0_i_113 ),
        .\i_/bdatw[15]_INST_0_i_24 (\i_/bdatw[15]_INST_0_i_24 ),
        .\i_/bdatw[15]_INST_0_i_24_0 (\i_/bdatw[15]_INST_0_i_24_0 ),
        .\i_/bdatw[15]_INST_0_i_44 (\i_/bdatw[15]_INST_0_i_44 ),
        .\i_/bdatw[15]_INST_0_i_77 (\i_/bdatw[15]_INST_0_i_77 ),
        .\i_/bdatw[15]_INST_0_i_9 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_9_0 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .\i_/bdatw[15]_INST_0_i_9_1 (\i_/bdatw[15]_INST_0_i_9_1 ),
        .\i_/bdatw[15]_INST_0_i_9_2 (\i_/bdatw[15]_INST_0_i_9_2 ),
        .\i_/bdatw[15]_INST_0_i_9_3 (\i_/bdatw[15]_INST_0_i_9_3 ),
        .out(out),
        .p_0_in(p_0_in),
        .p_0_in0_in(p_0_in0_in),
        .p_1_in(p_1_in),
        .p_1_in1_in(p_1_in1_in),
        .\rgf_c0bus_wb[0]_i_14 (\rgf_c0bus_wb[0]_i_14 ),
        .\rgf_c0bus_wb[10]_i_4 (\rgf_c0bus_wb[10]_i_4 ),
        .\rgf_c0bus_wb[10]_i_8 (\rgf_c0bus_wb[10]_i_8 ),
        .\rgf_c0bus_wb[11]_i_11 (\rgf_c0bus_wb[11]_i_11 ),
        .\rgf_c0bus_wb[11]_i_11_0 (\rgf_c0bus_wb[11]_i_11_0 ),
        .\rgf_c0bus_wb[11]_i_11_1 (\rgf_c0bus_wb[11]_i_11_1 ),
        .\rgf_c0bus_wb[11]_i_11_2 (\rgf_c0bus_wb[11]_i_11_2 ),
        .\rgf_c0bus_wb[11]_i_22 (\rgf_c0bus_wb[11]_i_22 ),
        .\rgf_c0bus_wb[11]_i_22_0 (\rgf_c0bus_wb[11]_i_22_0 ),
        .\rgf_c0bus_wb[11]_i_3 (\rgf_c0bus_wb[11]_i_3 ),
        .\rgf_c0bus_wb[11]_i_3_0 (\rgf_c0bus_wb[11]_i_3_0 ),
        .\rgf_c0bus_wb[11]_i_3_1 (\rgf_c0bus_wb[11]_i_3_1 ),
        .\rgf_c0bus_wb[11]_i_3_2 (\rgf_c0bus_wb[11]_i_3_2 ),
        .\rgf_c0bus_wb[11]_i_3_3 (\rgf_c0bus_wb[11]_i_3_3 ),
        .\rgf_c0bus_wb[11]_i_8 (\rgf_c0bus_wb[11]_i_8 ),
        .\rgf_c0bus_wb[11]_i_9 (\rgf_c0bus_wb[11]_i_9_1 ),
        .\rgf_c0bus_wb[11]_i_9_0 (\rgf_c0bus_wb[11]_i_9_0 ),
        .\rgf_c0bus_wb[11]_i_9_1 (\rgf_c0bus_wb[11]_i_9_2 ),
        .\rgf_c0bus_wb[11]_i_9_2 (\rgf_c0bus_wb[11]_i_9_3 ),
        .\rgf_c0bus_wb[11]_i_9_3 (\rgf_c0bus_wb[11]_i_9 ),
        .\rgf_c0bus_wb[11]_i_9_4 (\rgf_c0bus_wb[11]_i_9_4 ),
        .\rgf_c0bus_wb[12]_i_10 (a0bus_0[15]),
        .\rgf_c0bus_wb[12]_i_2 (\rgf_c0bus_wb[12]_i_2 ),
        .\rgf_c0bus_wb[12]_i_22_0 (bank02_n_264),
        .\rgf_c0bus_wb[12]_i_24 (\rgf_c0bus_wb[12]_i_24 ),
        .\rgf_c0bus_wb[12]_i_25_0 (\rgf_c0bus_wb[12]_i_25 ),
        .\rgf_c0bus_wb[12]_i_7 (bank13_n_164),
        .\rgf_c0bus_wb[13]_i_28 (\rgf_c0bus_wb[13]_i_28 ),
        .\rgf_c0bus_wb[13]_i_29 (\rgf_c0bus_wb[13]_i_29 ),
        .\rgf_c0bus_wb[13]_i_4 (\rgf_c0bus_wb[13]_i_4 ),
        .\rgf_c0bus_wb[14]_i_13 (a0bus_0[7]),
        .\rgf_c0bus_wb[14]_i_13_0 (a0bus_0[11]),
        .\rgf_c0bus_wb[14]_i_13_1 (a0bus_0[9]),
        .\rgf_c0bus_wb[14]_i_13_2 (a0bus_0[8]),
        .\rgf_c0bus_wb[14]_i_13_3 (a0bus_0[10]),
        .\rgf_c0bus_wb[14]_i_13_4 (a0bus_0[13]),
        .\rgf_c0bus_wb[14]_i_13_5 (a0bus_0[12]),
        .\rgf_c0bus_wb[14]_i_13_6 (a0bus_0[14]),
        .\rgf_c0bus_wb[14]_i_2 (\rgf_c0bus_wb[14]_i_2 ),
        .\rgf_c0bus_wb[15]_i_14 (\rgf_c0bus_wb[15]_i_14 ),
        .\rgf_c0bus_wb[15]_i_18 (\rgf_c0bus_wb[15]_i_18 ),
        .\rgf_c0bus_wb[15]_i_25_0 (\rgf_c0bus_wb[15]_i_25 ),
        .\rgf_c0bus_wb[15]_i_26 (\rgf_c0bus_wb[15]_i_26 ),
        .\rgf_c0bus_wb[15]_i_6 (\rgf_c0bus_wb[15]_i_6 ),
        .\rgf_c0bus_wb[15]_i_6_0 (\rgf_c0bus_wb[15]_i_6_0 ),
        .\rgf_c0bus_wb[15]_i_6_1 (\rgf_c0bus_wb[15]_i_6_1 ),
        .\rgf_c0bus_wb[3]_i_18 (a0bus_0[6]),
        .\rgf_c0bus_wb[3]_i_18_0 (a0bus_0[5]),
        .\rgf_c0bus_wb[3]_i_7 (a0bus_0[3]),
        .\rgf_c0bus_wb[3]_i_7_0 (\rgf_c0bus_wb[3]_i_7 ),
        .\rgf_c0bus_wb[3]_i_7_1 (\rgf_c0bus_wb[3]_i_7_0 ),
        .\rgf_c0bus_wb[3]_i_7_2 (a0bus_0[1]),
        .\rgf_c0bus_wb[3]_i_7_3 (a0bus_0[0]),
        .\rgf_c0bus_wb[3]_i_7_4 (a0bus_0[2]),
        .\rgf_c0bus_wb[4]_i_3 (bank13_n_156),
        .\rgf_c0bus_wb[4]_i_7 (a0bus_out_n_7),
        .\rgf_c0bus_wb[4]_i_7_0 (a0bus_out_n_3),
        .\rgf_c0bus_wb[4]_i_7_1 (a0bus_out_n_1),
        .\rgf_c0bus_wb[4]_i_7_2 (a0bus_out_n_2),
        .\rgf_c0bus_wb[4]_i_7_3 (a0bus_out_n_65),
        .\rgf_c0bus_wb[6]_i_11 (\rgf_c0bus_wb[6]_i_11 ),
        .\rgf_c0bus_wb[7]_i_7 (\rgf_c0bus_wb[7]_i_7 ),
        .\rgf_c0bus_wb[7]_i_7_0 (\rgf_c0bus_wb[7]_i_7_0 ),
        .\rgf_c0bus_wb[8]_i_2 (a0bus_0[4]),
        .\rgf_c0bus_wb[8]_i_6_0 (\rgf_c0bus_wb[8]_i_6 ),
        .\rgf_c0bus_wb_reg[10] (\rgf_c0bus_wb_reg[10]_1 ),
        .\rgf_c0bus_wb_reg[10]_0 (\rgf_c0bus_wb_reg[10] ),
        .\rgf_c0bus_wb_reg[10]_1 (\rgf_c0bus_wb_reg[10]_0 ),
        .\rgf_c0bus_wb_reg[7]_i_11 (\rgf_c0bus_wb_reg[7]_i_11 ),
        .\rgf_c1bus_wb[11]_i_10 (\rgf_c1bus_wb[11]_i_10 ),
        .\rgf_c1bus_wb[11]_i_10_0 (\rgf_c1bus_wb[11]_i_10_0 ),
        .\rgf_c1bus_wb[11]_i_10_1 (\rgf_c1bus_wb[11]_i_10_1 ),
        .\rgf_c1bus_wb[11]_i_10_2 (\rgf_c1bus_wb[11]_i_10_2 ),
        .\rgf_c1bus_wb[11]_i_10_3 (\rgf_c1bus_wb[11]_i_10_3 ),
        .\rgf_c1bus_wb[11]_i_10_4 (\rgf_c1bus_wb[11]_i_10_4 ),
        .\rgf_c1bus_wb[11]_i_10_5 (\rgf_c1bus_wb[11]_i_10_5 ),
        .\rgf_c1bus_wb[11]_i_13 (\rgf_c1bus_wb[11]_i_13 ),
        .\rgf_c1bus_wb[12]_i_2 (\rgf_c1bus_wb[12]_i_2 ),
        .\rgf_c1bus_wb[12]_i_20_0 (\rgf_c1bus_wb[12]_i_20 ),
        .\rgf_c1bus_wb[13]_i_16 (\rgf_c1bus_wb[13]_i_16 ),
        .\rgf_c1bus_wb[13]_i_9 (\rgf_c1bus_wb[13]_i_9 ),
        .\rgf_c1bus_wb[14]_i_11 (\rgf_c1bus_wb[14]_i_11 ),
        .\rgf_c1bus_wb[14]_i_11_0 (\rgf_c1bus_wb[14]_i_11_0 ),
        .\rgf_c1bus_wb[14]_i_11_1 (b1bus_out_n_23),
        .\rgf_c1bus_wb[14]_i_11_2 (b1bus_out_n_10),
        .\rgf_c1bus_wb[14]_i_28 (\rgf_c1bus_wb[14]_i_28 ),
        .\rgf_c1bus_wb[14]_i_28_0 (\rgf_c1bus_wb[14]_i_28_0 ),
        .\rgf_c1bus_wb[14]_i_28_1 (\rgf_c1bus_wb[14]_i_28_1 ),
        .\rgf_c1bus_wb[14]_i_28_2 (\rgf_c1bus_wb[14]_i_28_2 ),
        .\rgf_c1bus_wb[14]_i_28_3 (\rgf_c1bus_wb[14]_i_28_4 ),
        .\rgf_c1bus_wb[14]_i_28_4 (\rgf_c1bus_wb[14]_i_28_5 ),
        .\rgf_c1bus_wb[14]_i_28_5 (\rgf_c1bus_wb[14]_i_28_6 ),
        .\rgf_c1bus_wb[14]_i_28_6 (\rgf_c1bus_wb[14]_i_28_7 ),
        .\rgf_c1bus_wb[14]_i_30 (\rgf_c1bus_wb[14]_i_30 ),
        .\rgf_c1bus_wb[14]_i_32 (\rgf_c1bus_wb[14]_i_32 ),
        .\rgf_c1bus_wb[14]_i_32_0 (\rgf_c1bus_wb[14]_i_32_0 ),
        .\rgf_c1bus_wb[15]_i_14 (\rgf_c1bus_wb[15]_i_14 ),
        .\rgf_c1bus_wb[15]_i_14_0 (\rgf_c1bus_wb[15]_i_14_0 ),
        .\rgf_c1bus_wb[15]_i_14_1 (\rgf_c1bus_wb[15]_i_14_1 ),
        .\rgf_c1bus_wb[15]_i_14_2 (\rgf_c1bus_wb[15]_i_14_2 ),
        .\rgf_c1bus_wb[15]_i_14_3 (\rgf_c1bus_wb[15]_i_14_3 ),
        .\rgf_c1bus_wb[15]_i_19 (\rgf_c1bus_wb[15]_i_19 ),
        .\rgf_c1bus_wb[15]_i_19_0 (\rgf_c1bus_wb[15]_i_19_0 ),
        .\rgf_c1bus_wb[15]_i_19_1 (b1bus_out_n_24),
        .\rgf_c1bus_wb[15]_i_19_2 (b1bus_out_n_9),
        .\rgf_c1bus_wb[15]_i_27 (\rgf_c1bus_wb[15]_i_27 ),
        .\rgf_c1bus_wb[1]_i_14_0 (\rgf_c1bus_wb[1]_i_14 ),
        .\rgf_c1bus_wb[4]_i_22 (sreg_n_96),
        .\rgf_c1bus_wb[4]_i_22_0 (sreg_n_127),
        .\rgf_c1bus_wb[4]_i_23 (sreg_n_97),
        .\rgf_c1bus_wb[4]_i_23_0 (sreg_n_126),
        .\rgf_c1bus_wb[4]_i_24 (sreg_n_99),
        .\rgf_c1bus_wb[4]_i_24_0 (sreg_n_124),
        .\rgf_c1bus_wb[4]_i_25 (sreg_n_107),
        .\rgf_c1bus_wb[4]_i_25_0 (sreg_n_116),
        .\rgf_c1bus_wb[4]_i_26 (sreg_n_105),
        .\rgf_c1bus_wb[4]_i_26_0 (sreg_n_118),
        .\rgf_c1bus_wb[4]_i_27 (sreg_n_103),
        .\rgf_c1bus_wb[4]_i_27_0 (sreg_n_120),
        .\rgf_c1bus_wb[4]_i_28 (sreg_n_101),
        .\rgf_c1bus_wb[4]_i_28_0 (sreg_n_122),
        .\rgf_c1bus_wb[4]_i_33 (\rgf_c1bus_wb[4]_i_33 ),
        .\rgf_c1bus_wb[4]_i_33_0 (sreg_n_87),
        .\rgf_c1bus_wb[4]_i_37 (\rgf_c1bus_wb[4]_i_37 ),
        .\rgf_c1bus_wb[4]_i_37_0 (sreg_n_89),
        .\rgf_c1bus_wb[4]_i_41 (\rgf_c1bus_wb[4]_i_41 ),
        .\rgf_c1bus_wb[4]_i_41_0 (sreg_n_77),
        .\rgf_c1bus_wb[4]_i_47 (\rgf_c1bus_wb[4]_i_47 ),
        .\rgf_c1bus_wb[4]_i_47_0 (sreg_n_76),
        .\rgf_c1bus_wb[4]_i_51 (\rgf_c1bus_wb[4]_i_51 ),
        .\rgf_c1bus_wb[4]_i_51_0 (sreg_n_78),
        .\rgf_c1bus_wb[4]_i_53 (\rgf_c1bus_wb[4]_i_53 ),
        .\rgf_c1bus_wb[4]_i_53_0 (sreg_n_85),
        .\rgf_c1bus_wb[4]_i_57 (\rgf_c1bus_wb[4]_i_57 ),
        .\rgf_c1bus_wb[4]_i_57_0 (sreg_n_83),
        .\rgf_c1bus_wb[4]_i_61 (\rgf_c1bus_wb[4]_i_61 ),
        .\rgf_c1bus_wb[4]_i_61_0 (sreg_n_82),
        .\rgf_c1bus_wb[4]_i_65 (\rgf_c1bus_wb[4]_i_65 ),
        .\rgf_c1bus_wb[4]_i_65_0 (sreg_n_80),
        .\rgf_c1bus_wb[4]_i_67 (\rgf_c1bus_wb[4]_i_67 ),
        .\rgf_c1bus_wb[4]_i_67_0 (sreg_n_88),
        .\rgf_c1bus_wb[4]_i_7 (\tr_reg[15]_0 ),
        .\rgf_c1bus_wb[4]_i_7_0 (a1bus_out_n_49),
        .\rgf_c1bus_wb[4]_i_7_1 (a1bus_out_n_6),
        .\rgf_c1bus_wb[4]_i_9 (\rgf_c1bus_wb[4]_i_9 ),
        .\rgf_c1bus_wb[4]_i_9_0 (\rgf_c1bus_wb[4]_i_9_0 ),
        .\rgf_c1bus_wb[5]_i_10 (\rgf_c1bus_wb[5]_i_10 ),
        .\rgf_c1bus_wb[7]_i_4 (\rgf_c1bus_wb[7]_i_4 ),
        .\rgf_c1bus_wb[7]_i_4_0 (\rgf_c1bus_wb[7]_i_4_0 ),
        .\rgf_c1bus_wb[9]_i_17_0 (\rgf_c1bus_wb[9]_i_17 ),
        .\rgf_c1bus_wb_reg[10] (\rgf_c1bus_wb_reg[10] ),
        .\rgf_c1bus_wb_reg[3] (\rgf_c1bus_wb_reg[3] ),
        .\rgf_c1bus_wb_reg[4] (\rgf_c1bus_wb_reg[4] ),
        .\rgf_c1bus_wb_reg[5] (\rgf_c1bus_wb_reg[5] ),
        .\rgf_c1bus_wb_reg[5]_0 (\rgf_c1bus_wb_reg[5]_0 ),
        .\rgf_c1bus_wb_reg[5]_1 (\rgf_c1bus_wb_reg[5]_1 ),
        .\rgf_c1bus_wb_reg[7] (\rgf_c1bus_wb_reg[7] ),
        .\sr[4]_i_102 (a1bus_0[11]),
        .\sr[4]_i_102_0 (bank13_n_138),
        .\sr[4]_i_111 (\tr_reg[3] ),
        .\sr[4]_i_119 (\sr_reg[6]_6 ),
        .\sr[4]_i_126 (\sr_reg[6]_33 ),
        .\sr[4]_i_139 (\sp_reg[4]_0 ),
        .\sr[4]_i_169_0 (a1bus_out_n_23),
        .\sr[4]_i_169_1 (a1bus_out_n_57),
        .\sr[4]_i_169_2 (a1bus_out_n_26),
        .\sr[4]_i_169_3 (a1bus_out_n_17),
        .\sr[4]_i_169_4 (a1bus_out_n_55),
        .\sr[4]_i_169_5 (a1bus_out_n_21),
        .\sr[4]_i_169_6 (a1bus_out_n_56),
        .\sr[4]_i_169_7 (a1bus_out_n_28),
        .\sr[4]_i_169_8 (a1bus_out_n_32),
        .\sr[4]_i_171 (a1bus_out_n_5),
        .\sr[4]_i_171_0 (a1bus_out_n_51),
        .\sr[4]_i_171_1 (a1bus_out_n_9),
        .\sr[4]_i_171_2 (a1bus_out_n_52),
        .\sr[4]_i_175_0 (a1bus_out_n_34),
        .\sr[4]_i_175_1 (a1bus_out_n_38),
        .\sr[4]_i_175_2 (a1bus_out_n_62),
        .\sr[4]_i_175_3 (a1bus_out_n_40),
        .\sr[4]_i_175_4 (a1bus_out_n_63),
        .\sr[4]_i_175_5 (a1bus_out_n_44),
        .\sr[4]_i_175_6 (a1bus_out_n_64),
        .\sr[4]_i_177 (a1bus_out_n_11),
        .\sr[4]_i_177_0 (a1bus_out_n_53),
        .\sr[4]_i_177_1 (a1bus_out_n_15),
        .\sr[4]_i_177_2 (a1bus_out_n_54),
        .\sr[4]_i_179_0 (a1bus_out_n_58),
        .\sr[4]_i_179_1 (a1bus_out_n_61),
        .\sr[4]_i_179_2 (a1bus_out_n_59),
        .\sr[4]_i_179_3 (a1bus_out_n_60),
        .\sr[4]_i_179_4 (a1bus_out_n_31),
        .\sr[4]_i_179_5 (a1bus_out_n_35),
        .\sr[4]_i_179_6 (a1bus_out_n_25),
        .\sr[4]_i_179_7 (a1bus_out_n_29),
        .\sr[4]_i_188 (a0bus_out_n_5),
        .\sr[4]_i_188_0 (a0bus_out_n_6),
        .\sr[4]_i_188_1 (a0bus_out_n_11),
        .\sr[4]_i_188_2 (a0bus_out_n_66),
        .\sr[4]_i_196_0 (a0bus_out_n_31),
        .\sr[4]_i_196_1 (a0bus_out_n_29),
        .\sr[4]_i_196_2 (a0bus_out_n_30),
        .\sr[4]_i_196_3 (a0bus_out_n_35),
        .\sr[4]_i_196_4 (a0bus_out_n_72),
        .\sr[4]_i_196_5 (a0bus_out_n_23),
        .\sr[4]_i_196_6 (a0bus_out_n_21),
        .\sr[4]_i_196_7 (a0bus_out_n_22),
        .\sr[4]_i_196_8 (a0bus_out_n_27),
        .\sr[4]_i_196_9 (a0bus_out_n_70),
        .\sr[4]_i_203_0 (a0bus_out_n_15),
        .\sr[4]_i_203_1 (a0bus_out_n_13),
        .\sr[4]_i_203_2 (a0bus_out_n_14),
        .\sr[4]_i_203_3 (a0bus_out_n_19),
        .\sr[4]_i_203_4 (a0bus_out_n_68),
        .\sr[4]_i_207 (sreg_n_100),
        .\sr[4]_i_207_0 (sreg_n_123),
        .\sr[4]_i_208 (sreg_n_102),
        .\sr[4]_i_208_0 (sreg_n_121),
        .\sr[4]_i_209 (sreg_n_98),
        .\sr[4]_i_209_0 (sreg_n_125),
        .\sr[4]_i_210 (sreg_n_111),
        .\sr[4]_i_210_0 (sreg_n_112),
        .\sr[4]_i_211 (sreg_n_109),
        .\sr[4]_i_211_0 (sreg_n_114),
        .\sr[4]_i_213 (sreg_n_110),
        .\sr[4]_i_213_0 (sreg_n_113),
        .\sr[4]_i_219_0 (\sr[4]_i_219 ),
        .\sr[4]_i_220 (\sr[4]_i_220 ),
        .\sr[4]_i_220_0 (sreg_n_108),
        .\sr[4]_i_220_1 (sreg_n_115),
        .\sr[4]_i_224_0 (sreg_n_106),
        .\sr[4]_i_224_1 (sreg_n_117),
        .\sr[4]_i_225_0 (sreg_n_104),
        .\sr[4]_i_225_1 (sreg_n_119),
        .\sr[4]_i_235 (\sr[4]_i_235 ),
        .\sr[4]_i_235_0 (sreg_n_79),
        .\sr[4]_i_237 (\sr[4]_i_237 ),
        .\sr[4]_i_237_0 (sreg_n_81),
        .\sr[4]_i_240 (\sr[4]_i_240 ),
        .\sr[4]_i_240_0 (sreg_n_90),
        .\sr[4]_i_243 (\sr[4]_i_243 ),
        .\sr[4]_i_243_0 (sreg_n_86),
        .\sr[4]_i_245 (\sr[4]_i_245 ),
        .\sr[4]_i_245_0 (sreg_n_84),
        .\sr[4]_i_30 (\sr[4]_i_30 ),
        .\sr[4]_i_30_0 (bank13_n_130),
        .\sr[4]_i_38 (\sr[4]_i_38 ),
        .\sr[4]_i_44 (\sr[4]_i_44 ),
        .\sr[4]_i_55 (\sr[4]_i_55 ),
        .\sr[4]_i_67 (\sr[4]_i_67 ),
        .\sr[4]_i_77 (a1bus_0[14]),
        .\sr[4]_i_77_0 (a1bus_0[13]),
        .\sr[4]_i_77_1 (a1bus_0[15]),
        .\sr[4]_i_77_2 (a1bus_0[12]),
        .\sr[4]_i_84 (\sr[4]_i_84 ),
        .\sr[4]_i_88 (\tr_reg[1] ),
        .\sr[4]_i_88_0 (\sr_reg[6]_8 ),
        .\sr[4]_i_99 (a1bus_0[7]),
        .\sr[4]_i_99_0 (a1bus_0[8]),
        .\sr[4]_i_99_1 (a1bus_0[9]),
        .\sr[4]_i_99_2 (a1bus_0[10]),
        .\sr[6]_i_11 (a1bus_0[6]),
        .\sr[6]_i_11_0 (a1bus_0[5]),
        .\sr[6]_i_11_1 (\sr[6]_i_11 ),
        .\sr[6]_i_11_2 (\sr[6]_i_11_0 ),
        .\sr[6]_i_11_3 (a1bus_0[0]),
        .\sr[6]_i_11_4 (\sr[6]_i_11_1 ),
        .\sr[6]_i_11_5 (a1bus_0[2]),
        .\sr[6]_i_11_6 (a1bus_0[1]),
        .\sr[6]_i_11_7 ({\sr_reg[15] [6],\sr_reg[15] [1:0]}),
        .\sr[6]_i_11_8 (a1bus_0[3]),
        .\sr[6]_i_11_9 (a1bus_0[4]),
        .\sr[6]_i_15 (\sr[6]_i_15 ),
        .\sr_reg[14] (\sr_reg[14] ),
        .\sr_reg[15] (bank02_n_281),
        .\sr_reg[6] (\sr_reg[6] ),
        .\sr_reg[6]_0 (\sr_reg[6]_0 ),
        .\sr_reg[6]_1 (\sr_reg[6]_1 ),
        .\sr_reg[6]_10 (\sr_reg[6]_12 ),
        .\sr_reg[6]_11 (\sr_reg[6]_13 ),
        .\sr_reg[6]_12 (\sr_reg[6]_14 ),
        .\sr_reg[6]_13 (\sr_reg[6]_15 ),
        .\sr_reg[6]_14 (\sr_reg[6]_17 ),
        .\sr_reg[6]_15 (\sr_reg[6]_20 ),
        .\sr_reg[6]_16 (\sr_reg[6]_21 ),
        .\sr_reg[6]_17 (\sr_reg[6]_22 ),
        .\sr_reg[6]_18 (\sr_reg[6]_23 ),
        .\sr_reg[6]_19 (\sr_reg[6]_24 ),
        .\sr_reg[6]_2 (\sr_reg[6]_2 ),
        .\sr_reg[6]_20 (\sr_reg[6]_28 ),
        .\sr_reg[6]_21 (\sr_reg[6]_30 ),
        .\sr_reg[6]_22 (\sr_reg[6]_31 ),
        .\sr_reg[6]_23 (\sr_reg[6]_32 ),
        .\sr_reg[6]_24 (\sr_reg[6]_34 ),
        .\sr_reg[6]_25 (\sr_reg[6]_36 ),
        .\sr_reg[6]_26 (\sr_reg[6]_37 ),
        .\sr_reg[6]_27 (\sr_reg[6]_38 ),
        .\sr_reg[6]_28 (\sr_reg[6]_42 ),
        .\sr_reg[6]_3 (\sr_reg[6]_3 ),
        .\sr_reg[6]_4 (\sr_reg[6]_4 ),
        .\sr_reg[6]_5 (\sr_reg[6]_5 ),
        .\sr_reg[6]_6 (\sr_reg[6]_7 ),
        .\sr_reg[6]_7 (\sr_reg[6]_9 ),
        .\sr_reg[6]_8 (\sr_reg[6]_10 ),
        .\sr_reg[6]_9 (\sr_reg[6]_11 ),
        .\stat_reg[1] (\stat_reg[1] ),
        .\stat_reg[1]_0 (\stat_reg[1]_0 ),
        .\stat_reg[1]_1 (\stat_reg[1]_1 ),
        .\stat_reg[2] (\stat_reg[2] ),
        .\stat_reg[2]_0 (\stat_reg[2]_0 ),
        .\stat_reg[2]_1 (\stat_reg[2]_1 ),
        .\stat_reg[2]_2 (\stat_reg[2]_2 ),
        .\stat_reg[2]_3 (\stat_reg[2]_3 ),
        .tout__1_carry__0_i_1__0_0(tout__1_carry__0_i_1__0),
        .tout__1_carry__0_i_7__0(tout__1_carry__0_i_7__0),
        .tout__1_carry__0_i_7__0_0(tout__1_carry__0_i_7__0_0),
        .tout__1_carry__0_i_7__0_1(b1bus_out_n_22),
        .tout__1_carry__0_i_7__0_2(b1bus_out_n_11),
        .tout__1_carry__1_i_1__0_0(tout__1_carry__1_i_1__0),
        .tout__1_carry__2(tout__1_carry__2),
        .tout__1_carry__2_0(tout__1_carry__2_0),
        .tout__1_carry__2_1(tout__1_carry__2_1),
        .\tr_reg[10] (\tr_reg[10] ),
        .\tr_reg[10]_0 (\tr_reg[10]_0 ),
        .\tr_reg[11] (\tr_reg[11] ),
        .\tr_reg[11]_0 (\tr_reg[11]_1 ),
        .\tr_reg[12] (\tr_reg[12] ),
        .\tr_reg[12]_0 (\tr_reg[12]_0 ),
        .\tr_reg[12]_1 (\tr_reg[12]_2 ),
        .\tr_reg[13] (\tr_reg[13] ),
        .\tr_reg[13]_0 (\tr_reg[13]_0 ),
        .\tr_reg[14] (\tr_reg[14] ),
        .\tr_reg[14]_0 (\tr_reg[14]_0 ),
        .\tr_reg[14]_1 (\tr_reg[14]_1 ),
        .\tr_reg[15] (\tr_reg[15]_1 ),
        .\tr_reg[5] (\tr_reg[5] ),
        .\tr_reg[5]_0 (\tr_reg[5]_0 ),
        .\tr_reg[6] (\tr_reg[6] ),
        .\tr_reg[6]_0 (\tr_reg[6]_0 ),
        .\tr_reg[7] (\tr_reg[7] ),
        .\tr_reg[7]_0 (\tr_reg[7]_0 ),
        .\tr_reg[8] (\tr_reg[8] ),
        .\tr_reg[8]_0 (\tr_reg[8]_0 ),
        .\tr_reg[9] (\tr_reg[9] ),
        .\tr_reg[9]_0 (\tr_reg[9]_0 ));
  mcss_rgf_bank_5 bank13
       (.SR(SR),
        .a0bus_sel_0(a0bus_sel_0),
        .a1bus_b13(a1bus_b13),
        .a1bus_sel_0({a1bus_sel_0[3:2],a1bus_sel_0[0]}),
        .b0bus_sel_0(b0bus_sel_0),
        .\badr[0]_INST_0_i_1 (sreg_n_128),
        .\badr[0]_INST_0_i_1_0 (sreg_n_144),
        .\badr[10]_INST_0_i_1 (sreg_n_138),
        .\badr[10]_INST_0_i_1_0 (sreg_n_154),
        .\badr[11]_INST_0_i_1 (sreg_n_139),
        .\badr[11]_INST_0_i_1_0 (sreg_n_155),
        .\badr[12]_INST_0_i_1 (sreg_n_140),
        .\badr[12]_INST_0_i_1_0 (sreg_n_156),
        .\badr[13]_INST_0_i_1 (sreg_n_141),
        .\badr[13]_INST_0_i_1_0 (sreg_n_157),
        .\badr[14]_INST_0_i_1 (sreg_n_142),
        .\badr[14]_INST_0_i_1_0 (sreg_n_158),
        .\badr[15]_INST_0_i_1 (\badr[15]_INST_0_i_1_1 ),
        .\badr[15]_INST_0_i_1_0 (sreg_n_143),
        .\badr[15]_INST_0_i_1_1 (sreg_n_159),
        .\badr[15]_INST_0_i_2 (\badr[15]_INST_0_i_2 ),
        .\badr[1]_INST_0_i_1 (sreg_n_129),
        .\badr[1]_INST_0_i_1_0 (sreg_n_145),
        .\badr[2]_INST_0_i_1 (sreg_n_130),
        .\badr[2]_INST_0_i_1_0 (sreg_n_146),
        .\badr[3]_INST_0_i_1 (sreg_n_131),
        .\badr[3]_INST_0_i_1_0 (sreg_n_147),
        .\badr[4]_INST_0_i_1 (sreg_n_132),
        .\badr[4]_INST_0_i_1_0 (sreg_n_148),
        .\badr[5]_INST_0_i_1 (sreg_n_133),
        .\badr[5]_INST_0_i_1_0 (sreg_n_149),
        .\badr[6]_INST_0_i_1 (sreg_n_134),
        .\badr[6]_INST_0_i_1_0 (sreg_n_150),
        .\badr[7]_INST_0_i_1 (sreg_n_135),
        .\badr[7]_INST_0_i_1_0 (sreg_n_151),
        .\badr[8]_INST_0_i_1 (sreg_n_136),
        .\badr[8]_INST_0_i_1_0 (sreg_n_152),
        .\badr[9]_INST_0_i_1 (sreg_n_137),
        .\badr[9]_INST_0_i_1_0 (sreg_n_153),
        .\bbus_o[0]_INST_0_i_7 (\bbus_o[0]_INST_0_i_7 ),
        .\bbus_o[0]_INST_0_i_7_0 (\bbus_o[0]_INST_0_i_7_0 ),
        .\bbus_o[0]_INST_0_i_7_1 (\bbus_o[0]_INST_0_i_7_1 ),
        .\bbus_o[0]_INST_0_i_7_2 (\bbus_o[0]_INST_0_i_7_2 ),
        .\bbus_o[0]_INST_0_i_7_3 (\bbus_o[0]_INST_0_i_7_3 ),
        .\bbus_o[0]_INST_0_i_7_4 (\bbus_o[0]_INST_0_i_7_4 ),
        .\bbus_o[0]_INST_0_i_7_5 (\bbus_o[0]_INST_0_i_7_5 ),
        .\bbus_o[0]_INST_0_i_7_6 (\bbus_o[0]_INST_0_i_7_6 ),
        .\bbus_o[1]_INST_0_i_7 (\bbus_o[1]_INST_0_i_7 ),
        .\bbus_o[1]_INST_0_i_7_0 (\bbus_o[1]_INST_0_i_7_0 ),
        .\bbus_o[1]_INST_0_i_7_1 (\bbus_o[1]_INST_0_i_7_1 ),
        .\bbus_o[1]_INST_0_i_7_2 (\bbus_o[1]_INST_0_i_7_2 ),
        .\bbus_o[1]_INST_0_i_7_3 (\bbus_o[1]_INST_0_i_7_3 ),
        .\bbus_o[1]_INST_0_i_7_4 (\bbus_o[1]_INST_0_i_7_4 ),
        .\bbus_o[1]_INST_0_i_7_5 (\bbus_o[1]_INST_0_i_7_5 ),
        .\bbus_o[1]_INST_0_i_7_6 (\bbus_o[1]_INST_0_i_7_6 ),
        .\bbus_o[2]_INST_0_i_7 (\bbus_o[2]_INST_0_i_7 ),
        .\bbus_o[2]_INST_0_i_7_0 (\bbus_o[2]_INST_0_i_7_0 ),
        .\bbus_o[2]_INST_0_i_7_1 (\bbus_o[2]_INST_0_i_7_1 ),
        .\bbus_o[2]_INST_0_i_7_2 (\bbus_o[2]_INST_0_i_7_2 ),
        .\bbus_o[2]_INST_0_i_7_3 (\bbus_o[2]_INST_0_i_7_3 ),
        .\bbus_o[2]_INST_0_i_7_4 (\bbus_o[2]_INST_0_i_7_4 ),
        .\bbus_o[2]_INST_0_i_7_5 (\bbus_o[2]_INST_0_i_7_5 ),
        .\bbus_o[2]_INST_0_i_7_6 (\bbus_o[2]_INST_0_i_7_6 ),
        .\bbus_o[3]_INST_0_i_7 (\bbus_o[3]_INST_0_i_7 ),
        .\bbus_o[3]_INST_0_i_7_0 (\bbus_o[3]_INST_0_i_7_0 ),
        .\bbus_o[3]_INST_0_i_7_1 (\bbus_o[3]_INST_0_i_7_1 ),
        .\bbus_o[3]_INST_0_i_7_2 (\bbus_o[3]_INST_0_i_7_2 ),
        .\bbus_o[3]_INST_0_i_7_3 (\bbus_o[3]_INST_0_i_7_3 ),
        .\bbus_o[3]_INST_0_i_7_4 (\bbus_o[3]_INST_0_i_7_4 ),
        .\bbus_o[3]_INST_0_i_7_5 (\bbus_o[3]_INST_0_i_7_5 ),
        .\bbus_o[3]_INST_0_i_7_6 (\bbus_o[3]_INST_0_i_7_6 ),
        .\bbus_o[4]_INST_0_i_7 (\bbus_o[4]_INST_0_i_7 ),
        .\bbus_o[4]_INST_0_i_7_0 (\bbus_o[4]_INST_0_i_7_0 ),
        .\bbus_o[4]_INST_0_i_7_1 (\bbus_o[4]_INST_0_i_7_1 ),
        .\bbus_o[4]_INST_0_i_7_2 (\bbus_o[4]_INST_0_i_7_2 ),
        .\bbus_o[4]_INST_0_i_7_3 (\bbus_o[4]_INST_0_i_7_3 ),
        .\bbus_o[4]_INST_0_i_7_4 (\bbus_o[4]_INST_0_i_7_4 ),
        .\bbus_o[4]_INST_0_i_7_5 (\bbus_o[4]_INST_0_i_7_5 ),
        .\bbus_o[4]_INST_0_i_7_6 (\bbus_o[4]_INST_0_i_7_6 ),
        .\bdatw[10]_INST_0_i_43 (\bdatw[10]_INST_0_i_43 ),
        .\bdatw[10]_INST_0_i_43_0 (\bdatw[10]_INST_0_i_43_0 ),
        .\bdatw[11]_INST_0_i_44 (\bdatw[11]_INST_0_i_44 ),
        .\bdatw[11]_INST_0_i_44_0 (\bdatw[11]_INST_0_i_44_0 ),
        .\bdatw[12]_INST_0_i_42 (\bdatw[12]_INST_0_i_42 ),
        .\bdatw[12]_INST_0_i_42_0 (\bdatw[12]_INST_0_i_42_0 ),
        .\bdatw[8]_INST_0_i_43 (\bdatw[8]_INST_0_i_43 ),
        .\bdatw[8]_INST_0_i_43_0 (\bdatw[8]_INST_0_i_43_0 ),
        .\bdatw[9]_INST_0_i_42 (\bdatw[9]_INST_0_i_42 ),
        .\bdatw[9]_INST_0_i_42_0 (\bdatw[9]_INST_0_i_42_0 ),
        .clk(clk),
        .ctl_sela0(ctl_sela0),
        .ctl_sela0_rn(ctl_sela0_rn),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .fdat(fdat),
        .\fdat[15] (\fdat[15] ),
        .fdat_12_sp_1(fdat_12_sn_1),
        .fdatx(fdatx),
        .\fdatx[15] (\fdatx[15] ),
        .gr6_bus1(\a1buso/gr6_bus1 ),
        .gr6_bus1_0(\a1buso2l/gr6_bus1_0 ),
        .\grn_reg[0] (bank13_n_183),
        .\grn_reg[0]_0 (bank13_n_199),
        .\grn_reg[0]_1 (bank13_n_215),
        .\grn_reg[0]_10 (bank13_n_350),
        .\grn_reg[0]_11 (bank13_n_366),
        .\grn_reg[0]_12 (bank13_n_382),
        .\grn_reg[0]_13 (bank13_n_399),
        .\grn_reg[0]_14 (bank13_n_415),
        .\grn_reg[0]_15 (bank13_n_431),
        .\grn_reg[0]_16 (bank13_n_446),
        .\grn_reg[0]_2 (bank13_n_231),
        .\grn_reg[0]_3 (bank13_n_247),
        .\grn_reg[0]_4 (bank13_n_265),
        .\grn_reg[0]_5 (bank13_n_266),
        .\grn_reg[0]_6 (bank13_n_282),
        .\grn_reg[0]_7 (bank13_n_297),
        .\grn_reg[0]_8 (bank13_n_302),
        .\grn_reg[0]_9 (bank13_n_334),
        .\grn_reg[10] (bank13_n_173),
        .\grn_reg[10]_0 (bank13_n_189),
        .\grn_reg[10]_1 (bank13_n_205),
        .\grn_reg[10]_10 (bank13_n_372),
        .\grn_reg[10]_11 (bank13_n_389),
        .\grn_reg[10]_12 (bank13_n_405),
        .\grn_reg[10]_13 (bank13_n_421),
        .\grn_reg[10]_14 (bank13_n_436),
        .\grn_reg[10]_2 (bank13_n_221),
        .\grn_reg[10]_3 (bank13_n_237),
        .\grn_reg[10]_4 (bank13_n_255),
        .\grn_reg[10]_5 (bank13_n_272),
        .\grn_reg[10]_6 (bank13_n_287),
        .\grn_reg[10]_7 (bank13_n_324),
        .\grn_reg[10]_8 (bank13_n_340),
        .\grn_reg[10]_9 (bank13_n_356),
        .\grn_reg[11] (bank13_n_172),
        .\grn_reg[11]_0 (bank13_n_188),
        .\grn_reg[11]_1 (bank13_n_204),
        .\grn_reg[11]_10 (bank13_n_371),
        .\grn_reg[11]_11 (bank13_n_388),
        .\grn_reg[11]_12 (bank13_n_404),
        .\grn_reg[11]_13 (bank13_n_420),
        .\grn_reg[11]_14 (bank13_n_435),
        .\grn_reg[11]_2 (bank13_n_220),
        .\grn_reg[11]_3 (bank13_n_236),
        .\grn_reg[11]_4 (bank13_n_254),
        .\grn_reg[11]_5 (bank13_n_271),
        .\grn_reg[11]_6 (bank13_n_286),
        .\grn_reg[11]_7 (bank13_n_323),
        .\grn_reg[11]_8 (bank13_n_339),
        .\grn_reg[11]_9 (bank13_n_355),
        .\grn_reg[12] (bank13_n_171),
        .\grn_reg[12]_0 (bank13_n_187),
        .\grn_reg[12]_1 (bank13_n_203),
        .\grn_reg[12]_10 (bank13_n_370),
        .\grn_reg[12]_11 (bank13_n_387),
        .\grn_reg[12]_12 (bank13_n_403),
        .\grn_reg[12]_13 (bank13_n_419),
        .\grn_reg[12]_14 (bank13_n_434),
        .\grn_reg[12]_2 (bank13_n_219),
        .\grn_reg[12]_3 (bank13_n_235),
        .\grn_reg[12]_4 (bank13_n_253),
        .\grn_reg[12]_5 (bank13_n_270),
        .\grn_reg[12]_6 (bank13_n_285),
        .\grn_reg[12]_7 (bank13_n_322),
        .\grn_reg[12]_8 (bank13_n_338),
        .\grn_reg[12]_9 (bank13_n_354),
        .\grn_reg[13] (bank13_n_170),
        .\grn_reg[13]_0 (bank13_n_186),
        .\grn_reg[13]_1 (bank13_n_202),
        .\grn_reg[13]_10 (bank13_n_369),
        .\grn_reg[13]_11 (bank13_n_386),
        .\grn_reg[13]_12 (bank13_n_402),
        .\grn_reg[13]_13 (bank13_n_418),
        .\grn_reg[13]_14 (bank13_n_433),
        .\grn_reg[13]_2 (bank13_n_218),
        .\grn_reg[13]_3 (bank13_n_234),
        .\grn_reg[13]_4 (bank13_n_252),
        .\grn_reg[13]_5 (bank13_n_269),
        .\grn_reg[13]_6 (bank13_n_284),
        .\grn_reg[13]_7 (bank13_n_321),
        .\grn_reg[13]_8 (bank13_n_337),
        .\grn_reg[13]_9 (bank13_n_353),
        .\grn_reg[14] (bank13_n_169),
        .\grn_reg[14]_0 (bank13_n_185),
        .\grn_reg[14]_1 (bank13_n_201),
        .\grn_reg[14]_10 (bank13_n_368),
        .\grn_reg[14]_11 (bank13_n_385),
        .\grn_reg[14]_12 (bank13_n_401),
        .\grn_reg[14]_13 (bank13_n_417),
        .\grn_reg[14]_14 (bank13_n_432),
        .\grn_reg[14]_2 (bank13_n_217),
        .\grn_reg[14]_3 (bank13_n_233),
        .\grn_reg[14]_4 (bank13_n_251),
        .\grn_reg[14]_5 (bank13_n_268),
        .\grn_reg[14]_6 (bank13_n_283),
        .\grn_reg[14]_7 (bank13_n_320),
        .\grn_reg[14]_8 (bank13_n_336),
        .\grn_reg[14]_9 (bank13_n_352),
        .\grn_reg[15] ({bank13_n_26,bank13_n_27,bank13_n_28,bank13_n_29,bank13_n_30,bank13_n_31,bank13_n_32,bank13_n_33,bank13_n_34,bank13_n_35,bank13_n_36,\grn_reg[4]_1 }),
        .\grn_reg[15]_0 ({bank13_n_42,bank13_n_43,bank13_n_44,bank13_n_45,bank13_n_46,bank13_n_47,bank13_n_48,bank13_n_49,bank13_n_50,bank13_n_51,bank13_n_52,\grn_reg[4]_2 }),
        .\grn_reg[15]_1 (\grn_reg[15]_0 ),
        .\grn_reg[15]_10 (bank13_n_250),
        .\grn_reg[15]_11 (bank13_n_267),
        .\grn_reg[15]_12 (bank13_n_319),
        .\grn_reg[15]_13 (bank13_n_335),
        .\grn_reg[15]_14 (bank13_n_351),
        .\grn_reg[15]_15 (bank13_n_367),
        .\grn_reg[15]_16 (bank13_n_383),
        .\grn_reg[15]_17 (bank13_n_400),
        .\grn_reg[15]_18 (bank13_n_416),
        .\grn_reg[15]_19 (\grn_reg[15]_34 ),
        .\grn_reg[15]_2 ({bank13_n_89,bank13_n_90,bank13_n_91,bank13_n_92,bank13_n_93,bank13_n_94,bank13_n_95,bank13_n_96,bank13_n_97,bank13_n_98,bank13_n_99,\grn_reg[4]_6 }),
        .\grn_reg[15]_20 (\grn_reg[15]_35 ),
        .\grn_reg[15]_21 (\grn_reg[15]_36 ),
        .\grn_reg[15]_22 (\grn_reg[15]_37 ),
        .\grn_reg[15]_23 (\grn_reg[15]_38 ),
        .\grn_reg[15]_24 (\grn_reg[15]_39 ),
        .\grn_reg[15]_25 (\grn_reg[15]_40 ),
        .\grn_reg[15]_26 (\grn_reg[15]_41 ),
        .\grn_reg[15]_27 (\grn_reg[15]_42 ),
        .\grn_reg[15]_28 (\grn_reg[15]_43 ),
        .\grn_reg[15]_29 (\grn_reg[15]_44 ),
        .\grn_reg[15]_3 ({bank13_n_105,bank13_n_106,bank13_n_107,bank13_n_108,bank13_n_109,bank13_n_110,bank13_n_111,bank13_n_112,bank13_n_113,bank13_n_114,bank13_n_115,bank13_n_116,bank13_n_117,bank13_n_118,bank13_n_119,bank13_n_120}),
        .\grn_reg[15]_30 (\grn_reg[15]_45 ),
        .\grn_reg[15]_31 (\grn_reg[15]_46 ),
        .\grn_reg[15]_32 (\grn_reg[15]_47 ),
        .\grn_reg[15]_33 (\grn_reg[15]_48 ),
        .\grn_reg[15]_34 (\grn_reg[15]_49 ),
        .\grn_reg[15]_35 (\grn_reg[15]_50 ),
        .\grn_reg[15]_36 (\grn_reg[15]_51 ),
        .\grn_reg[15]_37 (\grn_reg[15]_52 ),
        .\grn_reg[15]_38 (\grn_reg[15]_53 ),
        .\grn_reg[15]_39 (\grn_reg[15]_54 ),
        .\grn_reg[15]_4 (bank13_n_168),
        .\grn_reg[15]_40 (\grn_reg[15]_55 ),
        .\grn_reg[15]_41 (\grn_reg[15]_56 ),
        .\grn_reg[15]_42 (\grn_reg[15]_57 ),
        .\grn_reg[15]_43 (\grn_reg[15]_58 ),
        .\grn_reg[15]_44 (\grn_reg[15]_59 ),
        .\grn_reg[15]_45 (\grn_reg[15]_60 ),
        .\grn_reg[15]_46 (\grn_reg[15]_61 ),
        .\grn_reg[15]_47 (\grn_reg[15]_62 ),
        .\grn_reg[15]_48 (\grn_reg[15]_63 ),
        .\grn_reg[15]_49 (\grn_reg[15]_64 ),
        .\grn_reg[15]_5 (bank13_n_184),
        .\grn_reg[15]_50 (\grn_reg[15]_65 ),
        .\grn_reg[15]_6 (bank13_n_200),
        .\grn_reg[15]_7 (bank13_n_216),
        .\grn_reg[15]_8 (bank13_n_232),
        .\grn_reg[15]_9 (bank13_n_248),
        .\grn_reg[1] (bank13_n_182),
        .\grn_reg[1]_0 (bank13_n_198),
        .\grn_reg[1]_1 (bank13_n_214),
        .\grn_reg[1]_10 (bank13_n_365),
        .\grn_reg[1]_11 (bank13_n_381),
        .\grn_reg[1]_12 (bank13_n_398),
        .\grn_reg[1]_13 (bank13_n_414),
        .\grn_reg[1]_14 (bank13_n_430),
        .\grn_reg[1]_15 (bank13_n_445),
        .\grn_reg[1]_2 (bank13_n_230),
        .\grn_reg[1]_3 (bank13_n_246),
        .\grn_reg[1]_4 (bank13_n_264),
        .\grn_reg[1]_5 (bank13_n_281),
        .\grn_reg[1]_6 (bank13_n_296),
        .\grn_reg[1]_7 (bank13_n_301),
        .\grn_reg[1]_8 (bank13_n_333),
        .\grn_reg[1]_9 (bank13_n_349),
        .\grn_reg[2] (bank13_n_181),
        .\grn_reg[2]_0 (bank13_n_197),
        .\grn_reg[2]_1 (bank13_n_213),
        .\grn_reg[2]_10 (bank13_n_364),
        .\grn_reg[2]_11 (bank13_n_380),
        .\grn_reg[2]_12 (bank13_n_397),
        .\grn_reg[2]_13 (bank13_n_413),
        .\grn_reg[2]_14 (bank13_n_429),
        .\grn_reg[2]_15 (bank13_n_444),
        .\grn_reg[2]_2 (bank13_n_229),
        .\grn_reg[2]_3 (bank13_n_245),
        .\grn_reg[2]_4 (bank13_n_263),
        .\grn_reg[2]_5 (bank13_n_280),
        .\grn_reg[2]_6 (bank13_n_295),
        .\grn_reg[2]_7 (bank13_n_300),
        .\grn_reg[2]_8 (bank13_n_332),
        .\grn_reg[2]_9 (bank13_n_348),
        .\grn_reg[3] (bank13_n_180),
        .\grn_reg[3]_0 (bank13_n_196),
        .\grn_reg[3]_1 (bank13_n_212),
        .\grn_reg[3]_10 (bank13_n_363),
        .\grn_reg[3]_11 (bank13_n_379),
        .\grn_reg[3]_12 (bank13_n_396),
        .\grn_reg[3]_13 (bank13_n_412),
        .\grn_reg[3]_14 (bank13_n_428),
        .\grn_reg[3]_15 (bank13_n_443),
        .\grn_reg[3]_2 (bank13_n_228),
        .\grn_reg[3]_3 (bank13_n_244),
        .\grn_reg[3]_4 (bank13_n_262),
        .\grn_reg[3]_5 (bank13_n_279),
        .\grn_reg[3]_6 (bank13_n_294),
        .\grn_reg[3]_7 (bank13_n_299),
        .\grn_reg[3]_8 (bank13_n_331),
        .\grn_reg[3]_9 (bank13_n_347),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (\grn_reg[4]_0 ),
        .\grn_reg[4]_1 (\grn_reg[4]_3 ),
        .\grn_reg[4]_10 (bank13_n_261),
        .\grn_reg[4]_11 (bank13_n_278),
        .\grn_reg[4]_12 (bank13_n_293),
        .\grn_reg[4]_13 (bank13_n_298),
        .\grn_reg[4]_14 (bank13_n_330),
        .\grn_reg[4]_15 (bank13_n_346),
        .\grn_reg[4]_16 (bank13_n_362),
        .\grn_reg[4]_17 (bank13_n_378),
        .\grn_reg[4]_18 (bank13_n_395),
        .\grn_reg[4]_19 (bank13_n_411),
        .\grn_reg[4]_2 (\grn_reg[4]_4 ),
        .\grn_reg[4]_20 (bank13_n_427),
        .\grn_reg[4]_21 (bank13_n_442),
        .\grn_reg[4]_3 (\grn_reg[4]_5 ),
        .\grn_reg[4]_4 (\grn_reg[4]_7 ),
        .\grn_reg[4]_5 (bank13_n_179),
        .\grn_reg[4]_6 (bank13_n_195),
        .\grn_reg[4]_7 (bank13_n_211),
        .\grn_reg[4]_8 (bank13_n_227),
        .\grn_reg[4]_9 (bank13_n_243),
        .\grn_reg[5] (bank13_n_178),
        .\grn_reg[5]_0 (bank13_n_194),
        .\grn_reg[5]_1 (bank13_n_210),
        .\grn_reg[5]_10 (bank13_n_377),
        .\grn_reg[5]_11 (bank13_n_394),
        .\grn_reg[5]_12 (bank13_n_410),
        .\grn_reg[5]_13 (bank13_n_426),
        .\grn_reg[5]_14 (bank13_n_441),
        .\grn_reg[5]_2 (bank13_n_226),
        .\grn_reg[5]_3 (bank13_n_242),
        .\grn_reg[5]_4 (bank13_n_260),
        .\grn_reg[5]_5 (bank13_n_277),
        .\grn_reg[5]_6 (bank13_n_292),
        .\grn_reg[5]_7 (bank13_n_329),
        .\grn_reg[5]_8 (bank13_n_345),
        .\grn_reg[5]_9 (bank13_n_361),
        .\grn_reg[6] (bank13_n_177),
        .\grn_reg[6]_0 (bank13_n_193),
        .\grn_reg[6]_1 (bank13_n_209),
        .\grn_reg[6]_10 (bank13_n_376),
        .\grn_reg[6]_11 (bank13_n_393),
        .\grn_reg[6]_12 (bank13_n_409),
        .\grn_reg[6]_13 (bank13_n_425),
        .\grn_reg[6]_14 (bank13_n_440),
        .\grn_reg[6]_2 (bank13_n_225),
        .\grn_reg[6]_3 (bank13_n_241),
        .\grn_reg[6]_4 (bank13_n_259),
        .\grn_reg[6]_5 (bank13_n_276),
        .\grn_reg[6]_6 (bank13_n_291),
        .\grn_reg[6]_7 (bank13_n_328),
        .\grn_reg[6]_8 (bank13_n_344),
        .\grn_reg[6]_9 (bank13_n_360),
        .\grn_reg[7] (bank13_n_176),
        .\grn_reg[7]_0 (bank13_n_192),
        .\grn_reg[7]_1 (bank13_n_208),
        .\grn_reg[7]_10 (bank13_n_375),
        .\grn_reg[7]_11 (bank13_n_392),
        .\grn_reg[7]_12 (bank13_n_408),
        .\grn_reg[7]_13 (bank13_n_424),
        .\grn_reg[7]_14 (bank13_n_439),
        .\grn_reg[7]_2 (bank13_n_224),
        .\grn_reg[7]_3 (bank13_n_240),
        .\grn_reg[7]_4 (bank13_n_258),
        .\grn_reg[7]_5 (bank13_n_275),
        .\grn_reg[7]_6 (bank13_n_290),
        .\grn_reg[7]_7 (bank13_n_327),
        .\grn_reg[7]_8 (bank13_n_343),
        .\grn_reg[7]_9 (bank13_n_359),
        .\grn_reg[8] (bank13_n_175),
        .\grn_reg[8]_0 (bank13_n_191),
        .\grn_reg[8]_1 (bank13_n_207),
        .\grn_reg[8]_10 (bank13_n_374),
        .\grn_reg[8]_11 (bank13_n_391),
        .\grn_reg[8]_12 (bank13_n_407),
        .\grn_reg[8]_13 (bank13_n_423),
        .\grn_reg[8]_14 (bank13_n_438),
        .\grn_reg[8]_2 (bank13_n_223),
        .\grn_reg[8]_3 (bank13_n_239),
        .\grn_reg[8]_4 (bank13_n_257),
        .\grn_reg[8]_5 (bank13_n_274),
        .\grn_reg[8]_6 (bank13_n_289),
        .\grn_reg[8]_7 (bank13_n_326),
        .\grn_reg[8]_8 (bank13_n_342),
        .\grn_reg[8]_9 (bank13_n_358),
        .\grn_reg[9] (bank13_n_174),
        .\grn_reg[9]_0 (bank13_n_190),
        .\grn_reg[9]_1 (bank13_n_206),
        .\grn_reg[9]_10 (bank13_n_373),
        .\grn_reg[9]_11 (bank13_n_390),
        .\grn_reg[9]_12 (bank13_n_406),
        .\grn_reg[9]_13 (bank13_n_422),
        .\grn_reg[9]_14 (bank13_n_437),
        .\grn_reg[9]_2 (bank13_n_222),
        .\grn_reg[9]_3 (bank13_n_238),
        .\grn_reg[9]_4 (bank13_n_256),
        .\grn_reg[9]_5 (bank13_n_273),
        .\grn_reg[9]_6 (bank13_n_288),
        .\grn_reg[9]_7 (bank13_n_325),
        .\grn_reg[9]_8 (bank13_n_341),
        .\grn_reg[9]_9 (bank13_n_357),
        .\i_/badr[0]_INST_0_i_18 (\i_/badr[15]_INST_0_i_19 ),
        .\i_/badr[0]_INST_0_i_18_0 (\i_/badr[15]_INST_0_i_19_0 ),
        .\i_/badr[0]_INST_0_i_18_1 (\i_/badr[15]_INST_0_i_19_1 ),
        .\i_/badr[15]_INST_0_i_135 (\sr_reg[0]_0 ),
        .\i_/badr[15]_INST_0_i_135_0 (\i_/badr[15]_INST_0_i_43 ),
        .\i_/badr[15]_INST_0_i_135_1 (\i_/badr[15]_INST_0_i_43_0 ),
        .\i_/badr[15]_INST_0_i_52 (\sr_reg[0]_1 ),
        .\i_/bbus_o[4]_INST_0_i_20 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .\i_/bbus_o[4]_INST_0_i_20_0 (\i_/bbus_o[4]_INST_0_i_20 ),
        .\i_/bbus_o[4]_INST_0_i_20_1 (\i_/bbus_o[4]_INST_0_i_20_0 ),
        .\i_/bbus_o[4]_INST_0_i_21 (\i_/bdatw[15]_INST_0_i_9_1 ),
        .\i_/bbus_o[4]_INST_0_i_21_0 (\i_/bdatw[15]_INST_0_i_9_2 ),
        .\i_/bbus_o[4]_INST_0_i_21_1 (\i_/bdatw[15]_INST_0_i_24 ),
        .\i_/bdatw[15]_INST_0_i_121 (\i_/bdatw[15]_INST_0_i_112 ),
        .\i_/bdatw[15]_INST_0_i_121_0 (\i_/bdatw[15]_INST_0_i_112_0 ),
        .\i_/bdatw[15]_INST_0_i_121_1 (\i_/bdatw[15]_INST_0_i_112_1 ),
        .\i_/bdatw[15]_INST_0_i_124 (\i_/bdatw[15]_INST_0_i_44 ),
        .\i_/bdatw[15]_INST_0_i_212 (\i_/bdatw[15]_INST_0_i_113 ),
        .\i_/bdatw[15]_INST_0_i_33 (\i_/bdatw[15]_INST_0_i_77 ),
        .\i_/bdatw[15]_INST_0_i_34 (\i_/bdatw[15]_INST_0_i_9_3 ),
        .\i_/bdatw[15]_INST_0_i_34_0 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_92 (\i_/bdatw[15]_INST_0_i_24_0 ),
        .\ir0_id_fl[20]_i_4 (\ir0_id_fl[20]_i_4 ),
        .\nir_id_reg[20] (\nir_id_reg[20] ),
        .out(\grn_reg[15] ),
        .p_0_in(p_0_in_1),
        .\rgf_c0bus_wb[12]_i_7 (bank02_n_281),
        .\rgf_c0bus_wb[13]_i_13 (\sr_reg[6]_33 ),
        .\rgf_c0bus_wb[13]_i_27_0 (\rgf_c0bus_wb[13]_i_27 ),
        .\rgf_c0bus_wb[13]_i_30_0 (\rgf_c0bus_wb[13]_i_30 ),
        .\rgf_c0bus_wb[15]_i_23_0 (a0bus_out_n_46),
        .\rgf_c0bus_wb[15]_i_23_1 (a0bus_out_n_45),
        .\rgf_c0bus_wb[15]_i_23_2 (a0bus_out_n_76),
        .\rgf_c0bus_wb[15]_i_23_3 (a0bus_out_n_74),
        .\rgf_c0bus_wb[15]_i_23_4 (a0bus_out_n_54),
        .\rgf_c0bus_wb[15]_i_23_5 (a0bus_out_n_53),
        .\rgf_c0bus_wb[15]_i_23_6 (a0bus_out_n_78),
        .\rgf_c0bus_wb[15]_i_23_7 (a0bus_out_n_3),
        .\rgf_c0bus_wb[15]_i_23_8 (a0bus_out_n_2),
        .\rgf_c0bus_wb[15]_i_23_9 (a0bus_out_n_1),
        .\rgf_c0bus_wb[4]_i_12 (a0bus_out_n_7),
        .\rgf_c0bus_wb[4]_i_12_0 (a0bus_out_n_6),
        .\rgf_c0bus_wb[4]_i_12_1 (a0bus_out_n_5),
        .\rgf_c0bus_wb[4]_i_12_2 (a0bus_out_n_64),
        .\rgf_c0bus_wb[4]_i_26_0 (\rgf_c0bus_wb[4]_i_26 ),
        .\rgf_c0bus_wb[4]_i_29_0 (\rgf_c0bus_wb[4]_i_29 ),
        .\rgf_c0bus_wb[4]_i_31_0 (\rgf_c0bus_wb[4]_i_31 ),
        .\rgf_c0bus_wb[4]_i_32_0 (\rgf_c0bus_wb[4]_i_32 ),
        .\rgf_c0bus_wb[4]_i_33_0 (\rgf_c0bus_wb[4]_i_33 ),
        .\rgf_c0bus_wb[4]_i_8_0 (a0bus_out_n_71),
        .\rgf_c0bus_wb[4]_i_8_1 (a0bus_out_n_31),
        .\rgf_c0bus_wb[4]_i_8_2 (a0bus_out_n_18),
        .\rgf_c0bus_wb[4]_i_8_3 (a0bus_out_n_17),
        .\rgf_c0bus_wb[4]_i_8_4 (a0bus_out_n_19),
        .\rgf_c0bus_wb[4]_i_8_5 (a0bus_out_n_26),
        .\rgf_c0bus_wb[4]_i_8_6 (a0bus_out_n_25),
        .\rgf_c0bus_wb[4]_i_8_7 (a0bus_out_n_27),
        .\rgf_c0bus_wb[4]_i_8_8 (a0bus_out_n_69),
        .\rgf_c0bus_wb[4]_i_8_9 (a0bus_out_n_23),
        .\rgf_c1bus_wb[14]_i_28 (\rgf_c1bus_wb[14]_i_28_3 ),
        .\rgf_c1bus_wb[4]_i_11 ({a1bus_b02[14:8],a1bus_b02[6],a1bus_b02[4:0]}),
        .\rgf_c1bus_wb[4]_i_11_0 (a1bus_out_n_52),
        .\rgf_c1bus_wb[4]_i_11_1 (a1bus_out_n_53),
        .\rgf_c1bus_wb[4]_i_11_2 (a1bus_out_n_5),
        .\rgf_c1bus_wb[4]_i_11_3 (a1bus_out_n_49),
        .\rgf_c1bus_wb[4]_i_11_4 (a1bus_out_n_3),
        .\rgf_c1bus_wb[4]_i_11_5 (a1bus_out_n_11),
        .\rgf_c1bus_wb[4]_i_11_6 (a1bus_out_n_9),
        .\rgf_c1bus_wb[4]_i_28_0 (\rgf_c1bus_wb[4]_i_28 ),
        .\rgf_c1bus_wb[4]_i_32 (\rgf_c1bus_wb[4]_i_32 ),
        .\rgf_c1bus_wb[4]_i_32_0 (sreg_n_71),
        .\rgf_c1bus_wb[4]_i_32_1 (\rgf_c1bus_wb[4]_i_32_0 ),
        .\rgf_c1bus_wb[4]_i_32_2 (sreg_n_50),
        .\rgf_c1bus_wb[4]_i_34 (\rgf_c1bus_wb[4]_i_34 ),
        .\rgf_c1bus_wb[4]_i_34_0 (sreg_n_72),
        .\rgf_c1bus_wb[4]_i_34_1 (\rgf_c1bus_wb[4]_i_34_0 ),
        .\rgf_c1bus_wb[4]_i_34_2 (sreg_n_51),
        .\rgf_c1bus_wb[4]_i_36 (\rgf_c1bus_wb[4]_i_36 ),
        .\rgf_c1bus_wb[4]_i_36_0 (sreg_n_73),
        .\rgf_c1bus_wb[4]_i_36_1 (\rgf_c1bus_wb[4]_i_36_0 ),
        .\rgf_c1bus_wb[4]_i_36_2 (sreg_n_52),
        .\rgf_c1bus_wb[4]_i_38 (\rgf_c1bus_wb[4]_i_38 ),
        .\rgf_c1bus_wb[4]_i_38_0 (sreg_n_74),
        .\rgf_c1bus_wb[4]_i_38_1 (\rgf_c1bus_wb[4]_i_38_0 ),
        .\rgf_c1bus_wb[4]_i_38_2 (sreg_n_53),
        .\rgf_c1bus_wb[4]_i_40 (\rgf_c1bus_wb[4]_i_40 ),
        .\rgf_c1bus_wb[4]_i_40_0 (sreg_n_60),
        .\rgf_c1bus_wb[4]_i_42 (\rgf_c1bus_wb[4]_i_42 ),
        .\rgf_c1bus_wb[4]_i_42_0 (sreg_n_61),
        .\rgf_c1bus_wb[4]_i_42_1 (\rgf_c1bus_wb[4]_i_42_0 ),
        .\rgf_c1bus_wb[4]_i_42_2 (sreg_n_40),
        .\rgf_c1bus_wb[4]_i_44 (\rgf_c1bus_wb[4]_i_44 ),
        .\rgf_c1bus_wb[4]_i_44_0 (sreg_n_54),
        .\rgf_c1bus_wb[4]_i_45 (\rgf_c1bus_wb[4]_i_45 ),
        .\rgf_c1bus_wb[4]_i_45_0 (sreg_n_39),
        .\rgf_c1bus_wb[4]_i_48 (\rgf_c1bus_wb[4]_i_48 ),
        .\rgf_c1bus_wb[4]_i_48_0 (sreg_n_63),
        .\rgf_c1bus_wb[4]_i_48_1 (\rgf_c1bus_wb[4]_i_48_0 ),
        .\rgf_c1bus_wb[4]_i_48_2 (sreg_n_42),
        .\rgf_c1bus_wb[4]_i_50 (\rgf_c1bus_wb[4]_i_50 ),
        .\rgf_c1bus_wb[4]_i_50_0 (sreg_n_62),
        .\rgf_c1bus_wb[4]_i_50_1 (\rgf_c1bus_wb[4]_i_50_0 ),
        .\rgf_c1bus_wb[4]_i_50_2 (sreg_n_41),
        .\rgf_c1bus_wb[4]_i_52 (\rgf_c1bus_wb[4]_i_52 ),
        .\rgf_c1bus_wb[4]_i_52_0 (sreg_n_70),
        .\rgf_c1bus_wb[4]_i_52_1 (\rgf_c1bus_wb[4]_i_52_0 ),
        .\rgf_c1bus_wb[4]_i_52_2 (sreg_n_49),
        .\rgf_c1bus_wb[4]_i_54 (\rgf_c1bus_wb[4]_i_54 ),
        .\rgf_c1bus_wb[4]_i_54_0 (sreg_n_69),
        .\rgf_c1bus_wb[4]_i_54_1 (\rgf_c1bus_wb[4]_i_54_0 ),
        .\rgf_c1bus_wb[4]_i_54_2 (sreg_n_48),
        .\rgf_c1bus_wb[4]_i_56 (\rgf_c1bus_wb[4]_i_56 ),
        .\rgf_c1bus_wb[4]_i_56_0 (sreg_n_68),
        .\rgf_c1bus_wb[4]_i_56_1 (\rgf_c1bus_wb[4]_i_56_0 ),
        .\rgf_c1bus_wb[4]_i_56_2 (sreg_n_47),
        .\rgf_c1bus_wb[4]_i_58 (\rgf_c1bus_wb[4]_i_58 ),
        .\rgf_c1bus_wb[4]_i_58_0 (sreg_n_67),
        .\rgf_c1bus_wb[4]_i_58_1 (\rgf_c1bus_wb[4]_i_58_0 ),
        .\rgf_c1bus_wb[4]_i_58_2 (sreg_n_46),
        .\rgf_c1bus_wb[4]_i_60 (\rgf_c1bus_wb[4]_i_60 ),
        .\rgf_c1bus_wb[4]_i_60_0 (sreg_n_66),
        .\rgf_c1bus_wb[4]_i_60_1 (\rgf_c1bus_wb[4]_i_60_0 ),
        .\rgf_c1bus_wb[4]_i_60_2 (sreg_n_45),
        .\rgf_c1bus_wb[4]_i_62 (\rgf_c1bus_wb[4]_i_62 ),
        .\rgf_c1bus_wb[4]_i_62_0 (sreg_n_65),
        .\rgf_c1bus_wb[4]_i_62_1 (\rgf_c1bus_wb[4]_i_62_0 ),
        .\rgf_c1bus_wb[4]_i_62_2 (sreg_n_44),
        .\rgf_c1bus_wb[4]_i_64 (\rgf_c1bus_wb[4]_i_64 ),
        .\rgf_c1bus_wb[4]_i_64_0 (sreg_n_64),
        .\rgf_c1bus_wb[4]_i_64_1 (\rgf_c1bus_wb[4]_i_64_0 ),
        .\rgf_c1bus_wb[4]_i_64_2 (sreg_n_43),
        .rst_n(rst_n),
        .\sp_reg[11] (\sp_reg[11]_0 ),
        .\sp_reg[13] (\sp_reg[13]_0 ),
        .\sp_reg[14] (bank13_n_156),
        .\sp_reg[1] (\sp_reg[1]_1 ),
        .\sp_reg[2] (\sp_reg[2]_0 ),
        .\sp_reg[4] (\sp_reg[4]_0 ),
        .\sp_reg[6] (bank13_n_164),
        .\sr[4]_i_129 (\sr[4]_i_129 ),
        .\sr[4]_i_133_0 (\sr[4]_i_133 ),
        .\sr[4]_i_138_0 (\sr_reg[6]_29 ),
        .\sr[4]_i_138_1 (a0bus_0[15]),
        .\sr[4]_i_139 (\rgf_c0bus_wb_reg[10]_1 ),
        .\sr[4]_i_139_0 (\rgf_c0bus_wb[3]_i_7 ),
        .\sr[4]_i_15 (\sr[4]_i_15 ),
        .\sr[4]_i_154_0 (a1bus_out_n_20),
        .\sr[4]_i_154_1 (a1bus_out_n_18),
        .\sr[4]_i_155_0 (a1bus_out_n_62),
        .\sr[4]_i_155_1 (a1bus_out_n_63),
        .\sr[4]_i_155_10 (a1bus_out_n_58),
        .\sr[4]_i_155_11 (a1bus_out_n_26),
        .\sr[4]_i_155_2 (a1bus_out_n_61),
        .\sr[4]_i_155_3 (a1bus_out_n_34),
        .\sr[4]_i_155_4 (a1bus_out_n_60),
        .\sr[4]_i_155_5 (a1bus_out_n_32),
        .\sr[4]_i_155_6 (a1bus_out_n_40),
        .\sr[4]_i_155_7 (a1bus_out_n_38),
        .\sr[4]_i_155_8 (a1bus_out_n_59),
        .\sr[4]_i_155_9 (a1bus_out_n_28),
        .\sr[4]_i_156_0 (\sr[4]_i_156 ),
        .\sr[4]_i_159_0 (a1bus_out_n_54),
        .\sr[4]_i_159_1 (a1bus_out_n_56),
        .\sr[4]_i_159_2 (a1bus_out_n_55),
        .\sr[4]_i_159_3 (a1bus_out_n_57),
        .\sr[4]_i_159_4 (a1bus_out_n_23),
        .\sr[4]_i_159_5 (a1bus_out_n_21),
        .\sr[4]_i_159_6 (a1bus_out_n_17),
        .\sr[4]_i_159_7 (a1bus_out_n_15),
        .\sr[4]_i_15_0 (\sr[4]_i_15_0 ),
        .\sr[4]_i_15_1 (\sr[4]_i_15_1 ),
        .\sr[4]_i_164_0 (a1bus_out_n_64),
        .\sr[4]_i_164_1 (a1bus_out_n_65),
        .\sr[4]_i_164_2 (a1bus_out_n_46),
        .\sr[4]_i_164_3 (a1bus_out_n_44),
        .\sr[4]_i_168 (a1bus_out_n_8),
        .\sr[4]_i_168_0 (a1bus_out_n_12),
        .\sr[4]_i_168_1 (a1bus_out_n_51),
        .\sr[4]_i_168_2 (a1bus_out_n_6),
        .\sr[4]_i_168_3 (a1bus_out_n_14),
        .\sr[4]_i_170 (a1bus_out_n_43),
        .\sr[4]_i_170_0 (\sr[6]_i_11 ),
        .\sr[4]_i_170_1 (a1bus_out_n_48),
        .\sr[4]_i_170_2 (a1bus_out_n_37),
        .\sr[4]_i_170_3 (a1bus_out_n_41),
        .\sr[4]_i_183_0 (a0bus_out_n_47),
        .\sr[4]_i_183_1 (a0bus_out_n_51),
        .\sr[4]_i_183_10 (a0bus_out_n_58),
        .\sr[4]_i_183_11 (a0bus_out_n_57),
        .\sr[4]_i_183_12 (a0bus_out_n_77),
        .\sr[4]_i_183_13 (a0bus_out_n_34),
        .\sr[4]_i_183_14 (a0bus_out_n_33),
        .\sr[4]_i_183_15 (a0bus_out_n_35),
        .\sr[4]_i_183_16 (a0bus_out_n_42),
        .\sr[4]_i_183_17 (a0bus_out_n_41),
        .\sr[4]_i_183_18 (a0bus_out_n_73),
        .\sr[4]_i_183_19 (a0bus_out_n_79),
        .\sr[4]_i_183_2 (a0bus_out_n_39),
        .\sr[4]_i_183_3 (a0bus_out_n_43),
        .\sr[4]_i_183_4 (a0bus_out_n_63),
        .\sr[4]_i_183_5 (a0bus_out_n_55),
        .\sr[4]_i_183_6 (a0bus_out_n_59),
        .\sr[4]_i_183_7 (a0bus_out_n_50),
        .\sr[4]_i_183_8 (a0bus_out_n_49),
        .\sr[4]_i_183_9 (a0bus_out_n_75),
        .\sr[4]_i_185 (\rgf_c0bus_wb[3]_i_7_0 ),
        .\sr[4]_i_185_0 (a0bus_out_n_65),
        .\sr[4]_i_186_0 (a0bus_out_n_38),
        .\sr[4]_i_186_1 (a0bus_out_n_37),
        .\sr[4]_i_186_2 (a0bus_out_n_30),
        .\sr[4]_i_186_3 (a0bus_out_n_29),
        .\sr[4]_i_186_4 (a0bus_out_n_70),
        .\sr[4]_i_186_5 (a0bus_out_n_72),
        .\sr[4]_i_194_0 (a0bus_out_n_14),
        .\sr[4]_i_194_1 (a0bus_out_n_13),
        .\sr[4]_i_194_2 (a0bus_out_n_66),
        .\sr[4]_i_194_3 (a0bus_out_n_22),
        .\sr[4]_i_194_4 (a0bus_out_n_21),
        .\sr[4]_i_194_5 (a0bus_out_n_68),
        .\sr[4]_i_195_0 (\sr[4]_i_195 ),
        .\sr[4]_i_197_0 (a0bus_out_n_10),
        .\sr[4]_i_197_1 (a0bus_out_n_9),
        .\sr[4]_i_197_2 (a0bus_out_n_11),
        .\sr[4]_i_197_3 (\sp_reg[0]_0 ),
        .\sr[4]_i_197_4 (\sr_reg[0] ),
        .\sr[4]_i_197_5 ({\sr_reg[15] [6],\sr_reg[15] [1:0]}),
        .\sr[4]_i_197_6 (a0bus_out_n_67),
        .\sr[4]_i_197_7 (a0bus_out_n_15),
        .\sr[4]_i_200_0 (\sr[4]_i_200 ),
        .\sr[4]_i_232_0 (\sr[4]_i_232 ),
        .\sr[4]_i_239 (\sr[4]_i_239 ),
        .\sr[4]_i_239_0 (sreg_n_75),
        .\sr[4]_i_27 (\sr[4]_i_27 ),
        .\sr[4]_i_27_0 (\rgf_c1bus_wb_reg[5]_1 ),
        .\sr[4]_i_27_1 (\rgf_c1bus_wb_reg[5] ),
        .\sr[4]_i_57_0 (\rgf_c0bus_wb[11]_i_9 ),
        .\sr[4]_i_57_1 (\rgf_c0bus_wb_reg[10] ),
        .\sr[4]_i_57_2 (\rgf_c0bus_wb[14]_i_2 ),
        .\sr[4]_i_57_3 (\rgf_c0bus_wb[11]_i_9_0 ),
        .\sr[4]_i_66 (\sr[4]_i_66 ),
        .\sr[4]_i_66_0 (\sr[4]_i_67 ),
        .\sr[4]_i_67 (bank02_n_264),
        .\sr[4]_i_67_0 (\rgf_c0bus_wb_reg[10]_0 ),
        .\sr[4]_i_80_0 (\sr[6]_i_11_0 ),
        .\sr[4]_i_80_1 (a1bus_0[15]),
        .\sr[4]_i_80_2 (\rgf_c1bus_wb_reg[7] ),
        .\sr[4]_i_83 (sreg_n_18),
        .\sr[4]_i_90 (\rgf_c1bus_wb[12]_i_2 ),
        .\sr_reg[6] (bank13_n_130),
        .\sr_reg[6]_0 (\sr_reg[6]_16 ),
        .\sr_reg[6]_1 (\sr_reg[6]_19 ),
        .\sr_reg[6]_2 (\sr_reg[6]_25 ),
        .\sr_reg[6]_3 (\sr_reg[6]_26 ),
        .\sr_reg[6]_4 (\sr_reg[6]_27 ),
        .\sr_reg[6]_5 (\sr_reg[6]_35 ),
        .\tr_reg[11] (\tr_reg[11]_0 ),
        .\tr_reg[12] (\tr_reg[12]_1 ),
        .\tr_reg[13] (\tr_reg[13]_1 ),
        .\tr_reg[13]_0 (bank13_n_138),
        .\tr_reg[14] (\tr_reg[14]_2 ),
        .\tr_reg[1] (\tr_reg[1] ),
        .\tr_reg[1]_0 (\tr_reg[1]_0 ),
        .\tr_reg[3] (\tr_reg[3] ));
  mcss_rgf_ivec ivec
       (.SR(SR),
        .clk(clk),
        .\iv_reg[15]_0 (\iv_reg[15]_1 ),
        .out(\iv_reg[15] ));
  mcss_rgf_pcnt pcnt
       (.D(D),
        .O(O),
        .S(S),
        .SR(SR),
        .clk(clk),
        .fadr(fadr),
        .\fadr[15] (\fadr[15] ),
        .\fadr[15]_0 (\fadr[15]_0 ),
        .out(\pc_reg[15] ),
        .\pc0_reg[15] (\pc0_reg[15] ),
        .\pc0_reg[15]_0 (\pc0_reg[15]_0 ),
        .\pc0_reg[15]_1 (fch_irq_req),
        .\pc0_reg[15]_2 (\pc0_reg[15]_1 ),
        .\pc_reg[13]_0 (\pc_reg[13] ),
        .\pc_reg[13]_1 (\pc_reg[13]_0 ),
        .\pc_reg[14]_0 (\pc_reg[14] ),
        .\pc_reg[15]_0 (\pc_reg[15]_0 ),
        .\pc_reg[15]_1 (\pc_reg[15]_1 ),
        .\pc_reg[15]_2 (\pc_reg[15]_2 ),
        .\pc_reg[1]_0 (\pc_reg[1] ));
  mcss_rgf_ctl rctl
       (.E(E),
        .bank_sel(bank_sel),
        .clk(clk),
        .out(\sr_reg[15] [1:0]),
        .p_2_in(p_2_in),
        .\rgf_c0bus_wb_reg[15]_0 (\rgf_c0bus_wb_reg[15] ),
        .\rgf_c0bus_wb_reg[15]_1 (\rgf_c0bus_wb_reg[15]_0 ),
        .\rgf_c1bus_wb_reg[0]_0 (\rgf_c1bus_wb_reg[0] ),
        .\rgf_c1bus_wb_reg[15]_0 (\rgf_c1bus_wb_reg[15] ),
        .\rgf_c1bus_wb_reg[15]_1 (\rgf_c1bus_wb_reg[15]_0 ),
        .\rgf_selc0_rn_wb_reg[2]_0 (\rgf_selc0_rn_wb_reg[2] ),
        .\rgf_selc0_rn_wb_reg[2]_1 (\rgf_selc0_rn_wb_reg[2]_0 ),
        .rgf_selc0_stat(rgf_selc0_stat),
        .\rgf_selc0_wb_reg[1]_0 (\rgf_selc0_wb_reg[1] ),
        .\rgf_selc0_wb_reg[1]_1 (\rgf_selc0_wb_reg[1]_0 ),
        .\rgf_selc1_rn_wb_reg[2]_0 (\rgf_selc1_rn_wb_reg[2] ),
        .\rgf_selc1_rn_wb_reg[2]_1 (\rgf_selc1_rn_wb_reg[2]_0 ),
        .rgf_selc1_stat(rgf_selc1_stat),
        .rgf_selc1_stat_reg_0(rgf_selc1_stat_reg),
        .\rgf_selc1_wb_reg[0]_0 (\rgf_selc1_wb_reg[0] ),
        .\rgf_selc1_wb_reg[1]_0 (\rgf_selc1_wb_reg[1] ),
        .\rgf_selc1_wb_reg[1]_1 (\rgf_selc1_wb_reg[1]_0 ),
        .rst_n(rst_n),
        .\sr_reg[0] (\sr_reg[0]_1 ));
  mcss_rgf_sptr sptr
       (.O(\sp_reg[1] ),
        .SR(SR),
        .clk(clk),
        .data3(data3),
        .out({p_0_in_2,\sp_reg[0] }),
        .\sp_reg[10]_0 (\sp_reg[10] ),
        .\sp_reg[11]_0 (\sp_reg[11] ),
        .\sp_reg[12]_0 (\sp_reg[12] ),
        .\sp_reg[13]_0 (\sp_reg[13] ),
        .\sp_reg[14]_0 (\sp_reg[14] ),
        .\sp_reg[14]_1 (\sp_reg[14]_0 ),
        .\sp_reg[14]_2 (\sp_reg[14]_1 ),
        .\sp_reg[15]_0 (\sp_reg[15] ),
        .\sp_reg[15]_1 (\sp_reg[15]_1 ),
        .\sp_reg[1]_0 (\sp_reg[1]_0 ),
        .\sp_reg[2]_0 (\sp_reg[2] ),
        .\sp_reg[3]_0 (\sp_reg[3] ),
        .\sp_reg[4]_0 (\sp_reg[4] ),
        .\sp_reg[5]_0 (\sp_reg[5] ),
        .\sp_reg[6]_0 (\sp_reg[6] ),
        .\sp_reg[7]_0 (\sp_reg[7] ),
        .\sp_reg[8]_0 (\sp_reg[8] ),
        .\sp_reg[9]_0 (\sp_reg[9] ));
  mcss_rgf_sreg sreg
       (.Q(Q),
        .a1bus_sel_0(a1bus_sel_0[2:1]),
        .b0bus_sel_0(b0bus_sel_0[0]),
        .\badr[15]_INST_0_i_208 (\badr[15]_INST_0_i_208 ),
        .\badr[15]_INST_0_i_7 ({bank13_n_26,bank13_n_27,bank13_n_28,bank13_n_29,bank13_n_30,bank13_n_31,bank13_n_32,bank13_n_33,bank13_n_34,bank13_n_35,bank13_n_36,\grn_reg[4]_1 }),
        .\badr[15]_INST_0_i_7_0 ({bank13_n_42,bank13_n_43,bank13_n_44,bank13_n_45,bank13_n_46,bank13_n_47,bank13_n_48,bank13_n_49,bank13_n_50,bank13_n_51,bank13_n_52,\grn_reg[4]_2 }),
        .clk(clk),
        .ctl_fetch1_fl_i_15(ctl_fetch1_fl_i_15),
        .fch_irq_req(fch_irq_req),
        .gr6_bus1(\a1buso2l/gr6_bus1 ),
        .gr6_bus1_0(\a1buso/gr6_bus1 ),
        .gr6_bus1_1(\a1buso2l/gr6_bus1_0 ),
        .\i_/bbus_o[4]_INST_0_i_5 ({bank02_n_52,bank02_n_53,bank02_n_54,bank02_n_55,bank02_n_56}),
        .\i_/bbus_o[4]_INST_0_i_6 ({bank02_n_15,bank02_n_16,bank02_n_17,bank02_n_18,bank02_n_19}),
        .irq(irq),
        .irq_0(irq_0),
        .irq_lev(irq_lev),
        .\rgf_c0bus_wb[0]_i_5 (\rgf_c0bus_wb_reg[10]_0 ),
        .\rgf_c0bus_wb[4]_i_10 (\sp_reg[0]_0 ),
        .\rgf_c0bus_wb[4]_i_10_0 (\sr_reg[0] ),
        .\rgf_c0bus_wb[4]_i_10_1 (a0bus_out_n_63),
        .\rgf_c1bus_wb[4]_i_39 ({bank02_n_20,bank02_n_21,bank02_n_22,bank02_n_23,bank02_n_24,bank02_n_25,bank02_n_26,bank02_n_27,bank02_n_28,bank02_n_29,bank02_n_30,bank02_n_31,bank02_n_32,bank02_n_33,bank02_n_34,bank02_n_35}),
        .\rgf_c1bus_wb[4]_i_39_0 ({bank02_n_36,bank02_n_37,bank02_n_38,bank02_n_39,bank02_n_40,bank02_n_41,bank02_n_42,bank02_n_43,bank02_n_44,bank02_n_45,bank02_n_46,bank02_n_47,bank02_n_48,bank02_n_49,bank02_n_50,bank02_n_51}),
        .\rgf_c1bus_wb[4]_i_45 ({bank13_n_89,bank13_n_90,bank13_n_91,bank13_n_92,bank13_n_93,bank13_n_94,bank13_n_95,bank13_n_96,bank13_n_97,bank13_n_98,bank13_n_99,\grn_reg[4]_6 }),
        .\rgf_c1bus_wb[4]_i_45_0 ({bank13_n_105,bank13_n_106,bank13_n_107,bank13_n_108,bank13_n_109,bank13_n_110,bank13_n_111,bank13_n_112,bank13_n_113,bank13_n_114,bank13_n_115,bank13_n_116,bank13_n_117,bank13_n_118,bank13_n_119,bank13_n_120}),
        .\rgf_c1bus_wb[4]_i_47 ({bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78,bank02_n_79,bank02_n_80,bank02_n_81,bank02_n_82,bank02_n_83,bank02_n_84,bank02_n_85,bank02_n_86,bank02_n_87,bank02_n_88}),
        .\rgf_c1bus_wb[4]_i_47_0 ({bank02_n_57,bank02_n_58,bank02_n_59,bank02_n_60,bank02_n_61,bank02_n_62,bank02_n_63,bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72}),
        .\rgf_selc1_wb[1]_i_16 (\rgf_selc1_wb[1]_i_16 ),
        .\sr[4]_i_160 (\sr[6]_i_11 ),
        .\sr[4]_i_160_0 (\tr_reg[15]_0 ),
        .\sr[4]_i_160_1 (\grn_reg[15]_1 ),
        .\sr[4]_i_160_2 (\sr_reg[15]_0 ),
        .\sr[4]_i_160_3 (\sp_reg[15]_0 ),
        .\sr[4]_i_172 (a1bus_out_n_46),
        .\sr[4]_i_172_0 (a1bus_b02[0]),
        .\sr[4]_i_172_1 (a1bus_out_n_66),
        .\sr[4]_i_172_2 (a1bus_out_n_47),
        .\sr[4]_i_188 (\rgf_c0bus_wb[3]_i_7_0 ),
        .\sr[4]_i_188_0 (a0bus_out_n_2),
        .\sr[4]_i_188_1 (a0bus_out_n_1),
        .\sr[4]_i_188_2 (a0bus_out_n_3),
        .\sr_reg[0]_0 (sreg_n_34),
        .\sr_reg[0]_1 (sreg_n_35),
        .\sr_reg[0]_10 (sreg_n_44),
        .\sr_reg[0]_11 (sreg_n_45),
        .\sr_reg[0]_12 (sreg_n_46),
        .\sr_reg[0]_13 (sreg_n_47),
        .\sr_reg[0]_14 (sreg_n_48),
        .\sr_reg[0]_15 (sreg_n_49),
        .\sr_reg[0]_16 (sreg_n_50),
        .\sr_reg[0]_17 (sreg_n_51),
        .\sr_reg[0]_18 (sreg_n_52),
        .\sr_reg[0]_19 (sreg_n_53),
        .\sr_reg[0]_2 (sreg_n_36),
        .\sr_reg[0]_20 (sreg_n_54),
        .\sr_reg[0]_21 (sreg_n_60),
        .\sr_reg[0]_22 (sreg_n_61),
        .\sr_reg[0]_23 (sreg_n_62),
        .\sr_reg[0]_24 (sreg_n_63),
        .\sr_reg[0]_25 (sreg_n_64),
        .\sr_reg[0]_26 (sreg_n_65),
        .\sr_reg[0]_27 (sreg_n_66),
        .\sr_reg[0]_28 (sreg_n_67),
        .\sr_reg[0]_29 (sreg_n_68),
        .\sr_reg[0]_3 (sreg_n_37),
        .\sr_reg[0]_30 (sreg_n_69),
        .\sr_reg[0]_31 (sreg_n_70),
        .\sr_reg[0]_32 (sreg_n_71),
        .\sr_reg[0]_33 (sreg_n_72),
        .\sr_reg[0]_34 (sreg_n_73),
        .\sr_reg[0]_35 (sreg_n_74),
        .\sr_reg[0]_36 (sreg_n_75),
        .\sr_reg[0]_37 (\sr_reg[0]_0 ),
        .\sr_reg[0]_38 (sreg_n_112),
        .\sr_reg[0]_39 (sreg_n_113),
        .\sr_reg[0]_4 (sreg_n_38),
        .\sr_reg[0]_40 (sreg_n_114),
        .\sr_reg[0]_41 (sreg_n_115),
        .\sr_reg[0]_42 (sreg_n_116),
        .\sr_reg[0]_43 (sreg_n_117),
        .\sr_reg[0]_44 (sreg_n_118),
        .\sr_reg[0]_45 (sreg_n_119),
        .\sr_reg[0]_46 (sreg_n_120),
        .\sr_reg[0]_47 (sreg_n_121),
        .\sr_reg[0]_48 (sreg_n_122),
        .\sr_reg[0]_49 (sreg_n_123),
        .\sr_reg[0]_5 (sreg_n_39),
        .\sr_reg[0]_50 (sreg_n_124),
        .\sr_reg[0]_51 (sreg_n_125),
        .\sr_reg[0]_52 (sreg_n_126),
        .\sr_reg[0]_53 (sreg_n_127),
        .\sr_reg[0]_6 (sreg_n_40),
        .\sr_reg[0]_7 (sreg_n_41),
        .\sr_reg[0]_8 (sreg_n_42),
        .\sr_reg[0]_9 (sreg_n_43),
        .\sr_reg[10]_0 (\sr_reg[10] ),
        .\sr_reg[15]_0 (\sr_reg[15] ),
        .\sr_reg[15]_1 (\sr_reg[15]_2 ),
        .\sr_reg[1]_0 (sreg_n_55),
        .\sr_reg[1]_1 (sreg_n_56),
        .\sr_reg[1]_10 (sreg_n_81),
        .\sr_reg[1]_11 (sreg_n_82),
        .\sr_reg[1]_12 (sreg_n_83),
        .\sr_reg[1]_13 (sreg_n_84),
        .\sr_reg[1]_14 (sreg_n_85),
        .\sr_reg[1]_15 (sreg_n_86),
        .\sr_reg[1]_16 (sreg_n_87),
        .\sr_reg[1]_17 (sreg_n_88),
        .\sr_reg[1]_18 (sreg_n_89),
        .\sr_reg[1]_19 (sreg_n_90),
        .\sr_reg[1]_2 (sreg_n_57),
        .\sr_reg[1]_20 (sreg_n_95),
        .\sr_reg[1]_21 (sreg_n_96),
        .\sr_reg[1]_22 (sreg_n_97),
        .\sr_reg[1]_23 (sreg_n_98),
        .\sr_reg[1]_24 (sreg_n_99),
        .\sr_reg[1]_25 (sreg_n_100),
        .\sr_reg[1]_26 (sreg_n_101),
        .\sr_reg[1]_27 (sreg_n_102),
        .\sr_reg[1]_28 (sreg_n_103),
        .\sr_reg[1]_29 (sreg_n_104),
        .\sr_reg[1]_3 (sreg_n_58),
        .\sr_reg[1]_30 (sreg_n_105),
        .\sr_reg[1]_31 (sreg_n_106),
        .\sr_reg[1]_32 (sreg_n_107),
        .\sr_reg[1]_33 (sreg_n_108),
        .\sr_reg[1]_34 (sreg_n_109),
        .\sr_reg[1]_35 (sreg_n_110),
        .\sr_reg[1]_36 (sreg_n_111),
        .\sr_reg[1]_37 (sreg_n_128),
        .\sr_reg[1]_38 (sreg_n_129),
        .\sr_reg[1]_39 (sreg_n_130),
        .\sr_reg[1]_4 (sreg_n_59),
        .\sr_reg[1]_40 (sreg_n_131),
        .\sr_reg[1]_41 (sreg_n_132),
        .\sr_reg[1]_42 (sreg_n_133),
        .\sr_reg[1]_43 (sreg_n_134),
        .\sr_reg[1]_44 (sreg_n_135),
        .\sr_reg[1]_45 (sreg_n_136),
        .\sr_reg[1]_46 (sreg_n_137),
        .\sr_reg[1]_47 (sreg_n_138),
        .\sr_reg[1]_48 (sreg_n_139),
        .\sr_reg[1]_49 (sreg_n_140),
        .\sr_reg[1]_5 (sreg_n_76),
        .\sr_reg[1]_50 (sreg_n_141),
        .\sr_reg[1]_51 (sreg_n_142),
        .\sr_reg[1]_52 (sreg_n_143),
        .\sr_reg[1]_53 (sreg_n_144),
        .\sr_reg[1]_54 (sreg_n_145),
        .\sr_reg[1]_55 (sreg_n_146),
        .\sr_reg[1]_56 (sreg_n_147),
        .\sr_reg[1]_57 (sreg_n_148),
        .\sr_reg[1]_58 (sreg_n_149),
        .\sr_reg[1]_59 (sreg_n_150),
        .\sr_reg[1]_6 (sreg_n_77),
        .\sr_reg[1]_60 (sreg_n_151),
        .\sr_reg[1]_61 (sreg_n_152),
        .\sr_reg[1]_62 (sreg_n_153),
        .\sr_reg[1]_63 (sreg_n_154),
        .\sr_reg[1]_64 (sreg_n_155),
        .\sr_reg[1]_65 (sreg_n_156),
        .\sr_reg[1]_66 (sreg_n_157),
        .\sr_reg[1]_67 (sreg_n_158),
        .\sr_reg[1]_68 (sreg_n_159),
        .\sr_reg[1]_7 (sreg_n_78),
        .\sr_reg[1]_8 (sreg_n_79),
        .\sr_reg[1]_9 (sreg_n_80),
        .\sr_reg[4]_0 (\sr_reg[4] ),
        .\sr_reg[4]_1 (\sr_reg[4]_0 ),
        .\sr_reg[4]_2 (\sr_reg[4]_1 ),
        .\sr_reg[5]_0 (\sr_reg[5] ),
        .\sr_reg[5]_1 (\sr_reg[5]_0 ),
        .\sr_reg[5]_2 (\sr_reg[5]_1 ),
        .\sr_reg[5]_3 (\sr_reg[5]_2 ),
        .\sr_reg[5]_4 (\sr_reg[5]_3 ),
        .\sr_reg[5]_5 (\sr_reg[5]_4 ),
        .\sr_reg[5]_6 (\sr_reg[5]_5 ),
        .\sr_reg[5]_7 (\sr_reg[5]_6 ),
        .\sr_reg[6]_0 (sreg_n_18),
        .\sr_reg[6]_1 (\sr_reg[6]_6 ),
        .\sr_reg[6]_2 (\sr_reg[6]_33 ),
        .\sr_reg[6]_3 (\sr_reg[6]_29 ),
        .\sr_reg[6]_4 (\sr_reg[6]_39 ),
        .\sr_reg[6]_5 (\sr_reg[6]_40 ),
        .\sr_reg[6]_6 (\sr_reg[6]_41 ),
        .\sr_reg[7]_0 (\sr_reg[7] ));
  mcss_rgf_treg treg
       (.SR(SR),
        .badrx(badrx),
        .badrx_15_sp_1(badrx_15_sn_1),
        .clk(clk),
        .out(\tr_reg[15] ),
        .\rgf_c1bus_wb[4]_i_13 (a1bus_out_n_46),
        .\rgf_c1bus_wb[4]_i_13_0 (a1bus_b02[0]),
        .\rgf_c1bus_wb[4]_i_13_1 (a1bus_out_n_66),
        .\rgf_c1bus_wb[4]_i_13_2 (a1bus_out_n_47),
        .\rgf_c1bus_wb[4]_i_13_3 (\sr[6]_i_11 ),
        .\rgf_c1bus_wb[4]_i_13_4 (\sr_reg[15] [6]),
        .\sr[4]_i_167 (\tr_reg[15]_0 ),
        .\sr[4]_i_167_0 (\grn_reg[15]_1 ),
        .\sr[4]_i_167_1 (\sr_reg[15]_0 ),
        .\sr[4]_i_167_2 (\sp_reg[15]_0 ),
        .\sr_reg[6] (\sr_reg[6]_18 ),
        .\sr_reg[6]_0 (\sr_reg[6]_8 ),
        .\tr_reg[15]_0 (\tr_reg[15]_2 ));
endmodule

module mcss_rgf_bank
   (.out({gr20[15],gr20[14],gr20[13],gr20[12],gr20[11],gr20[10],gr20[9],gr20[7],gr20[6],gr20[5],gr20[4],gr20[3],gr20[2],gr20[1],gr20[0]}),
    .\grn_reg[4] ({gr21[4],gr21[3],gr21[2],gr21[1],gr21[0]}),
    .\grn_reg[15] ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_0 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[4]_0 ({gr01[4],gr01[3],gr01[2],gr01[1],gr01[0]}),
    .\grn_reg[15]_1 ({gr05[15],gr05[14],gr05[13],gr05[12],gr05[11],gr05[10],gr05[9],gr05[8],gr05[7],gr05[6],gr05[5],gr05[4],gr05[3],gr05[2],gr05[1],gr05[0]}),
    .\grn_reg[15]_2 ({gr06[15],gr06[14],gr06[13],gr06[12],gr06[11],gr06[10],gr06[9],gr06[8],gr06[7],gr06[6],gr06[5],gr06[4],gr06[3],gr06[2],gr06[1],gr06[0]}),
    bdatw,
    \tr_reg[14] ,
    \tr_reg[14]_0 ,
    \stat_reg[1] ,
    \tr_reg[13] ,
    \tr_reg[13]_0 ,
    \stat_reg[1]_0 ,
    \tr_reg[12] ,
    \tr_reg[11] ,
    \tr_reg[10] ,
    \tr_reg[9] ,
    \tr_reg[8] ,
    \stat_reg[1]_1 ,
    \tr_reg[7] ,
    \tr_reg[7]_0 ,
    \stat_reg[2] ,
    \tr_reg[6] ,
    \badr[6]_INST_0_i_1 ,
    \tr_reg[6]_0 ,
    \stat_reg[2]_0 ,
    \tr_reg[5] ,
    \badr[5]_INST_0_i_1 ,
    \tr_reg[5]_0 ,
    \rgf_c1bus_wb[13]_i_9 ,
    \rgf_c1bus_wb[14]_i_30 ,
    \sr_reg[6] ,
    \badr[15]_INST_0_i_1 ,
    \sr_reg[6]_0 ,
    \sr_reg[6]_1 ,
    \badr[3]_INST_0_i_1 ,
    \badr[15]_INST_0_i_1_0 ,
    \badr[1]_INST_0_i_1 ,
    \sr_reg[6]_2 ,
    \badr[9]_INST_0_i_1 ,
    \sr_reg[6]_3 ,
    \rgf_c1bus_wb[15]_i_14 ,
    \badr[10]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1_0 ,
    \badr[2]_INST_0_i_1 ,
    \rgf_c1bus_wb[11]_i_13 ,
    \badr[10]_INST_0_i_1_0 ,
    \badr[14]_INST_0_i_1 ,
    \rgf_c1bus_wb[15]_i_14_0 ,
    \badr[3]_INST_0_i_1_0 ,
    \badr[7]_INST_0_i_1 ,
    \sr_reg[6]_4 ,
    \badr[6]_INST_0_i_1_1 ,
    \sr_reg[6]_5 ,
    \rgf_c1bus_wb[12]_i_20_0 ,
    \rgf_c1bus_wb[11]_i_10 ,
    \badr[15]_INST_0_i_1_1 ,
    \rgf_c1bus_wb[14]_i_28 ,
    \rgf_c1bus_wb[15]_i_14_1 ,
    \rgf_c1bus_wb[14]_i_28_0 ,
    \rgf_c1bus_wb[7]_i_4 ,
    \badr[5]_INST_0_i_1_0 ,
    \sr[4]_i_219_0 ,
    \tr_reg[12]_0 ,
    \rgf_c1bus_wb[11]_i_10_0 ,
    \rgf_c1bus_wb[4]_i_9 ,
    \badr[12]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_28_1 ,
    \badr[0]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_28_2 ,
    \rgf_c1bus_wb[9]_i_17_0 ,
    \badr[10]_INST_0_i_1_1 ,
    \rgf_c1bus_wb[14]_i_28_3 ,
    \rgf_c1bus_wb[13]_i_16 ,
    \rgf_c1bus_wb[14]_i_28_4 ,
    \rgf_c1bus_wb[4]_i_9_0 ,
    \sr_reg[6]_6 ,
    \tr_reg[14]_1 ,
    \sr_reg[6]_7 ,
    \sr_reg[6]_8 ,
    \rgf_c1bus_wb[15]_i_14_2 ,
    \badr[11]_INST_0_i_1 ,
    \sr_reg[6]_9 ,
    \sr_reg[6]_10 ,
    \badr[2]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[15]_i_14_3 ,
    \rgf_c1bus_wb[14]_i_28_5 ,
    \badr[9]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[14]_i_28_6 ,
    \rgf_c1bus_wb[14]_i_32 ,
    \badr[13]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1_1 ,
    \rgf_c1bus_wb[14]_i_32_0 ,
    \sr_reg[6]_11 ,
    \sr_reg[6]_12 ,
    \badr[14]_INST_0_i_1_0 ,
    \stat_reg[2]_1 ,
    \sr_reg[6]_13 ,
    \rgf_c1bus_wb[11]_i_10_1 ,
    \rgf_c1bus_wb[1]_i_14_0 ,
    \badr[6]_INST_0_i_1_2 ,
    \rgf_c1bus_wb[11]_i_10_2 ,
    \sr_reg[6]_14 ,
    \sr[4]_i_220 ,
    \rgf_c1bus_wb[11]_i_10_3 ,
    \rgf_c1bus_wb[11]_i_10_4 ,
    \rgf_c1bus_wb[15]_i_27 ,
    \grn_reg[14] ,
    \grn_reg[15]_3 ,
    \stat_reg[2]_2 ,
    \stat_reg[2]_3 ,
    \tr_reg[15] ,
    \tr_reg[12]_1 ,
    \tr_reg[11]_0 ,
    \tr_reg[10]_0 ,
    \tr_reg[9]_0 ,
    \tr_reg[8]_0 ,
    \rgf_c0bus_wb[15]_i_18 ,
    \rgf_c0bus_wb[11]_i_3 ,
    \rgf_c0bus_wb[11]_i_3_0 ,
    \badr[6]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_11 ,
    \badr[5]_INST_0_i_2 ,
    \badr[1]_INST_0_i_2 ,
    \badr[13]_INST_0_i_2 ,
    \badr[9]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_11_0 ,
    \rgf_c0bus_wb[11]_i_22 ,
    \badr[8]_INST_0_i_2 ,
    \badr[3]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_9 ,
    \badr[10]_INST_0_i_2 ,
    \badr[6]_INST_0_i_2_0 ,
    \badr[2]_INST_0_i_2 ,
    \rgf_c0bus_wb[15]_i_25_0 ,
    \rgf_c0bus_wb[11]_i_8 ,
    \badr[4]_INST_0_i_2 ,
    \rgf_c0bus_wb[0]_i_14 ,
    \sr_reg[6]_15 ,
    \sr_reg[6]_16 ,
    \badr[10]_INST_0_i_2_0 ,
    \badr[14]_INST_0_i_2 ,
    \rgf_c0bus_wb[13]_i_29 ,
    \badr[4]_INST_0_i_2_0 ,
    \badr[12]_INST_0_i_2 ,
    \badr[8]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[7]_i_7 ,
    \rgf_c0bus_wb[7]_i_7_0 ,
    \sr_reg[6]_17 ,
    \sr_reg[6]_18 ,
    \badr[14]_INST_0_i_2_0 ,
    \sr_reg[6]_19 ,
    \rgf_c0bus_wb[11]_i_11_1 ,
    \rgf_c0bus_wb[11]_i_9_0 ,
    \badr[6]_INST_0_i_2_1 ,
    \rgf_c0bus_wb[11]_i_11_2 ,
    \badr[13]_INST_0_i_2_0 ,
    \badr[5]_INST_0_i_2_0 ,
    \badr[9]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[15]_i_26 ,
    \sr_reg[6]_20 ,
    \badr[3]_INST_0_i_2_0 ,
    \badr[11]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_22_0 ,
    \badr[2]_INST_0_i_2_0 ,
    \sr_reg[6]_21 ,
    \rgf_c0bus_wb[12]_i_24 ,
    \rgf_c0bus_wb[12]_i_22_0 ,
    \sr_reg[14] ,
    \sr_reg[6]_22 ,
    \sr_reg[6]_23 ,
    \rgf_c0bus_wb[10]_i_8 ,
    \rgf_c0bus_wb[11]_i_9_1 ,
    \badr[1]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[13]_i_28 ,
    \badr[14]_INST_0_i_2_1 ,
    \rgf_c0bus_wb[8]_i_6_0 ,
    \rgf_c0bus_wb[12]_i_25_0 ,
    \sr_reg[6]_24 ,
    \sr_reg[6]_25 ,
    \sr_reg[6]_26 ,
    \badr[8]_INST_0_i_2_1 ,
    \badr[12]_INST_0_i_2_0 ,
    \sr_reg[6]_27 ,
    \sr_reg[15] ,
    \rgf_c0bus_wb[11]_i_3_1 ,
    \rgf_c1bus_wb[7]_i_4_0 ,
    \sr_reg[6]_28 ,
    \rgf_c1bus_wb[11]_i_10_5 ,
    \rgf_c0bus_wb[15]_i_6 ,
    \rgf_c0bus_wb[15]_i_6_0 ,
    \rgf_c0bus_wb[15]_i_6_1 ,
    bbus_o,
    \rgf_c0bus_wb[11]_i_3_2 ,
    \rgf_c0bus_wb[11]_i_9_2 ,
    \rgf_c0bus_wb[11]_i_9_3 ,
    \rgf_c0bus_wb[11]_i_9_4 ,
    \rgf_c0bus_wb[11]_i_3_3 ,
    \badr[14]_INST_0_i_1_1 ,
    \badr[13]_INST_0_i_1_0 ,
    \badr[14]_INST_0_i_2_2 ,
    \badr[6]_INST_0_i_1_3 ,
    tout__1_carry__0_i_1__0_0,
    \badr[10]_INST_0_i_1_2 ,
    tout__1_carry__1_i_1__0_0,
    p_1_in,
    \grn_reg[15]_4 ,
    \grn_reg[15]_5 ,
    \grn_reg[14]_0 ,
    \grn_reg[14]_1 ,
    \grn_reg[13] ,
    \grn_reg[13]_0 ,
    \grn_reg[12] ,
    \grn_reg[12]_0 ,
    \grn_reg[11] ,
    \grn_reg[11]_0 ,
    \grn_reg[10] ,
    \grn_reg[10]_0 ,
    \grn_reg[9] ,
    \grn_reg[9]_0 ,
    \grn_reg[8] ,
    \grn_reg[8]_0 ,
    \grn_reg[7] ,
    \grn_reg[7]_0 ,
    \grn_reg[6] ,
    \grn_reg[6]_0 ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[4]_2 ,
    \grn_reg[3] ,
    \grn_reg[3]_0 ,
    \grn_reg[2] ,
    \grn_reg[2]_0 ,
    \grn_reg[1] ,
    \grn_reg[1]_0 ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[0]_1 ,
    \grn_reg[4]_3 ,
    p_1_in1_in,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[14]_2 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_1 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_1 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_1 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_1 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_1 ,
    \grn_reg[9]_2 ,
    \grn_reg[7]_1 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_1 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_1 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_4 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_1 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_1 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_1 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_8 ,
    p_0_in,
    \grn_reg[15]_9 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_4 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_10 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_6 ,
    \grn_reg[4]_8 ,
    p_0_in0_in,
    \grn_reg[15]_11 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_9 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_7 ,
    \grn_reg[15]_12 ,
    gr6_bus1,
    \grn_reg[14]_7 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_8 ,
    \grn_reg[15]_13 ,
    b1bus_b02,
    \bdatw[13] ,
    \bdatw[13]_0 ,
    \bdatw[13]_1 ,
    \bdatw[14] ,
    \bdatw[14]_0 ,
    \bdatw[14]_1 ,
    \bdatw[14]_2 ,
    \bdatw[13]_2 ,
    \bdatw[13]_3 ,
    \bdatw[13]_4 ,
    \bdatw[13]_5 ,
    \bdatw[12] ,
    \bdatw[12]_0 ,
    \bdatw[12]_1 ,
    \bdatw[12]_2 ,
    \bdatw[11] ,
    \bdatw[11]_0 ,
    \bdatw[11]_1 ,
    \bdatw[11]_2 ,
    \bdatw[10] ,
    \bdatw[10]_0 ,
    \bdatw[10]_1 ,
    \bdatw[10]_2 ,
    \bdatw[9] ,
    \bdatw[9]_0 ,
    \bdatw[9]_1 ,
    \bdatw[9]_2 ,
    \bdatw[8] ,
    \bdatw[8]_0 ,
    \bdatw[8]_1 ,
    \bdatw[8]_2 ,
    \rgf_c1bus_wb[15]_i_19 ,
    \rgf_c1bus_wb[15]_i_19_0 ,
    \rgf_c1bus_wb[15]_i_19_1 ,
    \rgf_c1bus_wb[15]_i_19_2 ,
    \sr[4]_i_77 ,
    \rgf_c1bus_wb_reg[5] ,
    \sr[6]_i_15 ,
    \sr[6]_i_11 ,
    \rgf_c1bus_wb[5]_i_10 ,
    \rgf_c1bus_wb[14]_i_11 ,
    \rgf_c1bus_wb[14]_i_11_0 ,
    \rgf_c1bus_wb[14]_i_11_1 ,
    \rgf_c1bus_wb[14]_i_11_2 ,
    \sr[6]_i_11_0 ,
    \sr[4]_i_77_0 ,
    tout__1_carry__0_i_7__0,
    tout__1_carry__0_i_7__0_0,
    tout__1_carry__0_i_7__0_1,
    tout__1_carry__0_i_7__0_2,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[5]_1 ,
    \rgf_c1bus_wb_reg[7] ,
    \sr[6]_i_11_1 ,
    \sr[6]_i_11_2 ,
    \sr[4]_i_77_1 ,
    \sr[6]_i_11_3 ,
    \sr[6]_i_11_4 ,
    \sr[6]_i_11_5 ,
    \sr[6]_i_11_6 ,
    \sr[4]_i_30 ,
    \sr[6]_i_11_7 ,
    \sr[4]_i_30_0 ,
    \sr[4]_i_102 ,
    \sr[4]_i_77_2 ,
    \rgf_c1bus_wb_reg[3] ,
    \sr[6]_i_11_8 ,
    \sr[6]_i_11_9 ,
    \sr[4]_i_99 ,
    \sr[4]_i_99_0 ,
    \sr[4]_i_99_1 ,
    \sr[4]_i_99_2 ,
    \sr[4]_i_38 ,
    \rgf_c1bus_wb_reg[4] ,
    \sr[4]_i_119 ,
    \rgf_c1bus_wb[12]_i_2 ,
    \sr[4]_i_88 ,
    \sr[4]_i_88_0 ,
    \sr[4]_i_44 ,
    \rgf_c1bus_wb_reg[10] ,
    \sr[4]_i_102_0 ,
    \sr[4]_i_111 ,
    \sr[4]_i_84 ,
    \sr[4]_i_177 ,
    \sr[4]_i_177_0 ,
    \sr[4]_i_177_1 ,
    \sr[4]_i_177_2 ,
    \sr[4]_i_171 ,
    \sr[4]_i_171_0 ,
    \sr[4]_i_171_1 ,
    \sr[4]_i_171_2 ,
    \sr[4]_i_169_0 ,
    \sr[4]_i_169_1 ,
    \sr[4]_i_169_2 ,
    \sr[4]_i_179_0 ,
    \sr[4]_i_169_3 ,
    \sr[4]_i_169_4 ,
    \sr[4]_i_169_5 ,
    \sr[4]_i_169_6 ,
    \sr[4]_i_175_0 ,
    \sr[4]_i_179_1 ,
    \sr[4]_i_175_1 ,
    \sr[4]_i_175_2 ,
    \sr[4]_i_169_7 ,
    \sr[4]_i_179_2 ,
    \sr[4]_i_169_8 ,
    \sr[4]_i_179_3 ,
    \sr[4]_i_175_3 ,
    \sr[4]_i_175_4 ,
    \sr[4]_i_175_5 ,
    \sr[4]_i_175_6 ,
    \sr[4]_i_179_4 ,
    \sr[4]_i_179_5 ,
    \sr[4]_i_179_6 ,
    \sr[4]_i_179_7 ,
    \rgf_c1bus_wb[4]_i_7 ,
    \rgf_c1bus_wb[4]_i_7_0 ,
    \rgf_c1bus_wb[4]_i_7_1 ,
    \bdatw[15] ,
    \bdatw[15]_0 ,
    \bdatw[15]_1 ,
    \bdatw[15]_2 ,
    \bdatw[14]_3 ,
    \bdatw[14]_4 ,
    \bdatw[14]_5 ,
    \bdatw[14]_6 ,
    \bdatw[13]_6 ,
    \bdatw[13]_7 ,
    \bdatw[13]_8 ,
    \bdatw[13]_9 ,
    \bdatw[12]_3 ,
    \bdatw[12]_4 ,
    \bdatw[12]_5 ,
    \bdatw[12]_6 ,
    \bdatw[11]_3 ,
    \bdatw[11]_4 ,
    \bdatw[11]_5 ,
    \bdatw[11]_6 ,
    \bdatw[10]_3 ,
    \bdatw[10]_4 ,
    \bdatw[10]_5 ,
    \bdatw[10]_6 ,
    \bdatw[9]_3 ,
    \bdatw[9]_4 ,
    \bdatw[9]_5 ,
    \bdatw[9]_6 ,
    \bdatw[8]_3 ,
    \bdatw[8]_4 ,
    \bdatw[8]_5 ,
    \bdatw[8]_6 ,
    \rgf_c0bus_wb_reg[7]_i_11 ,
    \sr[4]_i_67 ,
    \rgf_c0bus_wb[6]_i_11 ,
    \rgf_c0bus_wb[14]_i_13 ,
    \rgf_c0bus_wb[3]_i_7 ,
    \rgf_c0bus_wb[14]_i_13_0 ,
    \rgf_c0bus_wb[14]_i_2 ,
    \bbus_o[7] ,
    \bbus_o[7]_0 ,
    \bbus_o[7]_1 ,
    \bbus_o[7]_2 ,
    \rgf_c0bus_wb[3]_i_18 ,
    \bbus_o[6] ,
    \bbus_o[6]_0 ,
    \bbus_o[6]_1 ,
    \bbus_o[6]_2 ,
    \bbus_o[5] ,
    \bbus_o[5]_0 ,
    \bbus_o[5]_1 ,
    \bbus_o[5]_2 ,
    \rgf_c0bus_wb_reg[10] ,
    \rgf_c0bus_wb_reg[10]_0 ,
    \rgf_c0bus_wb[12]_i_2 ,
    \sr[4]_i_55 ,
    \rgf_c0bus_wb[13]_i_4 ,
    \rgf_c0bus_wb[10]_i_4 ,
    \rgf_c0bus_wb_reg[10]_1 ,
    \rgf_c0bus_wb[14]_i_13_1 ,
    \rgf_c0bus_wb[14]_i_13_2 ,
    \rgf_c0bus_wb[3]_i_7_0 ,
    \rgf_c0bus_wb[3]_i_7_1 ,
    \rgf_c0bus_wb[14]_i_13_3 ,
    \rgf_c0bus_wb[14]_i_13_4 ,
    \rgf_c0bus_wb[14]_i_13_5 ,
    \rgf_c0bus_wb[12]_i_10 ,
    \rgf_c0bus_wb[14]_i_13_6 ,
    \rgf_c0bus_wb[3]_i_7_2 ,
    \rgf_c0bus_wb[3]_i_7_3 ,
    \rgf_c0bus_wb[3]_i_7_4 ,
    \rgf_c0bus_wb[3]_i_18_0 ,
    \rgf_c0bus_wb[8]_i_2 ,
    \sr[4]_i_139 ,
    \rgf_c0bus_wb[12]_i_7 ,
    \sr[4]_i_126 ,
    \rgf_c0bus_wb[15]_i_14 ,
    \sr[4]_i_203_0 ,
    \sr[4]_i_203_1 ,
    \sr[4]_i_203_2 ,
    \sr[4]_i_203_3 ,
    \sr[4]_i_203_4 ,
    \rgf_c0bus_wb[4]_i_7 ,
    \sr[4]_i_188 ,
    \sr[4]_i_188_0 ,
    \sr[4]_i_188_1 ,
    \sr[4]_i_188_2 ,
    \sr[4]_i_196_0 ,
    \sr[4]_i_196_1 ,
    \sr[4]_i_196_2 ,
    \sr[4]_i_196_3 ,
    \sr[4]_i_196_4 ,
    \sr[4]_i_196_5 ,
    \sr[4]_i_196_6 ,
    \sr[4]_i_196_7 ,
    \sr[4]_i_196_8 ,
    \sr[4]_i_196_9 ,
    \rgf_c0bus_wb[4]_i_7_0 ,
    \rgf_c0bus_wb[4]_i_7_1 ,
    \rgf_c0bus_wb[4]_i_7_2 ,
    \rgf_c0bus_wb[4]_i_7_3 ,
    \bbus_o[5]_3 ,
    \rgf_c0bus_wb[4]_i_3 ,
    tout__1_carry__2,
    tout__1_carry__2_0,
    tout__1_carry__2_1,
    a0bus_sel_0,
    bank_sel,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_43 ,
    ctl_sela0,
    \i_/badr[15]_INST_0_i_43_0 ,
    \bbus_o[4]_INST_0_i_1 ,
    \bbus_o[3]_INST_0_i_1 ,
    \bbus_o[2]_INST_0_i_1 ,
    \bbus_o[1]_INST_0_i_1 ,
    \bbus_o[0]_INST_0_i_1 ,
    \i_/bdatw[15]_INST_0_i_9 ,
    \i_/bdatw[15]_INST_0_i_9_0 ,
    \i_/bdatw[15]_INST_0_i_9_1 ,
    \i_/bdatw[15]_INST_0_i_9_2 ,
    ctl_selb0_0,
    \i_/bdatw[15]_INST_0_i_24 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_77 ,
    b0bus_sel_0,
    \i_/bdatw[15]_INST_0_i_9_3 ,
    \i_/bdatw[15]_INST_0_i_24_0 ,
    \rgf_c1bus_wb[4]_i_22 ,
    \rgf_c1bus_wb[4]_i_23 ,
    \sr[4]_i_209 ,
    \rgf_c1bus_wb[4]_i_24 ,
    \sr[4]_i_207 ,
    \rgf_c1bus_wb[4]_i_28 ,
    \sr[4]_i_208 ,
    \rgf_c1bus_wb[4]_i_27 ,
    \sr[4]_i_225_0 ,
    \rgf_c1bus_wb[4]_i_26 ,
    \sr[4]_i_224_0 ,
    \rgf_c1bus_wb[4]_i_25 ,
    \sr[4]_i_220_0 ,
    \sr[4]_i_211 ,
    \sr[4]_i_213 ,
    \sr[4]_i_210 ,
    \i_/badr[15]_INST_0_i_19 ,
    \i_/badr[15]_INST_0_i_19_0 ,
    \i_/badr[15]_INST_0_i_19_1 ,
    a1bus_sel_0,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_113 ,
    \i_/bdatw[15]_INST_0_i_44 ,
    \i_/bdatw[15]_INST_0_i_112 ,
    \i_/bdatw[15]_INST_0_i_112_0 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_112_1 ,
    \i_/badr[15]_INST_0_i_47 ,
    \bbus_o[4]_INST_0_i_1_0 ,
    \bbus_o[3]_INST_0_i_1_0 ,
    \bbus_o[2]_INST_0_i_1_0 ,
    \bbus_o[1]_INST_0_i_1_0 ,
    \bbus_o[0]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[4]_i_22_0 ,
    \rgf_c1bus_wb[4]_i_23_0 ,
    \sr[4]_i_209_0 ,
    \rgf_c1bus_wb[4]_i_24_0 ,
    \sr[4]_i_207_0 ,
    \rgf_c1bus_wb[4]_i_28_0 ,
    \sr[4]_i_208_0 ,
    \rgf_c1bus_wb[4]_i_27_0 ,
    \sr[4]_i_225_1 ,
    \rgf_c1bus_wb[4]_i_26_0 ,
    \sr[4]_i_224_1 ,
    \rgf_c1bus_wb[4]_i_25_0 ,
    \sr[4]_i_220_1 ,
    \sr[4]_i_211_0 ,
    \sr[4]_i_213_0 ,
    \sr[4]_i_210_0 ,
    \rgf_c1bus_wb[4]_i_47 ,
    \rgf_c1bus_wb[4]_i_47_0 ,
    \rgf_c1bus_wb[4]_i_41 ,
    \rgf_c1bus_wb[4]_i_41_0 ,
    \rgf_c1bus_wb[4]_i_51 ,
    \rgf_c1bus_wb[4]_i_51_0 ,
    \sr[4]_i_235 ,
    \sr[4]_i_235_0 ,
    \rgf_c1bus_wb[4]_i_65 ,
    \rgf_c1bus_wb[4]_i_65_0 ,
    \sr[4]_i_237 ,
    \sr[4]_i_237_0 ,
    \rgf_c1bus_wb[4]_i_61 ,
    \rgf_c1bus_wb[4]_i_61_0 ,
    \rgf_c1bus_wb[4]_i_57 ,
    \rgf_c1bus_wb[4]_i_57_0 ,
    \sr[4]_i_245 ,
    \sr[4]_i_245_0 ,
    \rgf_c1bus_wb[4]_i_53 ,
    \rgf_c1bus_wb[4]_i_53_0 ,
    \sr[4]_i_243 ,
    \sr[4]_i_243_0 ,
    \rgf_c1bus_wb[4]_i_33 ,
    \rgf_c1bus_wb[4]_i_33_0 ,
    \rgf_c1bus_wb[4]_i_67 ,
    \rgf_c1bus_wb[4]_i_67_0 ,
    \rgf_c1bus_wb[4]_i_37 ,
    \rgf_c1bus_wb[4]_i_37_0 ,
    \sr[4]_i_240 ,
    \sr[4]_i_240_0 ,
    SR,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    clk,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 );
  output [1:0]bdatw;
  output \tr_reg[14] ;
  output \tr_reg[14]_0 ;
  output \stat_reg[1] ;
  output \tr_reg[13] ;
  output \tr_reg[13]_0 ;
  output \stat_reg[1]_0 ;
  output \tr_reg[12] ;
  output \tr_reg[11] ;
  output \tr_reg[10] ;
  output \tr_reg[9] ;
  output \tr_reg[8] ;
  output \stat_reg[1]_1 ;
  output \tr_reg[7] ;
  output \tr_reg[7]_0 ;
  output \stat_reg[2] ;
  output \tr_reg[6] ;
  output \badr[6]_INST_0_i_1 ;
  output \tr_reg[6]_0 ;
  output \stat_reg[2]_0 ;
  output \tr_reg[5] ;
  output \badr[5]_INST_0_i_1 ;
  output \tr_reg[5]_0 ;
  output \rgf_c1bus_wb[13]_i_9 ;
  output \rgf_c1bus_wb[14]_i_30 ;
  output \sr_reg[6] ;
  output \badr[15]_INST_0_i_1 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[6]_1 ;
  output \badr[3]_INST_0_i_1 ;
  output \badr[15]_INST_0_i_1_0 ;
  output \badr[1]_INST_0_i_1 ;
  output \sr_reg[6]_2 ;
  output \badr[9]_INST_0_i_1 ;
  output \sr_reg[6]_3 ;
  output \rgf_c1bus_wb[15]_i_14 ;
  output \badr[10]_INST_0_i_1 ;
  output \badr[6]_INST_0_i_1_0 ;
  output \badr[2]_INST_0_i_1 ;
  output \rgf_c1bus_wb[11]_i_13 ;
  output \badr[10]_INST_0_i_1_0 ;
  output \badr[14]_INST_0_i_1 ;
  output \rgf_c1bus_wb[15]_i_14_0 ;
  output \badr[3]_INST_0_i_1_0 ;
  output \badr[7]_INST_0_i_1 ;
  output \sr_reg[6]_4 ;
  output \badr[6]_INST_0_i_1_1 ;
  output \sr_reg[6]_5 ;
  output \rgf_c1bus_wb[12]_i_20_0 ;
  output \rgf_c1bus_wb[11]_i_10 ;
  output \badr[15]_INST_0_i_1_1 ;
  output \rgf_c1bus_wb[14]_i_28 ;
  output \rgf_c1bus_wb[15]_i_14_1 ;
  output \rgf_c1bus_wb[14]_i_28_0 ;
  output \rgf_c1bus_wb[7]_i_4 ;
  output \badr[5]_INST_0_i_1_0 ;
  output \sr[4]_i_219_0 ;
  output \tr_reg[12]_0 ;
  output \rgf_c1bus_wb[11]_i_10_0 ;
  output \rgf_c1bus_wb[4]_i_9 ;
  output \badr[12]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_28_1 ;
  output \badr[0]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_28_2 ;
  output \rgf_c1bus_wb[9]_i_17_0 ;
  output \badr[10]_INST_0_i_1_1 ;
  output \rgf_c1bus_wb[14]_i_28_3 ;
  output \rgf_c1bus_wb[13]_i_16 ;
  output \rgf_c1bus_wb[14]_i_28_4 ;
  output \rgf_c1bus_wb[4]_i_9_0 ;
  output \sr_reg[6]_6 ;
  output \tr_reg[14]_1 ;
  output \sr_reg[6]_7 ;
  output \sr_reg[6]_8 ;
  output \rgf_c1bus_wb[15]_i_14_2 ;
  output \badr[11]_INST_0_i_1 ;
  output \sr_reg[6]_9 ;
  output \sr_reg[6]_10 ;
  output \badr[2]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[15]_i_14_3 ;
  output \rgf_c1bus_wb[14]_i_28_5 ;
  output \badr[9]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[14]_i_28_6 ;
  output \rgf_c1bus_wb[14]_i_32 ;
  output \badr[13]_INST_0_i_1 ;
  output \badr[2]_INST_0_i_1_1 ;
  output \rgf_c1bus_wb[14]_i_32_0 ;
  output \sr_reg[6]_11 ;
  output \sr_reg[6]_12 ;
  output \badr[14]_INST_0_i_1_0 ;
  output \stat_reg[2]_1 ;
  output \sr_reg[6]_13 ;
  output \rgf_c1bus_wb[11]_i_10_1 ;
  output \rgf_c1bus_wb[1]_i_14_0 ;
  output \badr[6]_INST_0_i_1_2 ;
  output \rgf_c1bus_wb[11]_i_10_2 ;
  output \sr_reg[6]_14 ;
  output \sr[4]_i_220 ;
  output \rgf_c1bus_wb[11]_i_10_3 ;
  output \rgf_c1bus_wb[11]_i_10_4 ;
  output \rgf_c1bus_wb[15]_i_27 ;
  output [12:0]\grn_reg[14] ;
  output \grn_reg[15]_3 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[2]_3 ;
  output \tr_reg[15] ;
  output \tr_reg[12]_1 ;
  output \tr_reg[11]_0 ;
  output \tr_reg[10]_0 ;
  output \tr_reg[9]_0 ;
  output \tr_reg[8]_0 ;
  output \rgf_c0bus_wb[15]_i_18 ;
  output \rgf_c0bus_wb[11]_i_3 ;
  output \rgf_c0bus_wb[11]_i_3_0 ;
  output \badr[6]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_11 ;
  output \badr[5]_INST_0_i_2 ;
  output \badr[1]_INST_0_i_2 ;
  output \badr[13]_INST_0_i_2 ;
  output \badr[9]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_11_0 ;
  output \rgf_c0bus_wb[11]_i_22 ;
  output \badr[8]_INST_0_i_2 ;
  output \badr[3]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_9 ;
  output \badr[10]_INST_0_i_2 ;
  output \badr[6]_INST_0_i_2_0 ;
  output \badr[2]_INST_0_i_2 ;
  output \rgf_c0bus_wb[15]_i_25_0 ;
  output \rgf_c0bus_wb[11]_i_8 ;
  output \badr[4]_INST_0_i_2 ;
  output \rgf_c0bus_wb[0]_i_14 ;
  output \sr_reg[6]_15 ;
  output \sr_reg[6]_16 ;
  output \badr[10]_INST_0_i_2_0 ;
  output \badr[14]_INST_0_i_2 ;
  output \rgf_c0bus_wb[13]_i_29 ;
  output \badr[4]_INST_0_i_2_0 ;
  output \badr[12]_INST_0_i_2 ;
  output \badr[8]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[7]_i_7 ;
  output \rgf_c0bus_wb[7]_i_7_0 ;
  output \sr_reg[6]_17 ;
  output \sr_reg[6]_18 ;
  output \badr[14]_INST_0_i_2_0 ;
  output \sr_reg[6]_19 ;
  output \rgf_c0bus_wb[11]_i_11_1 ;
  output \rgf_c0bus_wb[11]_i_9_0 ;
  output \badr[6]_INST_0_i_2_1 ;
  output \rgf_c0bus_wb[11]_i_11_2 ;
  output \badr[13]_INST_0_i_2_0 ;
  output \badr[5]_INST_0_i_2_0 ;
  output \badr[9]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[15]_i_26 ;
  output \sr_reg[6]_20 ;
  output \badr[3]_INST_0_i_2_0 ;
  output \badr[11]_INST_0_i_2 ;
  output \badr[7]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_22_0 ;
  output \badr[2]_INST_0_i_2_0 ;
  output \sr_reg[6]_21 ;
  output \rgf_c0bus_wb[12]_i_24 ;
  output \rgf_c0bus_wb[12]_i_22_0 ;
  output \sr_reg[14] ;
  output \sr_reg[6]_22 ;
  output \sr_reg[6]_23 ;
  output \rgf_c0bus_wb[10]_i_8 ;
  output \rgf_c0bus_wb[11]_i_9_1 ;
  output \badr[1]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[13]_i_28 ;
  output \badr[14]_INST_0_i_2_1 ;
  output \rgf_c0bus_wb[8]_i_6_0 ;
  output \rgf_c0bus_wb[12]_i_25_0 ;
  output \sr_reg[6]_24 ;
  output \sr_reg[6]_25 ;
  output \sr_reg[6]_26 ;
  output \badr[8]_INST_0_i_2_1 ;
  output \badr[12]_INST_0_i_2_0 ;
  output \sr_reg[6]_27 ;
  output \sr_reg[15] ;
  output \rgf_c0bus_wb[11]_i_3_1 ;
  output \rgf_c1bus_wb[7]_i_4_0 ;
  output \sr_reg[6]_28 ;
  output \rgf_c1bus_wb[11]_i_10_5 ;
  output \rgf_c0bus_wb[15]_i_6 ;
  output \rgf_c0bus_wb[15]_i_6_0 ;
  output \rgf_c0bus_wb[15]_i_6_1 ;
  output [0:0]bbus_o;
  output \rgf_c0bus_wb[11]_i_3_2 ;
  output \rgf_c0bus_wb[11]_i_9_2 ;
  output \rgf_c0bus_wb[11]_i_9_3 ;
  output \rgf_c0bus_wb[11]_i_9_4 ;
  output \rgf_c0bus_wb[11]_i_3_3 ;
  output [3:0]\badr[14]_INST_0_i_1_1 ;
  output [2:0]\badr[13]_INST_0_i_1_0 ;
  output [0:0]\badr[14]_INST_0_i_2_2 ;
  output [1:0]\badr[6]_INST_0_i_1_3 ;
  output [1:0]tout__1_carry__0_i_1__0_0;
  output [3:0]\badr[10]_INST_0_i_1_2 ;
  output [3:0]tout__1_carry__1_i_1__0_0;
  output [14:0]p_1_in;
  output \grn_reg[15]_4 ;
  output \grn_reg[15]_5 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13] ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12] ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11] ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10] ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9] ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8] ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7] ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6] ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3] ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2] ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1] ;
  output \grn_reg[1]_0 ;
  output [0:0]\grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[0]_1 ;
  output [4:0]\grn_reg[4]_3 ;
  output [15:0]p_1_in1_in;
  output \grn_reg[15]_6 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_8 ;
  output [14:0]p_0_in;
  output \grn_reg[15]_9 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output [0:0]\grn_reg[0]_4 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_6 ;
  output [4:0]\grn_reg[4]_8 ;
  output [15:0]p_0_in0_in;
  output \grn_reg[15]_11 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_7 ;
  output \grn_reg[15]_12 ;
  output gr6_bus1;
  output \grn_reg[14]_7 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_8 ;
  output \grn_reg[15]_13 ;
  output [4:0]b1bus_b02;
  input \bdatw[13] ;
  input \bdatw[13]_0 ;
  input \bdatw[13]_1 ;
  input \bdatw[14] ;
  input \bdatw[14]_0 ;
  input \bdatw[14]_1 ;
  input \bdatw[14]_2 ;
  input \bdatw[13]_2 ;
  input \bdatw[13]_3 ;
  input \bdatw[13]_4 ;
  input \bdatw[13]_5 ;
  input \bdatw[12] ;
  input \bdatw[12]_0 ;
  input \bdatw[12]_1 ;
  input \bdatw[12]_2 ;
  input \bdatw[11] ;
  input \bdatw[11]_0 ;
  input \bdatw[11]_1 ;
  input \bdatw[11]_2 ;
  input \bdatw[10] ;
  input \bdatw[10]_0 ;
  input \bdatw[10]_1 ;
  input \bdatw[10]_2 ;
  input \bdatw[9] ;
  input \bdatw[9]_0 ;
  input \bdatw[9]_1 ;
  input \bdatw[9]_2 ;
  input \bdatw[8] ;
  input \bdatw[8]_0 ;
  input \bdatw[8]_1 ;
  input \bdatw[8]_2 ;
  input \rgf_c1bus_wb[15]_i_19 ;
  input \rgf_c1bus_wb[15]_i_19_0 ;
  input \rgf_c1bus_wb[15]_i_19_1 ;
  input \rgf_c1bus_wb[15]_i_19_2 ;
  input \sr[4]_i_77 ;
  input \rgf_c1bus_wb_reg[5] ;
  input \sr[6]_i_15 ;
  input \sr[6]_i_11 ;
  input \rgf_c1bus_wb[5]_i_10 ;
  input \rgf_c1bus_wb[14]_i_11 ;
  input \rgf_c1bus_wb[14]_i_11_0 ;
  input \rgf_c1bus_wb[14]_i_11_1 ;
  input \rgf_c1bus_wb[14]_i_11_2 ;
  input \sr[6]_i_11_0 ;
  input \sr[4]_i_77_0 ;
  input tout__1_carry__0_i_7__0;
  input tout__1_carry__0_i_7__0_0;
  input tout__1_carry__0_i_7__0_1;
  input tout__1_carry__0_i_7__0_2;
  input \rgf_c1bus_wb_reg[5]_0 ;
  input \rgf_c1bus_wb_reg[5]_1 ;
  input \rgf_c1bus_wb_reg[7] ;
  input \sr[6]_i_11_1 ;
  input \sr[6]_i_11_2 ;
  input \sr[4]_i_77_1 ;
  input \sr[6]_i_11_3 ;
  input \sr[6]_i_11_4 ;
  input \sr[6]_i_11_5 ;
  input \sr[6]_i_11_6 ;
  input \sr[4]_i_30 ;
  input [2:0]\sr[6]_i_11_7 ;
  input \sr[4]_i_30_0 ;
  input \sr[4]_i_102 ;
  input \sr[4]_i_77_2 ;
  input \rgf_c1bus_wb_reg[3] ;
  input \sr[6]_i_11_8 ;
  input \sr[6]_i_11_9 ;
  input \sr[4]_i_99 ;
  input \sr[4]_i_99_0 ;
  input \sr[4]_i_99_1 ;
  input \sr[4]_i_99_2 ;
  input \sr[4]_i_38 ;
  input \rgf_c1bus_wb_reg[4] ;
  input \sr[4]_i_119 ;
  input \rgf_c1bus_wb[12]_i_2 ;
  input \sr[4]_i_88 ;
  input \sr[4]_i_88_0 ;
  input \sr[4]_i_44 ;
  input \rgf_c1bus_wb_reg[10] ;
  input \sr[4]_i_102_0 ;
  input \sr[4]_i_111 ;
  input \sr[4]_i_84 ;
  input \sr[4]_i_177 ;
  input \sr[4]_i_177_0 ;
  input \sr[4]_i_177_1 ;
  input \sr[4]_i_177_2 ;
  input \sr[4]_i_171 ;
  input \sr[4]_i_171_0 ;
  input \sr[4]_i_171_1 ;
  input \sr[4]_i_171_2 ;
  input \sr[4]_i_169_0 ;
  input \sr[4]_i_169_1 ;
  input \sr[4]_i_169_2 ;
  input \sr[4]_i_179_0 ;
  input \sr[4]_i_169_3 ;
  input \sr[4]_i_169_4 ;
  input \sr[4]_i_169_5 ;
  input \sr[4]_i_169_6 ;
  input \sr[4]_i_175_0 ;
  input \sr[4]_i_179_1 ;
  input \sr[4]_i_175_1 ;
  input \sr[4]_i_175_2 ;
  input \sr[4]_i_169_7 ;
  input \sr[4]_i_179_2 ;
  input \sr[4]_i_169_8 ;
  input \sr[4]_i_179_3 ;
  input \sr[4]_i_175_3 ;
  input \sr[4]_i_175_4 ;
  input \sr[4]_i_175_5 ;
  input \sr[4]_i_175_6 ;
  input \sr[4]_i_179_4 ;
  input \sr[4]_i_179_5 ;
  input \sr[4]_i_179_6 ;
  input \sr[4]_i_179_7 ;
  input \rgf_c1bus_wb[4]_i_7 ;
  input \rgf_c1bus_wb[4]_i_7_0 ;
  input \rgf_c1bus_wb[4]_i_7_1 ;
  input \bdatw[15] ;
  input \bdatw[15]_0 ;
  input \bdatw[15]_1 ;
  input \bdatw[15]_2 ;
  input \bdatw[14]_3 ;
  input \bdatw[14]_4 ;
  input \bdatw[14]_5 ;
  input \bdatw[14]_6 ;
  input \bdatw[13]_6 ;
  input \bdatw[13]_7 ;
  input \bdatw[13]_8 ;
  input \bdatw[13]_9 ;
  input \bdatw[12]_3 ;
  input \bdatw[12]_4 ;
  input \bdatw[12]_5 ;
  input \bdatw[12]_6 ;
  input \bdatw[11]_3 ;
  input \bdatw[11]_4 ;
  input \bdatw[11]_5 ;
  input \bdatw[11]_6 ;
  input \bdatw[10]_3 ;
  input \bdatw[10]_4 ;
  input \bdatw[10]_5 ;
  input \bdatw[10]_6 ;
  input \bdatw[9]_3 ;
  input \bdatw[9]_4 ;
  input \bdatw[9]_5 ;
  input \bdatw[9]_6 ;
  input \bdatw[8]_3 ;
  input \bdatw[8]_4 ;
  input \bdatw[8]_5 ;
  input \bdatw[8]_6 ;
  input \rgf_c0bus_wb_reg[7]_i_11 ;
  input \sr[4]_i_67 ;
  input \rgf_c0bus_wb[6]_i_11 ;
  input \rgf_c0bus_wb[14]_i_13 ;
  input \rgf_c0bus_wb[3]_i_7 ;
  input \rgf_c0bus_wb[14]_i_13_0 ;
  input \rgf_c0bus_wb[14]_i_2 ;
  input \bbus_o[7] ;
  input \bbus_o[7]_0 ;
  input \bbus_o[7]_1 ;
  input \bbus_o[7]_2 ;
  input \rgf_c0bus_wb[3]_i_18 ;
  input \bbus_o[6] ;
  input \bbus_o[6]_0 ;
  input \bbus_o[6]_1 ;
  input \bbus_o[6]_2 ;
  input \bbus_o[5] ;
  input \bbus_o[5]_0 ;
  input \bbus_o[5]_1 ;
  input \bbus_o[5]_2 ;
  input \rgf_c0bus_wb_reg[10] ;
  input \rgf_c0bus_wb_reg[10]_0 ;
  input \rgf_c0bus_wb[12]_i_2 ;
  input \sr[4]_i_55 ;
  input \rgf_c0bus_wb[13]_i_4 ;
  input \rgf_c0bus_wb[10]_i_4 ;
  input \rgf_c0bus_wb_reg[10]_1 ;
  input \rgf_c0bus_wb[14]_i_13_1 ;
  input \rgf_c0bus_wb[14]_i_13_2 ;
  input \rgf_c0bus_wb[3]_i_7_0 ;
  input \rgf_c0bus_wb[3]_i_7_1 ;
  input \rgf_c0bus_wb[14]_i_13_3 ;
  input \rgf_c0bus_wb[14]_i_13_4 ;
  input \rgf_c0bus_wb[14]_i_13_5 ;
  input \rgf_c0bus_wb[12]_i_10 ;
  input \rgf_c0bus_wb[14]_i_13_6 ;
  input \rgf_c0bus_wb[3]_i_7_2 ;
  input \rgf_c0bus_wb[3]_i_7_3 ;
  input \rgf_c0bus_wb[3]_i_7_4 ;
  input \rgf_c0bus_wb[3]_i_18_0 ;
  input \rgf_c0bus_wb[8]_i_2 ;
  input \sr[4]_i_139 ;
  input \rgf_c0bus_wb[12]_i_7 ;
  input \sr[4]_i_126 ;
  input \rgf_c0bus_wb[15]_i_14 ;
  input \sr[4]_i_203_0 ;
  input \sr[4]_i_203_1 ;
  input \sr[4]_i_203_2 ;
  input \sr[4]_i_203_3 ;
  input \sr[4]_i_203_4 ;
  input \rgf_c0bus_wb[4]_i_7 ;
  input \sr[4]_i_188 ;
  input \sr[4]_i_188_0 ;
  input \sr[4]_i_188_1 ;
  input \sr[4]_i_188_2 ;
  input \sr[4]_i_196_0 ;
  input \sr[4]_i_196_1 ;
  input \sr[4]_i_196_2 ;
  input \sr[4]_i_196_3 ;
  input \sr[4]_i_196_4 ;
  input \sr[4]_i_196_5 ;
  input \sr[4]_i_196_6 ;
  input \sr[4]_i_196_7 ;
  input \sr[4]_i_196_8 ;
  input \sr[4]_i_196_9 ;
  input \rgf_c0bus_wb[4]_i_7_0 ;
  input \rgf_c0bus_wb[4]_i_7_1 ;
  input \rgf_c0bus_wb[4]_i_7_2 ;
  input \rgf_c0bus_wb[4]_i_7_3 ;
  input \bbus_o[5]_3 ;
  input \rgf_c0bus_wb[4]_i_3 ;
  input tout__1_carry__2;
  input tout__1_carry__2_0;
  input tout__1_carry__2_1;
  input [3:0]a0bus_sel_0;
  input [0:0]bank_sel;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_43 ;
  input [0:0]ctl_sela0;
  input \i_/badr[15]_INST_0_i_43_0 ;
  input \bbus_o[4]_INST_0_i_1 ;
  input \bbus_o[3]_INST_0_i_1 ;
  input \bbus_o[2]_INST_0_i_1 ;
  input \bbus_o[1]_INST_0_i_1 ;
  input \bbus_o[0]_INST_0_i_1 ;
  input \i_/bdatw[15]_INST_0_i_9 ;
  input \i_/bdatw[15]_INST_0_i_9_0 ;
  input \i_/bdatw[15]_INST_0_i_9_1 ;
  input \i_/bdatw[15]_INST_0_i_9_2 ;
  input [0:0]ctl_selb0_0;
  input \i_/bdatw[15]_INST_0_i_24 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_77 ;
  input [1:0]b0bus_sel_0;
  input \i_/bdatw[15]_INST_0_i_9_3 ;
  input \i_/bdatw[15]_INST_0_i_24_0 ;
  input \rgf_c1bus_wb[4]_i_22 ;
  input \rgf_c1bus_wb[4]_i_23 ;
  input \sr[4]_i_209 ;
  input \rgf_c1bus_wb[4]_i_24 ;
  input \sr[4]_i_207 ;
  input \rgf_c1bus_wb[4]_i_28 ;
  input \sr[4]_i_208 ;
  input \rgf_c1bus_wb[4]_i_27 ;
  input \sr[4]_i_225_0 ;
  input \rgf_c1bus_wb[4]_i_26 ;
  input \sr[4]_i_224_0 ;
  input \rgf_c1bus_wb[4]_i_25 ;
  input \sr[4]_i_220_0 ;
  input \sr[4]_i_211 ;
  input \sr[4]_i_213 ;
  input \sr[4]_i_210 ;
  input \i_/badr[15]_INST_0_i_19 ;
  input \i_/badr[15]_INST_0_i_19_0 ;
  input \i_/badr[15]_INST_0_i_19_1 ;
  input [2:0]a1bus_sel_0;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_113 ;
  input \i_/bdatw[15]_INST_0_i_44 ;
  input \i_/bdatw[15]_INST_0_i_112 ;
  input \i_/bdatw[15]_INST_0_i_112_0 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_112_1 ;
  input \i_/badr[15]_INST_0_i_47 ;
  input \bbus_o[4]_INST_0_i_1_0 ;
  input \bbus_o[3]_INST_0_i_1_0 ;
  input \bbus_o[2]_INST_0_i_1_0 ;
  input \bbus_o[1]_INST_0_i_1_0 ;
  input \bbus_o[0]_INST_0_i_1_0 ;
  input \rgf_c1bus_wb[4]_i_22_0 ;
  input \rgf_c1bus_wb[4]_i_23_0 ;
  input \sr[4]_i_209_0 ;
  input \rgf_c1bus_wb[4]_i_24_0 ;
  input \sr[4]_i_207_0 ;
  input \rgf_c1bus_wb[4]_i_28_0 ;
  input \sr[4]_i_208_0 ;
  input \rgf_c1bus_wb[4]_i_27_0 ;
  input \sr[4]_i_225_1 ;
  input \rgf_c1bus_wb[4]_i_26_0 ;
  input \sr[4]_i_224_1 ;
  input \rgf_c1bus_wb[4]_i_25_0 ;
  input \sr[4]_i_220_1 ;
  input \sr[4]_i_211_0 ;
  input \sr[4]_i_213_0 ;
  input \sr[4]_i_210_0 ;
  input \rgf_c1bus_wb[4]_i_47 ;
  input \rgf_c1bus_wb[4]_i_47_0 ;
  input \rgf_c1bus_wb[4]_i_41 ;
  input \rgf_c1bus_wb[4]_i_41_0 ;
  input \rgf_c1bus_wb[4]_i_51 ;
  input \rgf_c1bus_wb[4]_i_51_0 ;
  input \sr[4]_i_235 ;
  input \sr[4]_i_235_0 ;
  input \rgf_c1bus_wb[4]_i_65 ;
  input \rgf_c1bus_wb[4]_i_65_0 ;
  input \sr[4]_i_237 ;
  input \sr[4]_i_237_0 ;
  input \rgf_c1bus_wb[4]_i_61 ;
  input \rgf_c1bus_wb[4]_i_61_0 ;
  input \rgf_c1bus_wb[4]_i_57 ;
  input \rgf_c1bus_wb[4]_i_57_0 ;
  input \sr[4]_i_245 ;
  input \sr[4]_i_245_0 ;
  input \rgf_c1bus_wb[4]_i_53 ;
  input \rgf_c1bus_wb[4]_i_53_0 ;
  input \sr[4]_i_243 ;
  input \sr[4]_i_243_0 ;
  input \rgf_c1bus_wb[4]_i_33 ;
  input \rgf_c1bus_wb[4]_i_33_0 ;
  input \rgf_c1bus_wb[4]_i_67 ;
  input \rgf_c1bus_wb[4]_i_67_0 ;
  input \rgf_c1bus_wb[4]_i_37 ;
  input \rgf_c1bus_wb[4]_i_37_0 ;
  input \sr[4]_i_240 ;
  input \sr[4]_i_240_0 ;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_14 ;
  input [15:0]\grn_reg[15]_15 ;
  input clk;
  input [0:0]\grn_reg[15]_16 ;
  input [15:0]\grn_reg[15]_17 ;
  input [0:0]\grn_reg[15]_18 ;
  input [15:0]\grn_reg[15]_19 ;
  input [0:0]\grn_reg[15]_20 ;
  input [15:0]\grn_reg[15]_21 ;
  input [0:0]\grn_reg[15]_22 ;
  input [15:0]\grn_reg[15]_23 ;
  input [0:0]\grn_reg[15]_24 ;
  input [15:0]\grn_reg[15]_25 ;
  input [0:0]\grn_reg[15]_26 ;
  input [15:0]\grn_reg[15]_27 ;
  input [0:0]\grn_reg[15]_28 ;
  input [15:0]\grn_reg[15]_29 ;
  input [0:0]\grn_reg[15]_30 ;
  input [15:0]\grn_reg[15]_31 ;
  input [0:0]\grn_reg[15]_32 ;
  input [15:0]\grn_reg[15]_33 ;
  input [0:0]\grn_reg[15]_34 ;
  input [15:0]\grn_reg[15]_35 ;
  input [0:0]\grn_reg[15]_36 ;
  input [15:0]\grn_reg[15]_37 ;
  input [0:0]\grn_reg[15]_38 ;
  input [15:0]\grn_reg[15]_39 ;
  input [0:0]\grn_reg[15]_40 ;
  input [15:0]\grn_reg[15]_41 ;
  input [0:0]\grn_reg[15]_42 ;
  input [15:0]\grn_reg[15]_43 ;
  input [0:0]\grn_reg[15]_44 ;
  input [15:0]\grn_reg[15]_45 ;
     output [15:0]gr20;
     output [15:0]gr21;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr01;
     output [15:0]gr05;
     output [15:0]gr06;

  wire [0:0]SR;
  wire [3:0]a0bus_sel_0;
  wire [7:5]a1bus_b02;
  wire [2:0]a1bus_sel_0;
  wire a1buso2l_n_23;
  wire a1buso2l_n_34;
  wire a1buso2l_n_36;
  wire a1buso2l_n_38;
  wire a1buso2l_n_40;
  wire a1buso2l_n_42;
  wire a1buso2l_n_44;
  wire a1buso2l_n_46;
  wire a1buso2l_n_47;
  wire a1buso2l_n_49;
  wire a1buso2l_n_51;
  wire a1buso2l_n_53;
  wire a1buso2l_n_55;
  wire a1buso2l_n_57;
  wire a1buso2l_n_59;
  wire a1buso2l_n_61;
  wire a1buso2l_n_63;
  wire a1buso_n_30;
  wire a1buso_n_31;
  wire [1:0]b0bus_sel_0;
  wire [4:0]b1bus_b02;
  wire b1buso2l_n_1;
  wire b1buso2l_n_10;
  wire b1buso2l_n_11;
  wire b1buso2l_n_12;
  wire b1buso2l_n_13;
  wire b1buso2l_n_14;
  wire b1buso2l_n_15;
  wire b1buso2l_n_16;
  wire b1buso2l_n_17;
  wire b1buso2l_n_18;
  wire b1buso2l_n_19;
  wire b1buso2l_n_2;
  wire b1buso2l_n_20;
  wire b1buso2l_n_21;
  wire b1buso2l_n_22;
  wire b1buso2l_n_23;
  wire b1buso2l_n_24;
  wire b1buso2l_n_25;
  wire b1buso2l_n_3;
  wire b1buso2l_n_4;
  wire b1buso2l_n_5;
  wire b1buso2l_n_6;
  wire b1buso2l_n_7;
  wire b1buso2l_n_8;
  wire b1buso2l_n_9;
  wire b1buso_n_1;
  wire b1buso_n_10;
  wire b1buso_n_11;
  wire b1buso_n_12;
  wire b1buso_n_13;
  wire b1buso_n_14;
  wire b1buso_n_15;
  wire b1buso_n_16;
  wire b1buso_n_17;
  wire b1buso_n_18;
  wire b1buso_n_19;
  wire b1buso_n_2;
  wire b1buso_n_20;
  wire b1buso_n_21;
  wire b1buso_n_22;
  wire b1buso_n_23;
  wire b1buso_n_24;
  wire b1buso_n_25;
  wire b1buso_n_3;
  wire b1buso_n_4;
  wire b1buso_n_5;
  wire b1buso_n_6;
  wire b1buso_n_7;
  wire b1buso_n_8;
  wire b1buso_n_9;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1_0 ;
  wire \badr[10]_INST_0_i_1_1 ;
  wire [3:0]\badr[10]_INST_0_i_1_2 ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[10]_INST_0_i_2_0 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2_0 ;
  wire \badr[13]_INST_0_i_1 ;
  wire [2:0]\badr[13]_INST_0_i_1_0 ;
  wire \badr[13]_INST_0_i_2 ;
  wire \badr[13]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire [3:0]\badr[14]_INST_0_i_1_1 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_2_1 ;
  wire [0:0]\badr[14]_INST_0_i_2_2 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_1_1 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2_0 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1_0 ;
  wire \badr[2]_INST_0_i_1_1 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[2]_INST_0_i_2_0 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1_0 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[3]_INST_0_i_2_0 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_2_0 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_2_0 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1_0 ;
  wire \badr[6]_INST_0_i_1_1 ;
  wire \badr[6]_INST_0_i_1_2 ;
  wire [1:0]\badr[6]_INST_0_i_1_3 ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2_0 ;
  wire \badr[6]_INST_0_i_2_1 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2_0 ;
  wire \badr[8]_INST_0_i_2_1 ;
  wire \badr[9]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1_0 ;
  wire \badr[9]_INST_0_i_2 ;
  wire \badr[9]_INST_0_i_2_0 ;
  wire [0:0]bank_sel;
  wire [0:0]bbus_o;
  wire \bbus_o[0]_INST_0_i_1 ;
  wire \bbus_o[0]_INST_0_i_1_0 ;
  wire \bbus_o[1]_INST_0_i_1 ;
  wire \bbus_o[1]_INST_0_i_1_0 ;
  wire \bbus_o[2]_INST_0_i_1 ;
  wire \bbus_o[2]_INST_0_i_1_0 ;
  wire \bbus_o[3]_INST_0_i_1 ;
  wire \bbus_o[3]_INST_0_i_1_0 ;
  wire \bbus_o[4]_INST_0_i_1 ;
  wire \bbus_o[4]_INST_0_i_1_0 ;
  wire \bbus_o[5] ;
  wire \bbus_o[5]_0 ;
  wire \bbus_o[5]_1 ;
  wire \bbus_o[5]_2 ;
  wire \bbus_o[5]_3 ;
  wire \bbus_o[6] ;
  wire \bbus_o[6]_0 ;
  wire \bbus_o[6]_1 ;
  wire \bbus_o[6]_2 ;
  wire \bbus_o[7] ;
  wire \bbus_o[7]_0 ;
  wire \bbus_o[7]_1 ;
  wire \bbus_o[7]_2 ;
  wire [1:0]bdatw;
  wire \bdatw[10] ;
  wire \bdatw[10]_0 ;
  wire \bdatw[10]_1 ;
  wire \bdatw[10]_2 ;
  wire \bdatw[10]_3 ;
  wire \bdatw[10]_4 ;
  wire \bdatw[10]_5 ;
  wire \bdatw[10]_6 ;
  wire \bdatw[11] ;
  wire \bdatw[11]_0 ;
  wire \bdatw[11]_1 ;
  wire \bdatw[11]_2 ;
  wire \bdatw[11]_3 ;
  wire \bdatw[11]_4 ;
  wire \bdatw[11]_5 ;
  wire \bdatw[11]_6 ;
  wire \bdatw[12] ;
  wire \bdatw[12]_0 ;
  wire \bdatw[12]_1 ;
  wire \bdatw[12]_2 ;
  wire \bdatw[12]_3 ;
  wire \bdatw[12]_4 ;
  wire \bdatw[12]_5 ;
  wire \bdatw[12]_6 ;
  wire \bdatw[13] ;
  wire \bdatw[13]_0 ;
  wire \bdatw[13]_1 ;
  wire \bdatw[13]_2 ;
  wire \bdatw[13]_3 ;
  wire \bdatw[13]_4 ;
  wire \bdatw[13]_5 ;
  wire \bdatw[13]_6 ;
  wire \bdatw[13]_7 ;
  wire \bdatw[13]_8 ;
  wire \bdatw[13]_9 ;
  wire \bdatw[14] ;
  wire \bdatw[14]_0 ;
  wire \bdatw[14]_1 ;
  wire \bdatw[14]_2 ;
  wire \bdatw[14]_3 ;
  wire \bdatw[14]_4 ;
  wire \bdatw[14]_5 ;
  wire \bdatw[14]_6 ;
  wire \bdatw[15] ;
  wire \bdatw[15]_0 ;
  wire \bdatw[15]_1 ;
  wire \bdatw[15]_2 ;
  wire \bdatw[8] ;
  wire \bdatw[8]_0 ;
  wire \bdatw[8]_1 ;
  wire \bdatw[8]_2 ;
  wire \bdatw[8]_3 ;
  wire \bdatw[8]_4 ;
  wire \bdatw[8]_5 ;
  wire \bdatw[8]_6 ;
  wire \bdatw[9] ;
  wire \bdatw[9]_0 ;
  wire \bdatw[9]_1 ;
  wire \bdatw[9]_2 ;
  wire \bdatw[9]_3 ;
  wire \bdatw[9]_4 ;
  wire \bdatw[9]_5 ;
  wire \bdatw[9]_6 ;
  wire clk;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire gr6_bus1;
  wire [0:0]\grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire [0:0]\grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire [12:0]\grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[14]_7 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire [0:0]\grn_reg[15]_14 ;
  wire [15:0]\grn_reg[15]_15 ;
  wire [0:0]\grn_reg[15]_16 ;
  wire [15:0]\grn_reg[15]_17 ;
  wire [0:0]\grn_reg[15]_18 ;
  wire [15:0]\grn_reg[15]_19 ;
  wire [0:0]\grn_reg[15]_20 ;
  wire [15:0]\grn_reg[15]_21 ;
  wire [0:0]\grn_reg[15]_22 ;
  wire [15:0]\grn_reg[15]_23 ;
  wire [0:0]\grn_reg[15]_24 ;
  wire [15:0]\grn_reg[15]_25 ;
  wire [0:0]\grn_reg[15]_26 ;
  wire [15:0]\grn_reg[15]_27 ;
  wire [0:0]\grn_reg[15]_28 ;
  wire [15:0]\grn_reg[15]_29 ;
  wire \grn_reg[15]_3 ;
  wire [0:0]\grn_reg[15]_30 ;
  wire [15:0]\grn_reg[15]_31 ;
  wire [0:0]\grn_reg[15]_32 ;
  wire [15:0]\grn_reg[15]_33 ;
  wire [0:0]\grn_reg[15]_34 ;
  wire [15:0]\grn_reg[15]_35 ;
  wire [0:0]\grn_reg[15]_36 ;
  wire [15:0]\grn_reg[15]_37 ;
  wire [0:0]\grn_reg[15]_38 ;
  wire [15:0]\grn_reg[15]_39 ;
  wire \grn_reg[15]_4 ;
  wire [0:0]\grn_reg[15]_40 ;
  wire [15:0]\grn_reg[15]_41 ;
  wire [0:0]\grn_reg[15]_42 ;
  wire [15:0]\grn_reg[15]_43 ;
  wire [0:0]\grn_reg[15]_44 ;
  wire [15:0]\grn_reg[15]_45 ;
  wire \grn_reg[15]_5 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_2 ;
  wire [4:0]\grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire [4:0]\grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire \i_/badr[15]_INST_0_i_19 ;
  wire \i_/badr[15]_INST_0_i_19_0 ;
  wire \i_/badr[15]_INST_0_i_19_1 ;
  wire \i_/badr[15]_INST_0_i_43 ;
  wire \i_/badr[15]_INST_0_i_43_0 ;
  wire \i_/badr[15]_INST_0_i_47 ;
  wire \i_/bdatw[15]_INST_0_i_112 ;
  wire \i_/bdatw[15]_INST_0_i_112_0 ;
  wire \i_/bdatw[15]_INST_0_i_112_1 ;
  wire \i_/bdatw[15]_INST_0_i_113 ;
  wire \i_/bdatw[15]_INST_0_i_24 ;
  wire \i_/bdatw[15]_INST_0_i_24_0 ;
  wire \i_/bdatw[15]_INST_0_i_44 ;
  wire \i_/bdatw[15]_INST_0_i_77 ;
  wire \i_/bdatw[15]_INST_0_i_9 ;
  wire \i_/bdatw[15]_INST_0_i_9_0 ;
  wire \i_/bdatw[15]_INST_0_i_9_1 ;
  wire \i_/bdatw[15]_INST_0_i_9_2 ;
  wire \i_/bdatw[15]_INST_0_i_9_3 ;
  wire [14:0]p_0_in;
  wire [15:0]p_0_in0_in;
  wire [15:5]p_0_in2_in;
  wire [14:0]p_1_in;
  wire [15:0]p_1_in1_in;
  wire [15:5]p_1_in3_in;
  wire \rgf_c0bus_wb[0]_i_14 ;
  wire \rgf_c0bus_wb[10]_i_4 ;
  wire \rgf_c0bus_wb[10]_i_8 ;
  wire \rgf_c0bus_wb[11]_i_11 ;
  wire \rgf_c0bus_wb[11]_i_11_0 ;
  wire \rgf_c0bus_wb[11]_i_11_1 ;
  wire \rgf_c0bus_wb[11]_i_11_2 ;
  wire \rgf_c0bus_wb[11]_i_22 ;
  wire \rgf_c0bus_wb[11]_i_22_0 ;
  wire \rgf_c0bus_wb[11]_i_3 ;
  wire \rgf_c0bus_wb[11]_i_3_0 ;
  wire \rgf_c0bus_wb[11]_i_3_1 ;
  wire \rgf_c0bus_wb[11]_i_3_2 ;
  wire \rgf_c0bus_wb[11]_i_3_3 ;
  wire \rgf_c0bus_wb[11]_i_8 ;
  wire \rgf_c0bus_wb[11]_i_9 ;
  wire \rgf_c0bus_wb[11]_i_9_0 ;
  wire \rgf_c0bus_wb[11]_i_9_1 ;
  wire \rgf_c0bus_wb[11]_i_9_2 ;
  wire \rgf_c0bus_wb[11]_i_9_3 ;
  wire \rgf_c0bus_wb[11]_i_9_4 ;
  wire \rgf_c0bus_wb[12]_i_10 ;
  wire \rgf_c0bus_wb[12]_i_2 ;
  wire \rgf_c0bus_wb[12]_i_22_0 ;
  wire \rgf_c0bus_wb[12]_i_22_n_0 ;
  wire \rgf_c0bus_wb[12]_i_23_n_0 ;
  wire \rgf_c0bus_wb[12]_i_24 ;
  wire \rgf_c0bus_wb[12]_i_25_0 ;
  wire \rgf_c0bus_wb[12]_i_25_n_0 ;
  wire \rgf_c0bus_wb[12]_i_7 ;
  wire \rgf_c0bus_wb[13]_i_28 ;
  wire \rgf_c0bus_wb[13]_i_29 ;
  wire \rgf_c0bus_wb[13]_i_4 ;
  wire \rgf_c0bus_wb[14]_i_13 ;
  wire \rgf_c0bus_wb[14]_i_13_0 ;
  wire \rgf_c0bus_wb[14]_i_13_1 ;
  wire \rgf_c0bus_wb[14]_i_13_2 ;
  wire \rgf_c0bus_wb[14]_i_13_3 ;
  wire \rgf_c0bus_wb[14]_i_13_4 ;
  wire \rgf_c0bus_wb[14]_i_13_5 ;
  wire \rgf_c0bus_wb[14]_i_13_6 ;
  wire \rgf_c0bus_wb[14]_i_2 ;
  wire \rgf_c0bus_wb[15]_i_14 ;
  wire \rgf_c0bus_wb[15]_i_18 ;
  wire \rgf_c0bus_wb[15]_i_25_0 ;
  wire \rgf_c0bus_wb[15]_i_26 ;
  wire \rgf_c0bus_wb[15]_i_6 ;
  wire \rgf_c0bus_wb[15]_i_6_0 ;
  wire \rgf_c0bus_wb[15]_i_6_1 ;
  wire \rgf_c0bus_wb[3]_i_18 ;
  wire \rgf_c0bus_wb[3]_i_18_0 ;
  wire \rgf_c0bus_wb[3]_i_7 ;
  wire \rgf_c0bus_wb[3]_i_7_0 ;
  wire \rgf_c0bus_wb[3]_i_7_1 ;
  wire \rgf_c0bus_wb[3]_i_7_2 ;
  wire \rgf_c0bus_wb[3]_i_7_3 ;
  wire \rgf_c0bus_wb[3]_i_7_4 ;
  wire \rgf_c0bus_wb[4]_i_3 ;
  wire \rgf_c0bus_wb[4]_i_7 ;
  wire \rgf_c0bus_wb[4]_i_7_0 ;
  wire \rgf_c0bus_wb[4]_i_7_1 ;
  wire \rgf_c0bus_wb[4]_i_7_2 ;
  wire \rgf_c0bus_wb[4]_i_7_3 ;
  wire \rgf_c0bus_wb[6]_i_11 ;
  wire \rgf_c0bus_wb[7]_i_7 ;
  wire \rgf_c0bus_wb[7]_i_7_0 ;
  wire \rgf_c0bus_wb[8]_i_2 ;
  wire \rgf_c0bus_wb[8]_i_6_0 ;
  wire \rgf_c0bus_wb_reg[10] ;
  wire \rgf_c0bus_wb_reg[10]_0 ;
  wire \rgf_c0bus_wb_reg[10]_1 ;
  wire \rgf_c0bus_wb_reg[7]_i_11 ;
  wire \rgf_c1bus_wb[11]_i_10 ;
  wire \rgf_c1bus_wb[11]_i_10_0 ;
  wire \rgf_c1bus_wb[11]_i_10_1 ;
  wire \rgf_c1bus_wb[11]_i_10_2 ;
  wire \rgf_c1bus_wb[11]_i_10_3 ;
  wire \rgf_c1bus_wb[11]_i_10_4 ;
  wire \rgf_c1bus_wb[11]_i_10_5 ;
  wire \rgf_c1bus_wb[11]_i_13 ;
  wire \rgf_c1bus_wb[12]_i_2 ;
  wire \rgf_c1bus_wb[12]_i_20_0 ;
  wire \rgf_c1bus_wb[13]_i_16 ;
  wire \rgf_c1bus_wb[13]_i_9 ;
  wire \rgf_c1bus_wb[14]_i_11 ;
  wire \rgf_c1bus_wb[14]_i_11_0 ;
  wire \rgf_c1bus_wb[14]_i_11_1 ;
  wire \rgf_c1bus_wb[14]_i_11_2 ;
  wire \rgf_c1bus_wb[14]_i_28 ;
  wire \rgf_c1bus_wb[14]_i_28_0 ;
  wire \rgf_c1bus_wb[14]_i_28_1 ;
  wire \rgf_c1bus_wb[14]_i_28_2 ;
  wire \rgf_c1bus_wb[14]_i_28_3 ;
  wire \rgf_c1bus_wb[14]_i_28_4 ;
  wire \rgf_c1bus_wb[14]_i_28_5 ;
  wire \rgf_c1bus_wb[14]_i_28_6 ;
  wire \rgf_c1bus_wb[14]_i_30 ;
  wire \rgf_c1bus_wb[14]_i_32 ;
  wire \rgf_c1bus_wb[14]_i_32_0 ;
  wire \rgf_c1bus_wb[15]_i_14 ;
  wire \rgf_c1bus_wb[15]_i_14_0 ;
  wire \rgf_c1bus_wb[15]_i_14_1 ;
  wire \rgf_c1bus_wb[15]_i_14_2 ;
  wire \rgf_c1bus_wb[15]_i_14_3 ;
  wire \rgf_c1bus_wb[15]_i_19 ;
  wire \rgf_c1bus_wb[15]_i_19_0 ;
  wire \rgf_c1bus_wb[15]_i_19_1 ;
  wire \rgf_c1bus_wb[15]_i_19_2 ;
  wire \rgf_c1bus_wb[15]_i_27 ;
  wire \rgf_c1bus_wb[1]_i_14_0 ;
  wire \rgf_c1bus_wb[4]_i_18_n_0 ;
  wire \rgf_c1bus_wb[4]_i_19_n_0 ;
  wire \rgf_c1bus_wb[4]_i_22 ;
  wire \rgf_c1bus_wb[4]_i_22_0 ;
  wire \rgf_c1bus_wb[4]_i_23 ;
  wire \rgf_c1bus_wb[4]_i_23_0 ;
  wire \rgf_c1bus_wb[4]_i_24 ;
  wire \rgf_c1bus_wb[4]_i_24_0 ;
  wire \rgf_c1bus_wb[4]_i_25 ;
  wire \rgf_c1bus_wb[4]_i_25_0 ;
  wire \rgf_c1bus_wb[4]_i_26 ;
  wire \rgf_c1bus_wb[4]_i_26_0 ;
  wire \rgf_c1bus_wb[4]_i_27 ;
  wire \rgf_c1bus_wb[4]_i_27_0 ;
  wire \rgf_c1bus_wb[4]_i_28 ;
  wire \rgf_c1bus_wb[4]_i_28_0 ;
  wire \rgf_c1bus_wb[4]_i_33 ;
  wire \rgf_c1bus_wb[4]_i_33_0 ;
  wire \rgf_c1bus_wb[4]_i_37 ;
  wire \rgf_c1bus_wb[4]_i_37_0 ;
  wire \rgf_c1bus_wb[4]_i_41 ;
  wire \rgf_c1bus_wb[4]_i_41_0 ;
  wire \rgf_c1bus_wb[4]_i_47 ;
  wire \rgf_c1bus_wb[4]_i_47_0 ;
  wire \rgf_c1bus_wb[4]_i_51 ;
  wire \rgf_c1bus_wb[4]_i_51_0 ;
  wire \rgf_c1bus_wb[4]_i_53 ;
  wire \rgf_c1bus_wb[4]_i_53_0 ;
  wire \rgf_c1bus_wb[4]_i_57 ;
  wire \rgf_c1bus_wb[4]_i_57_0 ;
  wire \rgf_c1bus_wb[4]_i_61 ;
  wire \rgf_c1bus_wb[4]_i_61_0 ;
  wire \rgf_c1bus_wb[4]_i_65 ;
  wire \rgf_c1bus_wb[4]_i_65_0 ;
  wire \rgf_c1bus_wb[4]_i_67 ;
  wire \rgf_c1bus_wb[4]_i_67_0 ;
  wire \rgf_c1bus_wb[4]_i_7 ;
  wire \rgf_c1bus_wb[4]_i_7_0 ;
  wire \rgf_c1bus_wb[4]_i_7_1 ;
  wire \rgf_c1bus_wb[4]_i_9 ;
  wire \rgf_c1bus_wb[4]_i_9_0 ;
  wire \rgf_c1bus_wb[5]_i_10 ;
  wire \rgf_c1bus_wb[7]_i_4 ;
  wire \rgf_c1bus_wb[7]_i_4_0 ;
  wire \rgf_c1bus_wb[9]_i_17_0 ;
  wire \rgf_c1bus_wb_reg[10] ;
  wire \rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[5]_0 ;
  wire \rgf_c1bus_wb_reg[5]_1 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire \sr[4]_i_102 ;
  wire \sr[4]_i_102_0 ;
  wire \sr[4]_i_111 ;
  wire \sr[4]_i_119 ;
  wire \sr[4]_i_126 ;
  wire \sr[4]_i_139 ;
  wire \sr[4]_i_169_0 ;
  wire \sr[4]_i_169_1 ;
  wire \sr[4]_i_169_2 ;
  wire \sr[4]_i_169_3 ;
  wire \sr[4]_i_169_4 ;
  wire \sr[4]_i_169_5 ;
  wire \sr[4]_i_169_6 ;
  wire \sr[4]_i_169_7 ;
  wire \sr[4]_i_169_8 ;
  wire \sr[4]_i_171 ;
  wire \sr[4]_i_171_0 ;
  wire \sr[4]_i_171_1 ;
  wire \sr[4]_i_171_2 ;
  wire \sr[4]_i_175_0 ;
  wire \sr[4]_i_175_1 ;
  wire \sr[4]_i_175_2 ;
  wire \sr[4]_i_175_3 ;
  wire \sr[4]_i_175_4 ;
  wire \sr[4]_i_175_5 ;
  wire \sr[4]_i_175_6 ;
  wire \sr[4]_i_177 ;
  wire \sr[4]_i_177_0 ;
  wire \sr[4]_i_177_1 ;
  wire \sr[4]_i_177_2 ;
  wire \sr[4]_i_179_0 ;
  wire \sr[4]_i_179_1 ;
  wire \sr[4]_i_179_2 ;
  wire \sr[4]_i_179_3 ;
  wire \sr[4]_i_179_4 ;
  wire \sr[4]_i_179_5 ;
  wire \sr[4]_i_179_6 ;
  wire \sr[4]_i_179_7 ;
  wire \sr[4]_i_188 ;
  wire \sr[4]_i_188_0 ;
  wire \sr[4]_i_188_1 ;
  wire \sr[4]_i_188_2 ;
  wire \sr[4]_i_196_0 ;
  wire \sr[4]_i_196_1 ;
  wire \sr[4]_i_196_2 ;
  wire \sr[4]_i_196_3 ;
  wire \sr[4]_i_196_4 ;
  wire \sr[4]_i_196_5 ;
  wire \sr[4]_i_196_6 ;
  wire \sr[4]_i_196_7 ;
  wire \sr[4]_i_196_8 ;
  wire \sr[4]_i_196_9 ;
  wire \sr[4]_i_203_0 ;
  wire \sr[4]_i_203_1 ;
  wire \sr[4]_i_203_2 ;
  wire \sr[4]_i_203_3 ;
  wire \sr[4]_i_203_4 ;
  wire \sr[4]_i_207 ;
  wire \sr[4]_i_207_0 ;
  wire \sr[4]_i_208 ;
  wire \sr[4]_i_208_0 ;
  wire \sr[4]_i_209 ;
  wire \sr[4]_i_209_0 ;
  wire \sr[4]_i_210 ;
  wire \sr[4]_i_210_0 ;
  wire \sr[4]_i_211 ;
  wire \sr[4]_i_211_0 ;
  wire \sr[4]_i_213 ;
  wire \sr[4]_i_213_0 ;
  wire \sr[4]_i_217_n_0 ;
  wire \sr[4]_i_218_n_0 ;
  wire \sr[4]_i_219_0 ;
  wire \sr[4]_i_219_n_0 ;
  wire \sr[4]_i_220 ;
  wire \sr[4]_i_220_0 ;
  wire \sr[4]_i_220_1 ;
  wire \sr[4]_i_224_0 ;
  wire \sr[4]_i_224_1 ;
  wire \sr[4]_i_224_n_0 ;
  wire \sr[4]_i_225_0 ;
  wire \sr[4]_i_225_1 ;
  wire \sr[4]_i_225_n_0 ;
  wire \sr[4]_i_235 ;
  wire \sr[4]_i_235_0 ;
  wire \sr[4]_i_237 ;
  wire \sr[4]_i_237_0 ;
  wire \sr[4]_i_240 ;
  wire \sr[4]_i_240_0 ;
  wire \sr[4]_i_243 ;
  wire \sr[4]_i_243_0 ;
  wire \sr[4]_i_245 ;
  wire \sr[4]_i_245_0 ;
  wire \sr[4]_i_30 ;
  wire \sr[4]_i_30_0 ;
  wire \sr[4]_i_38 ;
  wire \sr[4]_i_44 ;
  wire \sr[4]_i_55 ;
  wire \sr[4]_i_67 ;
  wire \sr[4]_i_77 ;
  wire \sr[4]_i_77_0 ;
  wire \sr[4]_i_77_1 ;
  wire \sr[4]_i_77_2 ;
  wire \sr[4]_i_84 ;
  wire \sr[4]_i_88 ;
  wire \sr[4]_i_88_0 ;
  wire \sr[4]_i_99 ;
  wire \sr[4]_i_99_0 ;
  wire \sr[4]_i_99_1 ;
  wire \sr[4]_i_99_2 ;
  wire \sr[6]_i_11 ;
  wire \sr[6]_i_11_0 ;
  wire \sr[6]_i_11_1 ;
  wire \sr[6]_i_11_2 ;
  wire \sr[6]_i_11_3 ;
  wire \sr[6]_i_11_4 ;
  wire \sr[6]_i_11_5 ;
  wire \sr[6]_i_11_6 ;
  wire [2:0]\sr[6]_i_11_7 ;
  wire \sr[6]_i_11_8 ;
  wire \sr[6]_i_11_9 ;
  wire \sr[6]_i_15 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_11 ;
  wire \sr_reg[6]_12 ;
  wire \sr_reg[6]_13 ;
  wire \sr_reg[6]_14 ;
  wire \sr_reg[6]_15 ;
  wire \sr_reg[6]_16 ;
  wire \sr_reg[6]_17 ;
  wire \sr_reg[6]_18 ;
  wire \sr_reg[6]_19 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_20 ;
  wire \sr_reg[6]_21 ;
  wire \sr_reg[6]_22 ;
  wire \sr_reg[6]_23 ;
  wire \sr_reg[6]_24 ;
  wire \sr_reg[6]_25 ;
  wire \sr_reg[6]_26 ;
  wire \sr_reg[6]_27 ;
  wire \sr_reg[6]_28 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_7 ;
  wire \sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[2] ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire [1:0]tout__1_carry__0_i_1__0_0;
  wire tout__1_carry__0_i_7__0;
  wire tout__1_carry__0_i_7__0_0;
  wire tout__1_carry__0_i_7__0_1;
  wire tout__1_carry__0_i_7__0_2;
  wire [3:0]tout__1_carry__1_i_1__0_0;
  wire tout__1_carry__2;
  wire tout__1_carry__2_0;
  wire tout__1_carry__2_1;
  wire \tr_reg[10] ;
  wire \tr_reg[10]_0 ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[12]_1 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire \tr_reg[14]_1 ;
  wire \tr_reg[15] ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[8] ;
  wire \tr_reg[8]_0 ;
  wire \tr_reg[9] ;
  wire \tr_reg[9]_0 ;

  mcss_rgf_bank_bus_28 a0buso
       (.a0bus_sel_0(a0bus_sel_0),
        .bank_sel(bank_sel),
        .ctl_sela0(ctl_sela0),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[0]_1 (\grn_reg[0]_1 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[10]_0 (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[11]_0 (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[12]_0 (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[13]_0 (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14]_0 ),
        .\grn_reg[14]_0 (\grn_reg[14]_1 ),
        .\grn_reg[15] (\grn_reg[15]_4 ),
        .\grn_reg[15]_0 (\grn_reg[15]_5 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4]_1 ),
        .\grn_reg[4]_0 (\grn_reg[4]_2 ),
        .\grn_reg[5] (\grn_reg[5] ),
        .\grn_reg[5]_0 (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[6]_0 (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[7]_0 (\grn_reg[7]_0 ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[8]_0 (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\grn_reg[9]_0 (\grn_reg[9]_0 ),
        .\i_/badr[15]_INST_0_i_10_0 (\sr[6]_i_11_7 [1:0]),
        .\i_/badr[15]_INST_0_i_10_1 (gr06),
        .\i_/badr[15]_INST_0_i_10_2 (gr05),
        .\i_/badr[15]_INST_0_i_43_0 (\i_/badr[15]_INST_0_i_43 ),
        .\i_/badr[15]_INST_0_i_43_1 (\i_/badr[15]_INST_0_i_43_0 ),
        .\i_/badr[15]_INST_0_i_46_0 (gr02),
        .\i_/badr[15]_INST_0_i_46_1 (gr01),
        .out(gr00),
        .p_1_in(p_1_in),
        .\rgf_c0bus_wb[4]_i_41 (gr07),
        .\rgf_c0bus_wb[4]_i_41_0 (gr03),
        .\rgf_c0bus_wb[4]_i_41_1 (gr04));
  mcss_rgf_bank_bus_29 a0buso2l
       (.a0bus_sel_0(a0bus_sel_0),
        .ctl_sela0(ctl_sela0),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (\grn_reg[0]_4 ),
        .\grn_reg[0]_0 (\grn_reg[0]_5 ),
        .\grn_reg[0]_1 (\grn_reg[0]_6 ),
        .\grn_reg[10] (\grn_reg[10]_3 ),
        .\grn_reg[10]_0 (\grn_reg[10]_4 ),
        .\grn_reg[11] (\grn_reg[11]_3 ),
        .\grn_reg[11]_0 (\grn_reg[11]_4 ),
        .\grn_reg[12] (\grn_reg[12]_3 ),
        .\grn_reg[12]_0 (\grn_reg[12]_4 ),
        .\grn_reg[13] (\grn_reg[13]_3 ),
        .\grn_reg[13]_0 (\grn_reg[13]_4 ),
        .\grn_reg[14] (\grn_reg[14]_4 ),
        .\grn_reg[14]_0 (\grn_reg[14]_5 ),
        .\grn_reg[15] (\grn_reg[15]_9 ),
        .\grn_reg[15]_0 (\grn_reg[15]_10 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[1]_0 (\grn_reg[1]_4 ),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[2]_0 (\grn_reg[2]_4 ),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[4] (\grn_reg[4]_6 ),
        .\grn_reg[4]_0 (\grn_reg[4]_7 ),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\grn_reg[6] (\grn_reg[6]_3 ),
        .\grn_reg[6]_0 (\grn_reg[6]_4 ),
        .\grn_reg[7] (\grn_reg[7]_3 ),
        .\grn_reg[7]_0 (\grn_reg[7]_4 ),
        .\grn_reg[8] (\grn_reg[8]_1 ),
        .\grn_reg[8]_0 (\grn_reg[8]_2 ),
        .\grn_reg[9] (\grn_reg[9]_3 ),
        .\grn_reg[9]_0 (\grn_reg[9]_4 ),
        .\i_/badr[15]_INST_0_i_11_0 (gr26),
        .\i_/badr[15]_INST_0_i_11_1 (gr25),
        .\i_/badr[15]_INST_0_i_47_0 (\i_/badr[15]_INST_0_i_47 ),
        .\i_/badr[15]_INST_0_i_47_1 (\i_/badr[15]_INST_0_i_43 ),
        .\i_/badr[15]_INST_0_i_47_2 (\i_/badr[15]_INST_0_i_43_0 ),
        .\i_/badr[15]_INST_0_i_50_0 (\sr[6]_i_11_7 [1:0]),
        .\i_/badr[15]_INST_0_i_50_1 (gr22),
        .\i_/badr[15]_INST_0_i_50_2 (gr21),
        .out(gr20),
        .p_0_in(p_0_in),
        .\rgf_c0bus_wb[4]_i_41 (gr27),
        .\rgf_c0bus_wb[4]_i_41_0 (gr23),
        .\rgf_c0bus_wb[4]_i_41_1 (gr24));
  mcss_rgf_bank_bus_30 a1buso
       (.a1bus_sel_0({a1bus_sel_0[2],a1bus_sel_0[0]}),
        .\badr[0]_INST_0_i_1 (\sr[4]_i_210 ),
        .\badr[10]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_28 ),
        .\badr[11]_INST_0_i_1 (\sr[4]_i_207 ),
        .\badr[12]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_24 ),
        .\badr[13]_INST_0_i_1 (\sr[4]_i_209 ),
        .\badr[14]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_23 ),
        .\badr[15]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_22 ),
        .\badr[1]_INST_0_i_1 (\sr[4]_i_213 ),
        .\badr[2]_INST_0_i_1 (\sr[4]_i_211 ),
        .\badr[3]_INST_0_i_1 (\sr[4]_i_220_0 ),
        .\badr[4]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_25 ),
        .\badr[5]_INST_0_i_1 (\sr[4]_i_224_0 ),
        .\badr[6]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_26 ),
        .\badr[7]_INST_0_i_1 (\sr[4]_i_225_0 ),
        .\badr[8]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_27 ),
        .\badr[9]_INST_0_i_1 (\sr[4]_i_208 ),
        .bank_sel(bank_sel),
        .\grn_reg[0] (\grn_reg[0]_2 ),
        .\grn_reg[0]_0 (\grn_reg[0]_3 ),
        .\grn_reg[10] (\grn_reg[10]_1 ),
        .\grn_reg[10]_0 (\grn_reg[10]_2 ),
        .\grn_reg[11] (\grn_reg[11]_1 ),
        .\grn_reg[11]_0 (\grn_reg[11]_2 ),
        .\grn_reg[12] (\grn_reg[12]_1 ),
        .\grn_reg[12]_0 (\grn_reg[12]_2 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[13]_0 (\grn_reg[13]_2 ),
        .\grn_reg[14] (\grn_reg[14]_2 ),
        .\grn_reg[14]_0 (\grn_reg[14]_3 ),
        .\grn_reg[15] (\grn_reg[15]_6 ),
        .\grn_reg[15]_0 (\grn_reg[15]_7 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (\grn_reg[1]_2 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (\grn_reg[2]_2 ),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (\grn_reg[3]_2 ),
        .\grn_reg[4] (\grn_reg[4]_4 ),
        .\grn_reg[4]_0 (\grn_reg[4]_5 ),
        .\grn_reg[5] (\grn_reg[5]_1 ),
        .\grn_reg[5]_0 (\grn_reg[5]_2 ),
        .\grn_reg[6] (\grn_reg[6]_1 ),
        .\grn_reg[6]_0 (\grn_reg[6]_2 ),
        .\grn_reg[7] (\grn_reg[7]_1 ),
        .\grn_reg[7]_0 (\grn_reg[7]_2 ),
        .\grn_reg[8] (a1buso_n_30),
        .\grn_reg[8]_0 (a1buso_n_31),
        .\grn_reg[9] (\grn_reg[9]_1 ),
        .\grn_reg[9]_0 (\grn_reg[9]_2 ),
        .\i_/badr[15]_INST_0_i_19_0 (\i_/badr[15]_INST_0_i_19 ),
        .\i_/badr[15]_INST_0_i_19_1 (\i_/badr[15]_INST_0_i_19_0 ),
        .\i_/badr[15]_INST_0_i_19_2 (\i_/badr[15]_INST_0_i_19_1 ),
        .\i_/badr[15]_INST_0_i_19_3 (gr02),
        .\i_/badr[15]_INST_0_i_19_4 (gr01),
        .\i_/badr[15]_INST_0_i_4_0 (\sr[6]_i_11_7 [1:0]),
        .out(gr00),
        .p_1_in1_in(p_1_in1_in),
        .\rgf_c1bus_wb[4]_i_47 (gr07),
        .\rgf_c1bus_wb[4]_i_47_0 (gr03),
        .\rgf_c1bus_wb[4]_i_47_1 (gr04));
  mcss_rgf_bank_bus_31 a1buso2l
       (.a1bus_sel_0(a1bus_sel_0),
        .\badr[0]_INST_0_i_1 (\sr[4]_i_210_0 ),
        .\badr[10]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_28_0 ),
        .\badr[11]_INST_0_i_1 (\sr[4]_i_207_0 ),
        .\badr[12]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_24_0 ),
        .\badr[13]_INST_0_i_1 (\sr[4]_i_209_0 ),
        .\badr[14]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_23_0 ),
        .\badr[15]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_22_0 ),
        .\badr[15]_INST_0_i_20 (\sr[6]_i_11_7 [1:0]),
        .\badr[1]_INST_0_i_1 (\sr[4]_i_213_0 ),
        .\badr[2]_INST_0_i_1 (\sr[4]_i_211_0 ),
        .\badr[3]_INST_0_i_1 (\sr[4]_i_220_1 ),
        .\badr[4]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_25_0 ),
        .\badr[5]_INST_0_i_1 (\sr[4]_i_224_1 ),
        .\badr[6]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_26_0 ),
        .\badr[7]_INST_0_i_1 (\sr[4]_i_225_1 ),
        .\badr[8]_INST_0_i_1 (\rgf_c1bus_wb[4]_i_27_0 ),
        .\badr[9]_INST_0_i_1 (\sr[4]_i_208_0 ),
        .\grn_reg[0] (\grn_reg[0]_7 ),
        .\grn_reg[0]_0 (\grn_reg[0]_8 ),
        .\grn_reg[0]_1 (a1buso2l_n_63),
        .\grn_reg[10] (\grn_reg[10]_5 ),
        .\grn_reg[10]_0 (\grn_reg[10]_6 ),
        .\grn_reg[10]_1 (a1buso2l_n_44),
        .\grn_reg[11] (\grn_reg[11]_5 ),
        .\grn_reg[11]_0 (\grn_reg[11]_6 ),
        .\grn_reg[11]_1 (a1buso2l_n_42),
        .\grn_reg[12] (\grn_reg[12]_5 ),
        .\grn_reg[12]_0 (\grn_reg[12]_6 ),
        .\grn_reg[12]_1 (a1buso2l_n_40),
        .\grn_reg[13] (\grn_reg[13]_5 ),
        .\grn_reg[13]_0 (\grn_reg[13]_6 ),
        .\grn_reg[13]_1 (a1buso2l_n_38),
        .\grn_reg[14] (\grn_reg[14]_6 ),
        .\grn_reg[14]_0 (\grn_reg[14]_7 ),
        .\grn_reg[14]_1 (a1buso2l_n_36),
        .\grn_reg[15] (\grn_reg[15]_11 ),
        .\grn_reg[15]_0 (\grn_reg[15]_12 ),
        .\grn_reg[15]_1 (a1buso2l_n_34),
        .\grn_reg[1] (\grn_reg[1]_5 ),
        .\grn_reg[1]_0 (\grn_reg[1]_6 ),
        .\grn_reg[1]_1 (a1buso2l_n_61),
        .\grn_reg[2] (\grn_reg[2]_5 ),
        .\grn_reg[2]_0 (\grn_reg[2]_6 ),
        .\grn_reg[2]_1 (a1buso2l_n_59),
        .\grn_reg[3] (\grn_reg[3]_5 ),
        .\grn_reg[3]_0 (\grn_reg[3]_6 ),
        .\grn_reg[3]_1 (a1buso2l_n_57),
        .\grn_reg[4] (\grn_reg[4]_9 ),
        .\grn_reg[4]_0 (\grn_reg[4]_10 ),
        .\grn_reg[4]_1 (a1buso2l_n_55),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\grn_reg[5]_1 (a1buso2l_n_53),
        .\grn_reg[6] (\grn_reg[6]_5 ),
        .\grn_reg[6]_0 (\grn_reg[6]_6 ),
        .\grn_reg[6]_1 (a1buso2l_n_51),
        .\grn_reg[7] (\grn_reg[7]_5 ),
        .\grn_reg[7]_0 (\grn_reg[7]_6 ),
        .\grn_reg[7]_1 (a1buso2l_n_49),
        .\grn_reg[8] (a1buso2l_n_23),
        .\grn_reg[8]_0 (a1buso2l_n_47),
        .\grn_reg[9] (\grn_reg[9]_5 ),
        .\grn_reg[9]_0 (\grn_reg[9]_6 ),
        .\grn_reg[9]_1 (a1buso2l_n_46),
        .\i_/badr[0]_INST_0_i_17_0 (\i_/badr[15]_INST_0_i_19 ),
        .\i_/badr[0]_INST_0_i_17_1 (\i_/badr[15]_INST_0_i_19_0 ),
        .\i_/badr[0]_INST_0_i_17_2 (\i_/badr[15]_INST_0_i_19_1 ),
        .\i_/badr[15]_INST_0_i_23_0 (gr22),
        .\i_/badr[15]_INST_0_i_23_1 (gr21),
        .\i_/badr[15]_INST_0_i_23_2 (\i_/badr[15]_INST_0_i_47 ),
        .out(gr20),
        .p_0_in0_in(p_0_in0_in),
        .\rgf_c1bus_wb[4]_i_33 (\rgf_c1bus_wb[4]_i_33 ),
        .\rgf_c1bus_wb[4]_i_33_0 (\rgf_c1bus_wb[4]_i_33_0 ),
        .\rgf_c1bus_wb[4]_i_37 (\rgf_c1bus_wb[4]_i_37 ),
        .\rgf_c1bus_wb[4]_i_37_0 (\rgf_c1bus_wb[4]_i_37_0 ),
        .\rgf_c1bus_wb[4]_i_39 (gr27),
        .\rgf_c1bus_wb[4]_i_41 (\rgf_c1bus_wb[4]_i_41 ),
        .\rgf_c1bus_wb[4]_i_41_0 (\rgf_c1bus_wb[4]_i_41_0 ),
        .\rgf_c1bus_wb[4]_i_47 (gr23),
        .\rgf_c1bus_wb[4]_i_47_0 (gr24),
        .\rgf_c1bus_wb[4]_i_47_1 (\rgf_c1bus_wb[4]_i_47 ),
        .\rgf_c1bus_wb[4]_i_47_2 (\rgf_c1bus_wb[4]_i_47_0 ),
        .\rgf_c1bus_wb[4]_i_47_3 ({gr26[15:9],gr26[7:0]}),
        .\rgf_c1bus_wb[4]_i_51 (\rgf_c1bus_wb[4]_i_51 ),
        .\rgf_c1bus_wb[4]_i_51_0 (\rgf_c1bus_wb[4]_i_51_0 ),
        .\rgf_c1bus_wb[4]_i_53 (\rgf_c1bus_wb[4]_i_53 ),
        .\rgf_c1bus_wb[4]_i_53_0 (\rgf_c1bus_wb[4]_i_53_0 ),
        .\rgf_c1bus_wb[4]_i_57 (\rgf_c1bus_wb[4]_i_57 ),
        .\rgf_c1bus_wb[4]_i_57_0 (\rgf_c1bus_wb[4]_i_57_0 ),
        .\rgf_c1bus_wb[4]_i_61 (\rgf_c1bus_wb[4]_i_61 ),
        .\rgf_c1bus_wb[4]_i_61_0 (\rgf_c1bus_wb[4]_i_61_0 ),
        .\rgf_c1bus_wb[4]_i_65 (\rgf_c1bus_wb[4]_i_65 ),
        .\rgf_c1bus_wb[4]_i_65_0 (\rgf_c1bus_wb[4]_i_65_0 ),
        .\rgf_c1bus_wb[4]_i_67 (\rgf_c1bus_wb[4]_i_67 ),
        .\rgf_c1bus_wb[4]_i_67_0 (\rgf_c1bus_wb[4]_i_67_0 ),
        .\sr[4]_i_235 (\sr[4]_i_235 ),
        .\sr[4]_i_235_0 (\sr[4]_i_235_0 ),
        .\sr[4]_i_237 (\sr[4]_i_237 ),
        .\sr[4]_i_237_0 (\sr[4]_i_237_0 ),
        .\sr[4]_i_240 (\sr[4]_i_240 ),
        .\sr[4]_i_240_0 (\sr[4]_i_240_0 ),
        .\sr[4]_i_243 (\sr[4]_i_243 ),
        .\sr[4]_i_243_0 (\sr[4]_i_243_0 ),
        .\sr[4]_i_245 (\sr[4]_i_245 ),
        .\sr[4]_i_245_0 (\sr[4]_i_245_0 ),
        .\sr_reg[0] (gr6_bus1));
  mcss_rgf_bank_bus_32 b0buso
       (.b0bus_sel_0(b0bus_sel_0),
        .bank_sel(bank_sel),
        .\bbus_o[0]_INST_0_i_1 (\bbus_o[0]_INST_0_i_1 ),
        .\bbus_o[1]_INST_0_i_1 (\bbus_o[1]_INST_0_i_1 ),
        .\bbus_o[2]_INST_0_i_1 (\bbus_o[2]_INST_0_i_1 ),
        .\bbus_o[3]_INST_0_i_1 (\bbus_o[3]_INST_0_i_1 ),
        .\bbus_o[4]_INST_0_i_1 (\bbus_o[4]_INST_0_i_1 ),
        .\bdatw[15]_INST_0_i_1 (gr07),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[4] (\grn_reg[4]_3 ),
        .\i_/bdatw[15]_INST_0_i_24_0 (\i_/bdatw[15]_INST_0_i_24 ),
        .\i_/bdatw[15]_INST_0_i_24_1 (\i_/bdatw[15]_INST_0_i_24_0 ),
        .\i_/bdatw[15]_INST_0_i_27_0 (gr04),
        .\i_/bdatw[15]_INST_0_i_27_1 (gr03),
        .\i_/bdatw[15]_INST_0_i_27_2 (\sr[6]_i_11_7 [1:0]),
        .\i_/bdatw[15]_INST_0_i_77_0 (\i_/bdatw[15]_INST_0_i_77 ),
        .\i_/bdatw[15]_INST_0_i_9_0 (gr02),
        .\i_/bdatw[15]_INST_0_i_9_1 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_9_2 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .\i_/bdatw[15]_INST_0_i_9_3 (\i_/bdatw[15]_INST_0_i_9_1 ),
        .\i_/bdatw[15]_INST_0_i_9_4 (\i_/bdatw[15]_INST_0_i_9_2 ),
        .\i_/bdatw[15]_INST_0_i_9_5 (gr06),
        .\i_/bdatw[15]_INST_0_i_9_6 (gr05),
        .\i_/bdatw[15]_INST_0_i_9_7 (gr01[15:5]),
        .\i_/bdatw[15]_INST_0_i_9_8 (\i_/bdatw[15]_INST_0_i_9_3 ),
        .out(gr00),
        .p_1_in3_in(p_1_in3_in));
  mcss_rgf_bank_bus_33 b0buso2l
       (.b0bus_sel_0(b0bus_sel_0),
        .\bbus_o[0]_INST_0_i_1 (\bbus_o[0]_INST_0_i_1_0 ),
        .\bbus_o[1]_INST_0_i_1 (\bbus_o[1]_INST_0_i_1_0 ),
        .\bbus_o[2]_INST_0_i_1 (\bbus_o[2]_INST_0_i_1_0 ),
        .\bbus_o[3]_INST_0_i_1 (\bbus_o[3]_INST_0_i_1_0 ),
        .\bbus_o[4]_INST_0_i_1 (\bbus_o[4]_INST_0_i_1_0 ),
        .\bdatw[15]_INST_0_i_1 (gr27),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[4] (\grn_reg[4]_8 ),
        .\i_/bdatw[15]_INST_0_i_10_0 (gr21[15:5]),
        .\i_/bdatw[15]_INST_0_i_10_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_10_2 (\i_/bdatw[15]_INST_0_i_9_3 ),
        .\i_/bdatw[15]_INST_0_i_10_3 (\i_/bdatw[15]_INST_0_i_9_0 ),
        .\i_/bdatw[15]_INST_0_i_10_4 (gr26),
        .\i_/bdatw[15]_INST_0_i_10_5 (gr25),
        .\i_/bdatw[15]_INST_0_i_10_6 (\i_/bdatw[15]_INST_0_i_9 ),
        .\i_/bdatw[15]_INST_0_i_28_0 (\i_/bdatw[15]_INST_0_i_9_1 ),
        .\i_/bdatw[15]_INST_0_i_28_1 (\i_/bdatw[15]_INST_0_i_9_2 ),
        .\i_/bdatw[15]_INST_0_i_28_2 (\i_/bdatw[15]_INST_0_i_24_0 ),
        .\i_/bdatw[15]_INST_0_i_28_3 (\i_/bdatw[15]_INST_0_i_24 ),
        .\i_/bdatw[15]_INST_0_i_31_0 (gr24),
        .\i_/bdatw[15]_INST_0_i_31_1 (gr23),
        .\i_/bdatw[15]_INST_0_i_31_2 (\sr[6]_i_11_7 [1:0]),
        .\i_/bdatw[15]_INST_0_i_82_0 (\i_/badr[15]_INST_0_i_47 ),
        .\i_/bdatw[15]_INST_0_i_82_1 (\i_/bdatw[15]_INST_0_i_77 ),
        .out(gr20),
        .p_0_in2_in(p_0_in2_in));
  mcss_rgf_bank_bus_34 b1buso
       (.bank_sel(bank_sel),
        .\bdatw[15]_INST_0_i_14 (gr07),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (b1buso_n_15),
        .\grn_reg[0]_0 (b1buso_n_20),
        .\grn_reg[0]_1 (b1buso_n_25),
        .\grn_reg[10] (b1buso_n_5),
        .\grn_reg[11] (b1buso_n_4),
        .\grn_reg[12] (b1buso_n_3),
        .\grn_reg[13] (b1buso_n_2),
        .\grn_reg[14] (b1buso_n_1),
        .\grn_reg[15] (\grn_reg[15]_8 ),
        .\grn_reg[1] (b1buso_n_14),
        .\grn_reg[1]_0 (b1buso_n_19),
        .\grn_reg[1]_1 (b1buso_n_24),
        .\grn_reg[2] (b1buso_n_13),
        .\grn_reg[2]_0 (b1buso_n_18),
        .\grn_reg[2]_1 (b1buso_n_23),
        .\grn_reg[3] (b1buso_n_12),
        .\grn_reg[3]_0 (b1buso_n_17),
        .\grn_reg[3]_1 (b1buso_n_22),
        .\grn_reg[4] (b1buso_n_11),
        .\grn_reg[4]_0 (b1buso_n_16),
        .\grn_reg[4]_1 (b1buso_n_21),
        .\grn_reg[5] (b1buso_n_10),
        .\grn_reg[6] (b1buso_n_9),
        .\grn_reg[7] (b1buso_n_8),
        .\grn_reg[8] (b1buso_n_7),
        .\grn_reg[9] (b1buso_n_6),
        .\i_/bdatw[15]_INST_0_i_112_0 (\i_/bdatw[15]_INST_0_i_112 ),
        .\i_/bdatw[15]_INST_0_i_112_1 (\i_/bdatw[15]_INST_0_i_112_0 ),
        .\i_/bdatw[15]_INST_0_i_112_2 (\i_/bdatw[15]_INST_0_i_112_1 ),
        .\i_/bdatw[15]_INST_0_i_113_0 (\i_/bdatw[15]_INST_0_i_113 ),
        .\i_/bdatw[15]_INST_0_i_113_1 (gr02),
        .\i_/bdatw[15]_INST_0_i_113_2 (gr01),
        .\i_/bdatw[15]_INST_0_i_44_0 (\sr[6]_i_11_7 [1:0]),
        .\i_/bdatw[15]_INST_0_i_44_1 (gr06),
        .\i_/bdatw[15]_INST_0_i_44_2 (gr05),
        .\i_/bdatw[15]_INST_0_i_44_3 (\i_/bdatw[15]_INST_0_i_44 ),
        .\i_/bdatw[15]_INST_0_i_44_4 (gr03),
        .\i_/bdatw[15]_INST_0_i_44_5 (gr04),
        .out(gr00));
  mcss_rgf_bank_bus_35 b1buso2l
       (.\bdatw[15]_INST_0_i_14 (gr27),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (b1buso2l_n_15),
        .\grn_reg[0]_0 (b1buso2l_n_20),
        .\grn_reg[0]_1 (b1buso2l_n_25),
        .\grn_reg[10] (b1buso2l_n_5),
        .\grn_reg[11] (b1buso2l_n_4),
        .\grn_reg[12] (b1buso2l_n_3),
        .\grn_reg[13] (b1buso2l_n_2),
        .\grn_reg[14] (b1buso2l_n_1),
        .\grn_reg[15] (\grn_reg[15]_13 ),
        .\grn_reg[1] (b1buso2l_n_14),
        .\grn_reg[1]_0 (b1buso2l_n_19),
        .\grn_reg[1]_1 (b1buso2l_n_24),
        .\grn_reg[2] (b1buso2l_n_13),
        .\grn_reg[2]_0 (b1buso2l_n_18),
        .\grn_reg[2]_1 (b1buso2l_n_23),
        .\grn_reg[3] (b1buso2l_n_12),
        .\grn_reg[3]_0 (b1buso2l_n_17),
        .\grn_reg[3]_1 (b1buso2l_n_22),
        .\grn_reg[4] (b1buso2l_n_11),
        .\grn_reg[4]_0 (b1buso2l_n_16),
        .\grn_reg[4]_1 (b1buso2l_n_21),
        .\grn_reg[5] (b1buso2l_n_10),
        .\grn_reg[6] (b1buso2l_n_9),
        .\grn_reg[7] (b1buso2l_n_8),
        .\grn_reg[8] (b1buso2l_n_7),
        .\grn_reg[9] (b1buso2l_n_6),
        .\i_/bdatw[15]_INST_0_i_110_0 (\i_/badr[15]_INST_0_i_47 ),
        .\i_/bdatw[15]_INST_0_i_110_1 (\i_/bdatw[15]_INST_0_i_112 ),
        .\i_/bdatw[15]_INST_0_i_110_2 (\i_/bdatw[15]_INST_0_i_112_0 ),
        .\i_/bdatw[15]_INST_0_i_110_3 (\i_/bdatw[15]_INST_0_i_112_1 ),
        .\i_/bdatw[15]_INST_0_i_111_0 (\i_/bdatw[15]_INST_0_i_44 ),
        .\i_/bdatw[15]_INST_0_i_111_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_111_2 (gr21),
        .\i_/bdatw[15]_INST_0_i_200_0 (\sr[6]_i_11_7 [1:0]),
        .\i_/bdatw[15]_INST_0_i_200_1 (\i_/bdatw[15]_INST_0_i_113 ),
        .\i_/bdatw[15]_INST_0_i_43_0 (gr23),
        .\i_/bdatw[15]_INST_0_i_43_1 (gr24),
        .\i_/bdatw[15]_INST_0_i_43_2 (gr26),
        .\i_/bdatw[15]_INST_0_i_43_3 (gr25),
        .out(gr20));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[5]_INST_0 
       (.I0(\tr_reg[5]_0 ),
        .I1(\bbus_o[5]_3 ),
        .O(bbus_o));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(\bdatw[10]_3 ),
        .I1(\bdatw[10]_4 ),
        .I2(\bdatw[10]_5 ),
        .I3(p_1_in3_in[10]),
        .I4(p_0_in2_in[10]),
        .I5(\bdatw[10]_6 ),
        .O(\tr_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(\bdatw[10] ),
        .I1(\bdatw[10]_0 ),
        .I2(\bdatw[10]_1 ),
        .I3(b1buso_n_5),
        .I4(b1buso2l_n_5),
        .I5(\bdatw[10]_2 ),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[10]_INST_0_i_42 
       (.I0(b1buso_n_23),
        .I1(b1buso_n_13),
        .I2(b1buso_n_18),
        .I3(b1buso2l_n_13),
        .I4(b1buso2l_n_18),
        .I5(b1buso2l_n_23),
        .O(b1bus_b02[2]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(\bdatw[11]_3 ),
        .I1(\bdatw[11]_4 ),
        .I2(\bdatw[11]_5 ),
        .I3(p_1_in3_in[11]),
        .I4(p_0_in2_in[11]),
        .I5(\bdatw[11]_6 ),
        .O(\tr_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(\bdatw[11] ),
        .I1(\bdatw[11]_0 ),
        .I2(\bdatw[11]_1 ),
        .I3(b1buso_n_4),
        .I4(b1buso2l_n_4),
        .I5(\bdatw[11]_2 ),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[11]_INST_0_i_43 
       (.I0(b1buso_n_22),
        .I1(b1buso_n_12),
        .I2(b1buso_n_17),
        .I3(b1buso2l_n_12),
        .I4(b1buso2l_n_17),
        .I5(b1buso2l_n_22),
        .O(b1bus_b02[3]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(\bdatw[12]_3 ),
        .I1(\bdatw[12]_4 ),
        .I2(\bdatw[12]_5 ),
        .I3(p_1_in3_in[12]),
        .I4(p_0_in2_in[12]),
        .I5(\bdatw[12]_6 ),
        .O(\tr_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(\bdatw[12] ),
        .I1(\bdatw[12]_0 ),
        .I2(\bdatw[12]_1 ),
        .I3(b1buso_n_3),
        .I4(b1buso2l_n_3),
        .I5(\bdatw[12]_2 ),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[12]_INST_0_i_41 
       (.I0(b1buso_n_21),
        .I1(b1buso_n_11),
        .I2(b1buso_n_16),
        .I3(b1buso2l_n_11),
        .I4(b1buso2l_n_16),
        .I5(b1buso2l_n_21),
        .O(b1bus_b02[4]));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[13]_INST_0 
       (.I0(\tr_reg[13] ),
        .I1(\bdatw[13] ),
        .I2(\tr_reg[13]_0 ),
        .I3(\bdatw[13]_0 ),
        .I4(\stat_reg[1]_0 ),
        .I5(\bdatw[13]_1 ),
        .O(bdatw[0]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(\bdatw[13]_6 ),
        .I1(\bdatw[13]_7 ),
        .I2(\bdatw[13]_8 ),
        .I3(p_1_in3_in[13]),
        .I4(p_0_in2_in[13]),
        .I5(\bdatw[13]_9 ),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13]_2 ),
        .I1(\bdatw[13]_3 ),
        .I2(\bdatw[13]_4 ),
        .I3(b1buso_n_2),
        .I4(b1buso2l_n_2),
        .I5(\bdatw[13]_5 ),
        .O(\tr_reg[13]_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(\tr_reg[5]_0 ),
        .I1(\bdatw[13] ),
        .I2(\tr_reg[5] ),
        .O(\stat_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[14]_INST_0 
       (.I0(\tr_reg[14] ),
        .I1(\bdatw[13] ),
        .I2(\tr_reg[14]_0 ),
        .I3(\bdatw[13]_0 ),
        .I4(\stat_reg[1] ),
        .I5(\bdatw[13]_1 ),
        .O(bdatw[1]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(\bdatw[14]_3 ),
        .I1(\bdatw[14]_4 ),
        .I2(\bdatw[14]_5 ),
        .I3(p_1_in3_in[14]),
        .I4(p_0_in2_in[14]),
        .I5(\bdatw[14]_6 ),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(\bdatw[14] ),
        .I1(\bdatw[14]_0 ),
        .I2(\bdatw[14]_1 ),
        .I3(b1buso_n_1),
        .I4(b1buso2l_n_1),
        .I5(\bdatw[14]_2 ),
        .O(\tr_reg[14]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(\tr_reg[6]_0 ),
        .I1(\bdatw[13] ),
        .I2(\tr_reg[6] ),
        .O(\stat_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(\bdatw[15] ),
        .I1(\bdatw[15]_0 ),
        .I2(\bdatw[15]_1 ),
        .I3(p_1_in3_in[15]),
        .I4(p_0_in2_in[15]),
        .I5(\bdatw[15]_2 ),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[15]_INST_0_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_19 ),
        .I1(\rgf_c1bus_wb[15]_i_19_0 ),
        .I2(\rgf_c1bus_wb[15]_i_19_1 ),
        .I3(b1buso_n_8),
        .I4(b1buso2l_n_8),
        .I5(\rgf_c1bus_wb[15]_i_19_2 ),
        .O(\tr_reg[7]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(\tr_reg[7] ),
        .I1(\bdatw[13] ),
        .I2(\tr_reg[7]_0 ),
        .O(\stat_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(\bdatw[8]_3 ),
        .I1(\bdatw[8]_4 ),
        .I2(\bdatw[8]_5 ),
        .I3(p_1_in3_in[8]),
        .I4(p_0_in2_in[8]),
        .I5(\bdatw[8]_6 ),
        .O(\tr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(\bdatw[8] ),
        .I1(\bdatw[8]_0 ),
        .I2(\bdatw[8]_1 ),
        .I3(b1buso_n_7),
        .I4(b1buso2l_n_7),
        .I5(\bdatw[8]_2 ),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_42 
       (.I0(b1buso_n_25),
        .I1(b1buso_n_15),
        .I2(b1buso_n_20),
        .I3(b1buso2l_n_15),
        .I4(b1buso2l_n_20),
        .I5(b1buso2l_n_25),
        .O(b1bus_b02[0]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(\bdatw[9]_3 ),
        .I1(\bdatw[9]_4 ),
        .I2(\bdatw[9]_5 ),
        .I3(p_1_in3_in[9]),
        .I4(p_0_in2_in[9]),
        .I5(\bdatw[9]_6 ),
        .O(\tr_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(\bdatw[9] ),
        .I1(\bdatw[9]_0 ),
        .I2(\bdatw[9]_1 ),
        .I3(b1buso_n_6),
        .I4(b1buso2l_n_6),
        .I5(\bdatw[9]_2 ),
        .O(\tr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[9]_INST_0_i_41 
       (.I0(b1buso_n_24),
        .I1(b1buso_n_14),
        .I2(b1buso_n_19),
        .I3(b1buso2l_n_14),
        .I4(b1buso2l_n_19),
        .I5(b1buso2l_n_24),
        .O(b1bus_b02[1]));
  mcss_rgf_grn_36 grn00
       (.Q(gr00),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ),
        .\grn_reg[15]_1 (\grn_reg[15]_15 ));
  mcss_rgf_grn_37 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_16 ),
        .\grn_reg[15]_1 (\grn_reg[15]_17 ));
  mcss_rgf_grn_38 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_18 ),
        .\grn_reg[15]_1 (\grn_reg[15]_19 ));
  mcss_rgf_grn_39 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_20 ),
        .\grn_reg[15]_1 (\grn_reg[15]_21 ));
  mcss_rgf_grn_40 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_22 ),
        .\grn_reg[15]_1 (\grn_reg[15]_23 ));
  mcss_rgf_grn_41 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_24 ),
        .\grn_reg[15]_1 (\grn_reg[15]_25 ));
  mcss_rgf_grn_42 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_26 ),
        .\grn_reg[15]_1 (\grn_reg[15]_27 ));
  mcss_rgf_grn_43 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_28 ),
        .\grn_reg[15]_1 (\grn_reg[15]_29 ));
  mcss_rgf_grn_44 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_30 ),
        .\grn_reg[15]_1 (\grn_reg[15]_31 ));
  mcss_rgf_grn_45 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_32 ),
        .\grn_reg[15]_1 (\grn_reg[15]_33 ));
  mcss_rgf_grn_46 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_34 ),
        .\grn_reg[15]_1 (\grn_reg[15]_35 ));
  mcss_rgf_grn_47 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_36 ),
        .\grn_reg[15]_1 (\grn_reg[15]_37 ));
  mcss_rgf_grn_48 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_38 ),
        .\grn_reg[15]_1 (\grn_reg[15]_39 ));
  mcss_rgf_grn_49 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_40 ),
        .\grn_reg[15]_1 (\grn_reg[15]_41 ));
  mcss_rgf_grn_50 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_42 ),
        .\grn_reg[15]_1 (\grn_reg[15]_43 ));
  mcss_rgf_grn_51 grn27
       (.Q(gr27),
        .SR(SR),
        .\badr[0]_INST_0_i_1 (\badr[0]_INST_0_i_1 ),
        .\badr[10]_INST_0_i_1 (\badr[10]_INST_0_i_1_1 ),
        .\badr[10]_INST_0_i_1_0 (\badr[10]_INST_0_i_1 ),
        .\badr[10]_INST_0_i_2 (\badr[10]_INST_0_i_2_0 ),
        .\badr[10]_INST_0_i_2_0 (\badr[10]_INST_0_i_2 ),
        .\badr[11]_INST_0_i_1 (\badr[11]_INST_0_i_1 ),
        .\badr[11]_INST_0_i_2 (\badr[11]_INST_0_i_2 ),
        .\badr[12]_INST_0_i_1 (\badr[12]_INST_0_i_1 ),
        .\badr[12]_INST_0_i_2 (\badr[12]_INST_0_i_2 ),
        .\badr[12]_INST_0_i_2_0 (\badr[12]_INST_0_i_2_0 ),
        .\badr[13]_INST_0_i_1 (\badr[13]_INST_0_i_1 ),
        .\badr[14]_INST_0_i_1 (\badr[14]_INST_0_i_1 ),
        .\badr[14]_INST_0_i_1_0 (\badr[14]_INST_0_i_1_0 ),
        .\badr[14]_INST_0_i_2 (\badr[14]_INST_0_i_2 ),
        .\badr[14]_INST_0_i_2_0 (\badr[14]_INST_0_i_2_0 ),
        .\badr[14]_INST_0_i_2_1 (\badr[14]_INST_0_i_2_1 ),
        .\badr[15]_INST_0_i_1 (\badr[15]_INST_0_i_1 ),
        .\badr[15]_INST_0_i_1_0 (\badr[15]_INST_0_i_1_0 ),
        .\badr[1]_INST_0_i_2 (\badr[1]_INST_0_i_2 ),
        .\badr[1]_INST_0_i_2_0 (\badr[1]_INST_0_i_2_0 ),
        .\badr[2]_INST_0_i_1 (\badr[2]_INST_0_i_1_1 ),
        .\badr[2]_INST_0_i_1_0 (\badr[2]_INST_0_i_1 ),
        .\badr[2]_INST_0_i_2 (\badr[2]_INST_0_i_2_0 ),
        .\badr[3]_INST_0_i_1 (\badr[3]_INST_0_i_1 ),
        .\badr[3]_INST_0_i_2 (\badr[3]_INST_0_i_2_0 ),
        .\badr[4]_INST_0_i_2 (\badr[4]_INST_0_i_2_0 ),
        .\badr[5]_INST_0_i_1 (\badr[5]_INST_0_i_1 ),
        .\badr[5]_INST_0_i_1_0 (\badr[5]_INST_0_i_1_0 ),
        .\badr[5]_INST_0_i_2 (\badr[5]_INST_0_i_2 ),
        .\badr[5]_INST_0_i_2_0 (\badr[5]_INST_0_i_2_0 ),
        .\badr[6]_INST_0_i_1 (\badr[6]_INST_0_i_1 ),
        .\badr[6]_INST_0_i_1_0 (\badr[6]_INST_0_i_1_0 ),
        .\badr[6]_INST_0_i_2 (\badr[6]_INST_0_i_2 ),
        .\badr[6]_INST_0_i_2_0 (\badr[6]_INST_0_i_2_0 ),
        .\badr[6]_INST_0_i_2_1 (\badr[6]_INST_0_i_2_1 ),
        .\badr[7]_INST_0_i_2 (\badr[7]_INST_0_i_2 ),
        .\badr[8]_INST_0_i_2 (\badr[8]_INST_0_i_2_0 ),
        .\badr[9]_INST_0_i_1 (\badr[9]_INST_0_i_1 ),
        .\badr[9]_INST_0_i_1_0 (\badr[9]_INST_0_i_1_0 ),
        .\bbus_o[5] (\bbus_o[5] ),
        .\bbus_o[5]_0 (\bbus_o[5]_0 ),
        .\bbus_o[5]_1 (\bbus_o[5]_1 ),
        .\bbus_o[5]_2 (\bbus_o[5]_2 ),
        .\bbus_o[6] (\bbus_o[6] ),
        .\bbus_o[6]_0 (\bbus_o[6]_0 ),
        .\bbus_o[6]_1 (\bbus_o[6]_1 ),
        .\bbus_o[6]_2 (\bbus_o[6]_2 ),
        .\bbus_o[7] (\bbus_o[7] ),
        .\bbus_o[7]_0 (\bbus_o[7]_0 ),
        .\bbus_o[7]_1 (\bbus_o[7]_1 ),
        .\bbus_o[7]_2 (\bbus_o[7]_2 ),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_44 ),
        .\grn_reg[15]_1 (\grn_reg[15]_45 ),
        .p_0_in2_in(p_0_in2_in[7:5]),
        .p_1_in3_in(p_1_in3_in[7:5]),
        .\rgf_c0bus_wb[0]_i_8 (\rgf_c0bus_wb[3]_i_7_3 ),
        .\rgf_c0bus_wb[10]_i_26 (\rgf_c0bus_wb[14]_i_2 ),
        .\rgf_c0bus_wb[10]_i_26_0 (\rgf_c0bus_wb[14]_i_13_3 ),
        .\rgf_c0bus_wb[10]_i_26_1 (\rgf_c0bus_wb[3]_i_7_4 ),
        .\rgf_c0bus_wb[10]_i_4 (\rgf_c0bus_wb[10]_i_4 ),
        .\rgf_c0bus_wb[10]_i_8_0 (\rgf_c0bus_wb[10]_i_8 ),
        .\rgf_c0bus_wb[11]_i_17 (\rgf_c0bus_wb[14]_i_13_0 ),
        .\rgf_c0bus_wb[11]_i_17_0 (\rgf_c0bus_wb[3]_i_7_0 ),
        .\rgf_c0bus_wb[11]_i_17_1 (\rgf_c0bus_wb[3]_i_7_1 ),
        .\rgf_c0bus_wb[11]_i_17_2 (\rgf_c0bus_wb[14]_i_13_4 ),
        .\rgf_c0bus_wb[11]_i_17_3 (\rgf_c0bus_wb[14]_i_13_5 ),
        .\rgf_c0bus_wb[11]_i_17_4 (\rgf_c0bus_wb[14]_i_13_6 ),
        .\rgf_c0bus_wb[11]_i_22 (\rgf_c0bus_wb[11]_i_22_0 ),
        .\rgf_c0bus_wb[11]_i_3 (\rgf_c0bus_wb[11]_i_3 ),
        .\rgf_c0bus_wb[11]_i_3_0 (\rgf_c0bus_wb[11]_i_3_0 ),
        .\rgf_c0bus_wb[11]_i_3_1 (\rgf_c0bus_wb[11]_i_3_1 ),
        .\rgf_c0bus_wb[11]_i_3_2 (\rgf_c0bus_wb[11]_i_3_3 ),
        .\rgf_c0bus_wb[11]_i_9 (\rgf_c0bus_wb[11]_i_9_0 ),
        .\rgf_c0bus_wb[11]_i_9_0 (\rgf_c0bus_wb[11]_i_9_2 ),
        .\rgf_c0bus_wb[11]_i_9_1 (\rgf_c0bus_wb[11]_i_9_3 ),
        .\rgf_c0bus_wb[11]_i_9_2 (\rgf_c0bus_wb[11]_i_9_4 ),
        .\rgf_c0bus_wb[13]_i_28_0 (\rgf_c0bus_wb[13]_i_28 ),
        .\rgf_c0bus_wb[13]_i_29_0 (\rgf_c0bus_wb[13]_i_29 ),
        .\rgf_c0bus_wb[13]_i_4 (\rgf_c0bus_wb[13]_i_4 ),
        .\rgf_c0bus_wb[15]_i_18_0 (\rgf_c0bus_wb[15]_i_18 ),
        .\rgf_c0bus_wb[15]_i_26_0 (\rgf_c0bus_wb[15]_i_26 ),
        .\rgf_c0bus_wb[15]_i_6 (\rgf_c0bus_wb[15]_i_6 ),
        .\rgf_c0bus_wb[15]_i_6_0 (\rgf_c0bus_wb[15]_i_6_0 ),
        .\rgf_c0bus_wb[15]_i_6_1 (\rgf_c0bus_wb[15]_i_6_1 ),
        .\rgf_c0bus_wb[1]_i_3 (\sr[4]_i_67 ),
        .\rgf_c0bus_wb[3]_i_7 (\sr[6]_i_11_7 [2]),
        .\rgf_c0bus_wb[4]_i_3 (\rgf_c0bus_wb[4]_i_3 ),
        .\rgf_c0bus_wb[5]_i_2 (\badr[9]_INST_0_i_2 ),
        .\rgf_c0bus_wb[5]_i_8 (\rgf_c0bus_wb[3]_i_7 ),
        .\rgf_c0bus_wb[5]_i_8_0 (\rgf_c0bus_wb[3]_i_18_0 ),
        .\rgf_c0bus_wb[5]_i_8_1 (\rgf_c0bus_wb[8]_i_2 ),
        .\rgf_c0bus_wb[5]_i_8_2 (\rgf_c0bus_wb[3]_i_7_2 ),
        .\rgf_c0bus_wb[6]_i_11 (\rgf_c0bus_wb[6]_i_11 ),
        .\rgf_c0bus_wb[7]_i_15_0 (\rgf_c0bus_wb[14]_i_13 ),
        .\rgf_c0bus_wb[7]_i_15_1 (\rgf_c0bus_wb[12]_i_10 ),
        .\rgf_c0bus_wb[7]_i_7 (\rgf_c0bus_wb[7]_i_7 ),
        .\rgf_c0bus_wb[7]_i_7_0 (\rgf_c0bus_wb[7]_i_7_0 ),
        .\rgf_c0bus_wb_reg[10] (\rgf_c0bus_wb_reg[10]_0 ),
        .\rgf_c0bus_wb_reg[10]_0 (\rgf_c0bus_wb_reg[10] ),
        .\rgf_c0bus_wb_reg[10]_1 (\rgf_c0bus_wb_reg[10]_1 ),
        .\rgf_c0bus_wb_reg[7]_i_11 (\rgf_c0bus_wb_reg[7]_i_11 ),
        .\rgf_c1bus_wb[10]_i_14 (\sr[6]_i_15 ),
        .\rgf_c1bus_wb[10]_i_14_0 (\sr[6]_i_11_5 ),
        .\rgf_c1bus_wb[11]_i_10 (\rgf_c1bus_wb[11]_i_10 ),
        .\rgf_c1bus_wb[11]_i_11 (\sr[6]_i_11_0 ),
        .\rgf_c1bus_wb[11]_i_11_0 (\sr[6]_i_11_2 ),
        .\rgf_c1bus_wb[11]_i_11_1 (\sr[4]_i_102 ),
        .\rgf_c1bus_wb[11]_i_11_2 (\sr[4]_i_99_2 ),
        .\rgf_c1bus_wb[11]_i_11_3 (\sr[4]_i_99_1 ),
        .\rgf_c1bus_wb[11]_i_11_4 (\sr[4]_i_99_0 ),
        .\rgf_c1bus_wb[11]_i_11_5 (\sr[4]_i_99 ),
        .\rgf_c1bus_wb[11]_i_11_6 (\sr[6]_i_11_9 ),
        .\rgf_c1bus_wb[11]_i_13_0 (\rgf_c1bus_wb[11]_i_13 ),
        .\rgf_c1bus_wb[11]_i_8 (\sr[6]_i_11_3 ),
        .\rgf_c1bus_wb[11]_i_8_0 (\sr[6]_i_11_6 ),
        .\rgf_c1bus_wb[11]_i_8_1 (\sr[6]_i_11_8 ),
        .\rgf_c1bus_wb[12]_i_2 (\rgf_c1bus_wb[14]_i_28_2 ),
        .\rgf_c1bus_wb[12]_i_20 (\rgf_c1bus_wb[12]_i_20_0 ),
        .\rgf_c1bus_wb[12]_i_2_0 (\rgf_c1bus_wb[12]_i_2 ),
        .\rgf_c1bus_wb[13]_i_16_0 (\rgf_c1bus_wb[13]_i_16 ),
        .\rgf_c1bus_wb[13]_i_9_0 (\rgf_c1bus_wb[13]_i_9 ),
        .\rgf_c1bus_wb[14]_i_11 (\rgf_c1bus_wb[14]_i_11 ),
        .\rgf_c1bus_wb[14]_i_11_0 (\rgf_c1bus_wb[14]_i_11_0 ),
        .\rgf_c1bus_wb[14]_i_11_1 (\rgf_c1bus_wb[14]_i_11_1 ),
        .\rgf_c1bus_wb[14]_i_11_2 (b1buso_n_9),
        .\rgf_c1bus_wb[14]_i_11_3 (b1buso2l_n_9),
        .\rgf_c1bus_wb[14]_i_11_4 (\rgf_c1bus_wb[14]_i_11_2 ),
        .\rgf_c1bus_wb[14]_i_28 (\rgf_c1bus_wb[14]_i_28 ),
        .\rgf_c1bus_wb[14]_i_28_0 (\rgf_c1bus_wb[14]_i_28_1 ),
        .\rgf_c1bus_wb[14]_i_28_1 (\rgf_c1bus_wb[14]_i_28_0 ),
        .\rgf_c1bus_wb[14]_i_28_2 (\rgf_c1bus_wb[14]_i_28_4 ),
        .\rgf_c1bus_wb[14]_i_28_3 (\rgf_c1bus_wb[14]_i_28_5 ),
        .\rgf_c1bus_wb[14]_i_3 (\sr[6]_i_11 ),
        .\rgf_c1bus_wb[14]_i_30_0 (\rgf_c1bus_wb[14]_i_30 ),
        .\rgf_c1bus_wb[14]_i_32_0 (\rgf_c1bus_wb[14]_i_32 ),
        .\rgf_c1bus_wb[14]_i_32_1 (\rgf_c1bus_wb[14]_i_32_0 ),
        .\rgf_c1bus_wb[15]_i_14 (\rgf_c1bus_wb[15]_i_14_3 ),
        .\rgf_c1bus_wb[1]_i_14 (\rgf_c1bus_wb[1]_i_14_0 ),
        .\rgf_c1bus_wb[1]_i_3 (\rgf_c1bus_wb[14]_i_28_3 ),
        .\rgf_c1bus_wb[2]_i_7 (\sr[4]_i_77 ),
        .\rgf_c1bus_wb[2]_i_7_0 (\sr[4]_i_77_0 ),
        .\rgf_c1bus_wb[2]_i_7_1 (\sr[4]_i_77_1 ),
        .\rgf_c1bus_wb[2]_i_7_2 (\sr[4]_i_77_2 ),
        .\rgf_c1bus_wb[3]_i_4 (\badr[10]_INST_0_i_1_0 ),
        .\rgf_c1bus_wb[3]_i_4_0 (\badr[6]_INST_0_i_1_1 ),
        .\rgf_c1bus_wb[4]_i_3_0 (\rgf_c1bus_wb[4]_i_18_n_0 ),
        .\rgf_c1bus_wb[4]_i_3_1 (\rgf_c1bus_wb[4]_i_19_n_0 ),
        .\rgf_c1bus_wb[4]_i_3_2 (\sr[4]_i_119 ),
        .\rgf_c1bus_wb[4]_i_7_0 (\sr[6]_i_11_1 ),
        .\rgf_c1bus_wb[4]_i_7_1 (\rgf_c1bus_wb[4]_i_7 ),
        .\rgf_c1bus_wb[4]_i_7_2 (\grn_reg[15]_3 ),
        .\rgf_c1bus_wb[4]_i_7_3 (\rgf_c1bus_wb[4]_i_7_0 ),
        .\rgf_c1bus_wb[4]_i_7_4 (\rgf_c1bus_wb[4]_i_7_1 ),
        .\rgf_c1bus_wb[4]_i_7_5 (\sr[4]_i_171_0 ),
        .\rgf_c1bus_wb[4]_i_9_0 (\rgf_c1bus_wb[4]_i_9 ),
        .\rgf_c1bus_wb[5]_i_10 (\rgf_c1bus_wb[5]_i_10 ),
        .\rgf_c1bus_wb[7]_i_4 (\rgf_c1bus_wb[7]_i_4 ),
        .\rgf_c1bus_wb[7]_i_4_0 (\rgf_c1bus_wb[7]_i_4_0 ),
        .\rgf_c1bus_wb[8]_i_3 (\sr_reg[6]_5 ),
        .\rgf_c1bus_wb[8]_i_3_0 (\badr[15]_INST_0_i_1_1 ),
        .\rgf_c1bus_wb[9]_i_17 (\rgf_c1bus_wb[9]_i_17_0 ),
        .\rgf_c1bus_wb_reg[10] (\rgf_c1bus_wb_reg[10] ),
        .\rgf_c1bus_wb_reg[1] (\badr[2]_INST_0_i_1_0 ),
        .\rgf_c1bus_wb_reg[1]_0 (\badr[6]_INST_0_i_1_2 ),
        .\rgf_c1bus_wb_reg[3] (\rgf_c1bus_wb_reg[3] ),
        .\rgf_c1bus_wb_reg[4] (\rgf_c1bus_wb_reg[4] ),
        .\rgf_c1bus_wb_reg[5] (\rgf_c1bus_wb_reg[5] ),
        .\rgf_c1bus_wb_reg[5]_0 (\rgf_c1bus_wb_reg[5]_0 ),
        .\rgf_c1bus_wb_reg[5]_1 (\rgf_c1bus_wb_reg[5]_1 ),
        .\rgf_c1bus_wb_reg[7] (\rgf_c1bus_wb_reg[7] ),
        .\sr[4]_i_144 (\rgf_c0bus_wb[3]_i_18 ),
        .\sr[4]_i_144_0 (\rgf_c0bus_wb[14]_i_13_1 ),
        .\sr[4]_i_144_1 (\rgf_c0bus_wb[14]_i_13_2 ),
        .\sr[4]_i_56 (\badr[13]_INST_0_i_2 ),
        .\sr_reg[6] (\sr_reg[6] ),
        .\sr_reg[6]_0 (\sr_reg[6]_2 ),
        .\sr_reg[6]_1 (\sr_reg[6]_3 ),
        .\sr_reg[6]_10 (\sr_reg[6]_14 ),
        .\sr_reg[6]_11 (\sr_reg[6]_15 ),
        .\sr_reg[6]_12 (\sr_reg[6]_16 ),
        .\sr_reg[6]_13 (\sr_reg[6]_17 ),
        .\sr_reg[6]_14 (\sr_reg[6]_18 ),
        .\sr_reg[6]_15 (\sr_reg[6]_19 ),
        .\sr_reg[6]_16 (\sr_reg[6]_20 ),
        .\sr_reg[6]_17 (\sr_reg[6]_21 ),
        .\sr_reg[6]_18 (\sr_reg[6]_22 ),
        .\sr_reg[6]_19 (\sr_reg[6]_23 ),
        .\sr_reg[6]_2 (\sr_reg[6]_4 ),
        .\sr_reg[6]_20 (\sr_reg[6]_25 ),
        .\sr_reg[6]_21 (\sr_reg[6]_27 ),
        .\sr_reg[6]_22 (\sr_reg[6]_28 ),
        .\sr_reg[6]_3 (\sr_reg[6]_1 ),
        .\sr_reg[6]_4 (\sr_reg[6]_7 ),
        .\sr_reg[6]_5 (\sr_reg[6]_8 ),
        .\sr_reg[6]_6 (\sr_reg[6]_9 ),
        .\sr_reg[6]_7 (\sr_reg[6]_10 ),
        .\sr_reg[6]_8 (\sr_reg[6]_12 ),
        .\sr_reg[6]_9 (\sr_reg[6]_13 ),
        .\stat_reg[2] (\stat_reg[2] ),
        .\stat_reg[2]_0 (\stat_reg[2]_0 ),
        .\stat_reg[2]_1 (\stat_reg[2]_2 ),
        .\stat_reg[2]_2 (\stat_reg[2]_3 ),
        .tout__1_carry__0_i_7__0(tout__1_carry__0_i_7__0),
        .tout__1_carry__0_i_7__0_0(tout__1_carry__0_i_7__0_0),
        .tout__1_carry__0_i_7__0_1(tout__1_carry__0_i_7__0_1),
        .tout__1_carry__0_i_7__0_2(b1buso_n_10),
        .tout__1_carry__0_i_7__0_3(b1buso2l_n_10),
        .tout__1_carry__0_i_7__0_4(tout__1_carry__0_i_7__0_2),
        .\tr_reg[5] (\tr_reg[5] ),
        .\tr_reg[5]_0 (\tr_reg[5]_0 ),
        .\tr_reg[6] (\tr_reg[6] ),
        .\tr_reg[6]_0 (\tr_reg[6]_0 ),
        .\tr_reg[7] (\tr_reg[7] ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[10]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_13_2 ),
        .I1(\rgf_c0bus_wb[14]_i_13 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[14]_i_13_3 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[14]_i_13_1 ),
        .O(\badr[9]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[11]_i_10 
       (.I0(\rgf_c0bus_wb[3]_i_7_2 ),
        .I1(\rgf_c0bus_wb[3]_i_7_3 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[3]_i_7 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[3]_i_7_4 ),
        .O(\badr[2]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[12]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_13_6 ),
        .I1(\rgf_c0bus_wb[12]_i_10 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[14]_i_13_5 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[14]_i_13_4 ),
        .O(\badr[13]_INST_0_i_2_0 ));
  LUT6 #(
    .INIT(64'h5F5030305F503F3F)) 
    \rgf_c0bus_wb[12]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\rgf_c0bus_wb[12]_i_7 ),
        .I4(\rgf_c0bus_wb[3]_i_7_0 ),
        .I5(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_25_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[12]_i_19 
       (.I0(\rgf_c0bus_wb[14]_i_13_1 ),
        .I1(\rgf_c0bus_wb[14]_i_13_3 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[14]_i_13 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[14]_i_13_2 ),
        .O(\badr[8]_INST_0_i_2_1 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[12]_i_20 
       (.I0(\rgf_c0bus_wb[3]_i_18_0 ),
        .I1(\rgf_c0bus_wb[3]_i_18 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[3]_i_7 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[8]_i_2 ),
        .O(\badr[4]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[12]_i_21 
       (.I0(\rgf_c0bus_wb[3]_i_7_2 ),
        .I1(\rgf_c0bus_wb[3]_i_7_4 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\sr[6]_i_11_7 [2]),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[3]_i_7_3 ),
        .O(\sr_reg[6]_26 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \rgf_c0bus_wb[12]_i_22 
       (.I0(\sr[4]_i_196_5 ),
        .I1(\sr[4]_i_196_6 ),
        .I2(\sr[4]_i_196_7 ),
        .I3(\rgf_c0bus_wb[3]_i_7_1 ),
        .I4(\sr[4]_i_196_8 ),
        .I5(\sr[4]_i_196_9 ),
        .O(\rgf_c0bus_wb[12]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \rgf_c0bus_wb[12]_i_23 
       (.I0(\sr[4]_i_203_0 ),
        .I1(\sr[4]_i_203_1 ),
        .I2(\sr[4]_i_203_2 ),
        .I3(\rgf_c0bus_wb[3]_i_7_1 ),
        .I4(\sr[4]_i_203_3 ),
        .I5(\sr[4]_i_203_4 ),
        .O(\rgf_c0bus_wb[12]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \rgf_c0bus_wb[12]_i_25 
       (.I0(\sr[4]_i_196_0 ),
        .I1(\sr[4]_i_196_1 ),
        .I2(\sr[4]_i_196_2 ),
        .I3(\rgf_c0bus_wb[3]_i_7_1 ),
        .I4(\sr[4]_i_196_3 ),
        .I5(\sr[4]_i_196_4 ),
        .O(\rgf_c0bus_wb[12]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000FFF53535353)) 
    \rgf_c0bus_wb[12]_i_8 
       (.I0(\rgf_c0bus_wb[11]_i_22 ),
        .I1(\badr[8]_INST_0_i_2 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\badr[3]_INST_0_i_2 ),
        .I4(\rgf_c0bus_wb[12]_i_2 ),
        .I5(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_11_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[13]_i_21 
       (.I0(\rgf_c0bus_wb[14]_i_13_3 ),
        .I1(\rgf_c0bus_wb[14]_i_13_0 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[14]_i_13_2 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[14]_i_13_1 ),
        .O(\badr[9]_INST_0_i_2_0 ));
  LUT6 #(
    .INIT(64'h55335533F0FFF000)) 
    \rgf_c0bus_wb[14]_i_12 
       (.I0(\badr[5]_INST_0_i_2 ),
        .I1(\badr[1]_INST_0_i_2 ),
        .I2(\badr[13]_INST_0_i_2 ),
        .I3(\rgf_c0bus_wb_reg[10] ),
        .I4(\badr[9]_INST_0_i_2 ),
        .I5(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_11 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[14]_i_6 
       (.I0(\rgf_c0bus_wb[11]_i_11 ),
        .I1(\rgf_c0bus_wb[14]_i_2 ),
        .O(\rgf_c0bus_wb[11]_i_3_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_25 
       (.I0(\rgf_c0bus_wb[12]_i_10 ),
        .I1(\rgf_c0bus_wb[15]_i_14 ),
        .O(\rgf_c0bus_wb[0]_i_14 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_21 
       (.I0(\rgf_c0bus_wb[4]_i_7_0 ),
        .I1(\rgf_c0bus_wb[4]_i_7_1 ),
        .I2(\rgf_c0bus_wb[4]_i_7_2 ),
        .I3(\rgf_c0bus_wb[3]_i_7_1 ),
        .I4(\rgf_c0bus_wb[4]_i_7 ),
        .I5(\rgf_c0bus_wb[4]_i_7_3 ),
        .O(\sr_reg[15] ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[7]_i_10 
       (.I0(\badr[8]_INST_0_i_2_1 ),
        .I1(\rgf_c0bus_wb_reg[10] ),
        .I2(\badr[12]_INST_0_i_2_0 ),
        .O(\rgf_c0bus_wb[11]_i_8 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \rgf_c0bus_wb[7]_i_8 
       (.I0(\rgf_c0bus_wb[14]_i_13_3 ),
        .I1(\rgf_c0bus_wb[14]_i_13_1 ),
        .I2(\rgf_c0bus_wb[14]_i_13_5 ),
        .I3(\rgf_c0bus_wb[3]_i_7_1 ),
        .I4(\rgf_c0bus_wb[14]_i_13_0 ),
        .I5(\rgf_c0bus_wb[3]_i_7_0 ),
        .O(\rgf_c0bus_wb[11]_i_22 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c0bus_wb[8]_i_12 
       (.I0(\badr[13]_INST_0_i_2_0 ),
        .I1(\badr[9]_INST_0_i_2_0 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .O(\rgf_c0bus_wb[11]_i_9_1 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[8]_i_6 
       (.I0(\rgf_c0bus_wb[3]_i_7_4 ),
        .I1(\rgf_c0bus_wb[3]_i_7_2 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[8]_i_2 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[3]_i_7 ),
        .O(\badr[3]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h5050303F5F5F303F)) 
    \rgf_c0bus_wb[8]_i_7 
       (.I0(\rgf_c0bus_wb[3]_i_18 ),
        .I1(\rgf_c0bus_wb[3]_i_18_0 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[14]_i_13 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[14]_i_13_2 ),
        .O(\badr[8]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[9]_i_20 
       (.I0(\rgf_c0bus_wb[14]_i_13_5 ),
        .I1(\rgf_c0bus_wb[14]_i_13_0 ),
        .I2(\rgf_c0bus_wb[3]_i_7_0 ),
        .I3(\rgf_c0bus_wb[14]_i_13_6 ),
        .I4(\rgf_c0bus_wb[3]_i_7_1 ),
        .I5(\rgf_c0bus_wb[14]_i_13_4 ),
        .O(\badr[13]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c1bus_wb[12]_i_17 
       (.I0(\sr[4]_i_77_2 ),
        .I1(\sr[4]_i_77_0 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[4]_i_77 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[4]_i_77_1 ),
        .O(\badr[15]_INST_0_i_1_1 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c1bus_wb[12]_i_19 
       (.I0(\sr[6]_i_11_8 ),
        .I1(\sr[6]_i_11_9 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[6]_i_11 ),
        .O(\badr[6]_INST_0_i_1_1 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c1bus_wb[12]_i_20 
       (.I0(\sr[4]_i_99 ),
        .I1(\sr[4]_i_99_0 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[4]_i_99_1 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[4]_i_99_2 ),
        .O(\badr[10]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h03F3050503F3F5F5)) 
    \rgf_c1bus_wb[12]_i_21 
       (.I0(\sr[6]_i_11_3 ),
        .I1(\sr[6]_i_11_7 [2]),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_11_6 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[6]_i_11_5 ),
        .O(\sr_reg[6]_5 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[13]_i_6 
       (.I0(\badr[12]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb[14]_i_28_1 ),
        .O(\rgf_c1bus_wb[4]_i_9_0 ));
  LUT3 #(
    .INIT(8'hA3)) 
    \rgf_c1bus_wb[15]_i_15 
       (.I0(\badr[14]_INST_0_i_1_0 ),
        .I1(\badr[10]_INST_0_i_1 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[11]_i_10_4 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_18 
       (.I0(\sr[4]_i_77_1 ),
        .I1(\sr[4]_i_84 ),
        .O(\rgf_c1bus_wb[15]_i_27 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[15]_i_21 
       (.I0(\sr[6]_i_11_9 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_11_5 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[6]_i_11_8 ),
        .O(\badr[3]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[15]_i_22 
       (.I0(\sr[4]_i_99_0 ),
        .I1(\sr[4]_i_99_1 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_11 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[4]_i_99 ),
        .O(\badr[7]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[1]_i_13 
       (.I0(\sr[6]_i_11_8 ),
        .I1(\sr[6]_i_11_9 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_11_6 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[6]_i_11_5 ),
        .O(\badr[2]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[1]_i_14 
       (.I0(\sr[4]_i_99 ),
        .I1(\sr[4]_i_99_0 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[6]_i_11 ),
        .O(\badr[6]_INST_0_i_1_2 ));
  LUT6 #(
    .INIT(64'h3347FF47FFFFFFFF)) 
    \rgf_c1bus_wb[2]_i_6 
       (.I0(\sr[6]_i_11_5 ),
        .I1(\sr[6]_i_11_1 ),
        .I2(\sr[6]_i_11_6 ),
        .I3(\sr[6]_i_11_2 ),
        .I4(\sr[6]_i_11_3 ),
        .I5(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[11]_i_10_5 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \rgf_c1bus_wb[4]_i_18 
       (.I0(\sr[4]_i_175_0 ),
        .I1(\grn_reg[14] [4]),
        .I2(\sr[4]_i_179_1 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_175_1 ),
        .I5(\sr[4]_i_175_2 ),
        .O(\rgf_c1bus_wb[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \rgf_c1bus_wb[4]_i_19 
       (.I0(\sr[4]_i_175_3 ),
        .I1(\grn_reg[14] [2]),
        .I2(\sr[4]_i_175_4 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_175_5 ),
        .I5(\sr[4]_i_175_6 ),
        .O(\rgf_c1bus_wb[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_31 
       (.I0(\grn_reg[4]_4 ),
        .I1(\grn_reg[4]_5 ),
        .I2(\rgf_c1bus_wb[4]_i_25 ),
        .I3(\grn_reg[4]_9 ),
        .I4(a1buso2l_n_55),
        .I5(\rgf_c1bus_wb[4]_i_25_0 ),
        .O(\grn_reg[14] [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_35 
       (.I0(\grn_reg[2]_1 ),
        .I1(\grn_reg[2]_2 ),
        .I2(\sr[4]_i_211 ),
        .I3(\grn_reg[2]_5 ),
        .I4(a1buso2l_n_59),
        .I5(\sr[4]_i_211_0 ),
        .O(\grn_reg[14] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_39 
       (.I0(\grn_reg[15]_6 ),
        .I1(\grn_reg[15]_7 ),
        .I2(\rgf_c1bus_wb[4]_i_22 ),
        .I3(\grn_reg[15]_11 ),
        .I4(a1buso2l_n_34),
        .I5(\rgf_c1bus_wb[4]_i_22_0 ),
        .O(\grn_reg[15]_3 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_43 
       (.I0(\grn_reg[0]_2 ),
        .I1(\grn_reg[0]_3 ),
        .I2(\sr[4]_i_210 ),
        .I3(\grn_reg[0]_7 ),
        .I4(a1buso2l_n_63),
        .I5(\sr[4]_i_210_0 ),
        .O(\grn_reg[14] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_46 
       (.I0(\grn_reg[14]_2 ),
        .I1(\grn_reg[14]_3 ),
        .I2(\rgf_c1bus_wb[4]_i_23 ),
        .I3(\grn_reg[14]_6 ),
        .I4(a1buso2l_n_36),
        .I5(\rgf_c1bus_wb[4]_i_23_0 ),
        .O(\grn_reg[14] [12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_49 
       (.I0(\grn_reg[12]_1 ),
        .I1(\grn_reg[12]_2 ),
        .I2(\rgf_c1bus_wb[4]_i_24 ),
        .I3(\grn_reg[12]_5 ),
        .I4(a1buso2l_n_40),
        .I5(\rgf_c1bus_wb[4]_i_24_0 ),
        .O(\grn_reg[14] [10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_55 
       (.I0(\grn_reg[6]_1 ),
        .I1(\grn_reg[6]_2 ),
        .I2(\rgf_c1bus_wb[4]_i_26 ),
        .I3(\grn_reg[6]_5 ),
        .I4(a1buso2l_n_51),
        .I5(\rgf_c1bus_wb[4]_i_26_0 ),
        .O(\grn_reg[14] [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_59 
       (.I0(a1buso_n_30),
        .I1(a1buso_n_31),
        .I2(\rgf_c1bus_wb[4]_i_27 ),
        .I3(a1buso2l_n_23),
        .I4(a1buso2l_n_47),
        .I5(\rgf_c1bus_wb[4]_i_27_0 ),
        .O(\grn_reg[14] [6]));
  LUT6 #(
    .INIT(64'hF0FFF000AACCAACC)) 
    \rgf_c1bus_wb[4]_i_6 
       (.I0(\sr[6]_i_11_9 ),
        .I1(\sr[6]_i_11_8 ),
        .I2(\sr[6]_i_11_5 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[6]_i_11_6 ),
        .I5(\sr[6]_i_11_2 ),
        .O(\rgf_c1bus_wb[14]_i_28_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_63 
       (.I0(\grn_reg[10]_1 ),
        .I1(\grn_reg[10]_2 ),
        .I2(\rgf_c1bus_wb[4]_i_28 ),
        .I3(\grn_reg[10]_5 ),
        .I4(a1buso2l_n_44),
        .I5(\rgf_c1bus_wb[4]_i_28_0 ),
        .O(\grn_reg[14] [8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_66 
       (.I0(\grn_reg[1]_1 ),
        .I1(\grn_reg[1]_2 ),
        .I2(\sr[4]_i_213 ),
        .I3(\grn_reg[1]_5 ),
        .I4(a1buso2l_n_61),
        .I5(\sr[4]_i_213_0 ),
        .O(\grn_reg[14] [1]));
  LUT5 #(
    .INIT(32'h0FFF5533)) 
    \rgf_c1bus_wb[9]_i_17 
       (.I0(\sr[4]_i_77_0 ),
        .I1(\sr[4]_i_77 ),
        .I2(\sr[4]_i_77_1 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[6]_i_11_2 ),
        .O(\rgf_c1bus_wb[14]_i_28_3 ));
  LUT6 #(
    .INIT(64'h0F000FFFDDCCDDCC)) 
    \sr[4]_i_105 
       (.I0(\badr[15]_INST_0_i_1_1 ),
        .I1(\sr[4]_i_38 ),
        .I2(\rgf_c1bus_wb[14]_i_28_0 ),
        .I3(\rgf_c1bus_wb_reg[7] ),
        .I4(\rgf_c1bus_wb[14]_i_28 ),
        .I5(\rgf_c1bus_wb_reg[5]_1 ),
        .O(\rgf_c1bus_wb[15]_i_14_1 ));
  LUT6 #(
    .INIT(64'h555533330F0FFF00)) 
    \sr[4]_i_115 
       (.I0(\badr[3]_INST_0_i_1_0 ),
        .I1(\badr[7]_INST_0_i_1 ),
        .I2(\badr[11]_INST_0_i_1 ),
        .I3(\sr[4]_i_44 ),
        .I4(\rgf_c1bus_wb_reg[7] ),
        .I5(\rgf_c1bus_wb_reg[5]_1 ),
        .O(\rgf_c1bus_wb[15]_i_14_2 ));
  LUT6 #(
    .INIT(64'hF055FF55F033F033)) 
    \sr[4]_i_128 
       (.I0(\badr[10]_INST_0_i_2 ),
        .I1(\badr[6]_INST_0_i_2_0 ),
        .I2(\sr[4]_i_55 ),
        .I3(\rgf_c0bus_wb_reg[10]_0 ),
        .I4(\badr[2]_INST_0_i_2 ),
        .I5(\rgf_c0bus_wb_reg[10] ),
        .O(\rgf_c0bus_wb[11]_i_9 ));
  LUT5 #(
    .INIT(32'h5050303F)) 
    \sr[4]_i_135 
       (.I0(\badr[13]_INST_0_i_2_0 ),
        .I1(\badr[5]_INST_0_i_2_0 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\badr[9]_INST_0_i_2_0 ),
        .I4(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_11_2 ));
  LUT6 #(
    .INIT(64'h888888880F000FFF)) 
    \sr[4]_i_146 
       (.I0(\rgf_c0bus_wb[11]_i_9_0 ),
        .I1(\sr[4]_i_67 ),
        .I2(\badr[6]_INST_0_i_2_1 ),
        .I3(\rgf_c0bus_wb_reg[10] ),
        .I4(\badr[10]_INST_0_i_2_0 ),
        .I5(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_11_1 ));
  LUT6 #(
    .INIT(64'hCCAACCAA0F000FFF)) 
    \sr[4]_i_161 
       (.I0(\sr[4]_i_88 ),
        .I1(\sr[4]_i_88_0 ),
        .I2(\tr_reg[12]_0 ),
        .I3(\sr[6]_i_11_2 ),
        .I4(\tr_reg[14]_1 ),
        .I5(\rgf_c1bus_wb_reg[7] ),
        .O(\sr_reg[6]_6 ));
  LUT6 #(
    .INIT(64'hAFA0AFA0CFCFC0C0)) 
    \sr[4]_i_162 
       (.I0(\sr[4]_i_217_n_0 ),
        .I1(\sr[4]_i_218_n_0 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .I3(\rgf_c1bus_wb[4]_i_18_n_0 ),
        .I4(\sr[4]_i_219_n_0 ),
        .I5(\sr[6]_i_11_2 ),
        .O(\rgf_c1bus_wb[14]_i_28_6 ));
  LUT6 #(
    .INIT(64'h222EEE2EFFFFFFFF)) 
    \sr[4]_i_165 
       (.I0(\sr[4]_i_111 ),
        .I1(\sr[6]_i_11_2 ),
        .I2(\sr[6]_i_11_3 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[6]_i_11_6 ),
        .I5(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[11]_i_10_3 ));
  LUT6 #(
    .INIT(64'hCFCFAFA0C0C0AFA0)) 
    \sr[4]_i_169 
       (.I0(\tr_reg[12]_0 ),
        .I1(\sr[4]_i_218_n_0 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .I3(\sr[4]_i_217_n_0 ),
        .I4(\sr[6]_i_11_2 ),
        .I5(\sr[4]_i_219_n_0 ),
        .O(\sr[4]_i_219_0 ));
  LUT6 #(
    .INIT(64'h00000000222EEE2E)) 
    \sr[4]_i_173 
       (.I0(\sr[4]_i_102_0 ),
        .I1(\sr[6]_i_11_2 ),
        .I2(\sr[4]_i_99_2 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_102 ),
        .I5(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[11]_i_10_1 ));
  LUT6 #(
    .INIT(64'h3333555500FF0F0F)) 
    \sr[4]_i_175 
       (.I0(\sr[4]_i_217_n_0 ),
        .I1(\sr[4]_i_219_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_19_n_0 ),
        .I4(\sr[6]_i_11_2 ),
        .I5(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[11]_i_10_0 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \sr[4]_i_179 
       (.I0(\sr[4]_i_224_n_0 ),
        .I1(\sr[4]_i_225_n_0 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .I3(\sr[4]_i_88 ),
        .I4(\sr[6]_i_11_2 ),
        .I5(\sr[4]_i_111 ),
        .O(\sr[4]_i_220 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \sr[4]_i_180 
       (.I0(\tr_reg[12]_0 ),
        .I1(\tr_reg[14]_1 ),
        .I2(\sr[4]_i_217_n_0 ),
        .I3(\sr[6]_i_11_2 ),
        .I4(\sr[4]_i_218_n_0 ),
        .I5(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[11]_i_10_2 ));
  LUT6 #(
    .INIT(64'h3F3F505F3030505F)) 
    \sr[4]_i_181 
       (.I0(\sr[4]_i_219_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .I3(\rgf_c1bus_wb[4]_i_19_n_0 ),
        .I4(\sr[6]_i_11_2 ),
        .I5(\sr[4]_i_119 ),
        .O(\sr_reg[6]_11 ));
  LUT6 #(
    .INIT(64'h303F303FA0A0AFAF)) 
    \sr[4]_i_184 
       (.I0(\sr[4]_i_126 ),
        .I1(\sr_reg[14] ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_7_0 ),
        .O(\sr_reg[6]_24 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \sr[4]_i_196 
       (.I0(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\sr[4]_i_139 ),
        .I4(\rgf_c0bus_wb[3]_i_7_0 ),
        .I5(\rgf_c0bus_wb[12]_i_7 ),
        .O(\rgf_c0bus_wb[12]_i_24 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_203 
       (.I0(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I1(\sr_reg[14] ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_7_0 ),
        .I5(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_22_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_215 
       (.I0(\sr[4]_i_177 ),
        .I1(\grn_reg[14] [10]),
        .I2(\sr[4]_i_177_0 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_177_1 ),
        .I5(\sr[4]_i_177_2 ),
        .O(\tr_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_216 
       (.I0(\sr[4]_i_171 ),
        .I1(\grn_reg[14] [12]),
        .I2(\sr[4]_i_171_0 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_171_1 ),
        .I5(\sr[4]_i_171_2 ),
        .O(\tr_reg[14]_1 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_217 
       (.I0(\sr[4]_i_169_0 ),
        .I1(\grn_reg[14] [6]),
        .I2(\sr[4]_i_169_1 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_169_2 ),
        .I5(\sr[4]_i_179_0 ),
        .O(\sr[4]_i_217_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_218 
       (.I0(\sr[4]_i_169_3 ),
        .I1(\grn_reg[14] [8]),
        .I2(\sr[4]_i_169_4 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_169_5 ),
        .I5(\sr[4]_i_169_6 ),
        .O(\sr[4]_i_218_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_219 
       (.I0(\sr[4]_i_169_7 ),
        .I1(\grn_reg[14] [5]),
        .I2(\sr[4]_i_179_2 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_169_8 ),
        .I5(\sr[4]_i_179_3 ),
        .O(\sr[4]_i_219_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_224 
       (.I0(\sr[4]_i_179_4 ),
        .I1(a1bus_b02[5]),
        .I2(\sr[4]_i_179_3 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_179_5 ),
        .I5(\sr[4]_i_179_1 ),
        .O(\sr[4]_i_224_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_225 
       (.I0(\sr[4]_i_179_6 ),
        .I1(a1bus_b02[7]),
        .I2(\sr[4]_i_179_0 ),
        .I3(\sr[6]_i_11_1 ),
        .I4(\sr[4]_i_179_7 ),
        .I5(\sr[4]_i_179_2 ),
        .O(\sr[4]_i_225_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFFFEFFFE00)) 
    \sr[4]_i_226 
       (.I0(\rgf_c0bus_wb[4]_i_7 ),
        .I1(\sr[4]_i_188 ),
        .I2(\sr[4]_i_188_0 ),
        .I3(\rgf_c0bus_wb[3]_i_7_1 ),
        .I4(\sr[4]_i_188_1 ),
        .I5(\sr[4]_i_188_2 ),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_234 
       (.I0(\grn_reg[11]_1 ),
        .I1(\grn_reg[11]_2 ),
        .I2(\sr[4]_i_207 ),
        .I3(\grn_reg[11]_5 ),
        .I4(a1buso2l_n_42),
        .I5(\sr[4]_i_207_0 ),
        .O(\grn_reg[14] [9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_236 
       (.I0(\grn_reg[9]_1 ),
        .I1(\grn_reg[9]_2 ),
        .I2(\sr[4]_i_208 ),
        .I3(\grn_reg[9]_5 ),
        .I4(a1buso2l_n_46),
        .I5(\sr[4]_i_208_0 ),
        .O(\grn_reg[14] [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_238 
       (.I0(\grn_reg[13]_1 ),
        .I1(\grn_reg[13]_2 ),
        .I2(\sr[4]_i_209 ),
        .I3(\grn_reg[13]_5 ),
        .I4(a1buso2l_n_38),
        .I5(\sr[4]_i_209_0 ),
        .O(\grn_reg[14] [11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_241 
       (.I0(\grn_reg[3]_1 ),
        .I1(\grn_reg[3]_2 ),
        .I2(\sr[4]_i_220_0 ),
        .I3(\grn_reg[3]_5 ),
        .I4(a1buso2l_n_57),
        .I5(\sr[4]_i_220_1 ),
        .O(\grn_reg[14] [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_242 
       (.I0(\grn_reg[5]_1 ),
        .I1(\grn_reg[5]_2 ),
        .I2(\sr[4]_i_224_0 ),
        .I3(\grn_reg[5]_5 ),
        .I4(a1buso2l_n_53),
        .I5(\sr[4]_i_224_1 ),
        .O(a1bus_b02[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_244 
       (.I0(\grn_reg[7]_1 ),
        .I1(\grn_reg[7]_2 ),
        .I2(\sr[4]_i_225_0 ),
        .I3(\grn_reg[7]_5 ),
        .I4(a1buso2l_n_49),
        .I5(\sr[4]_i_225_1 ),
        .O(a1bus_b02[7]));
  LUT6 #(
    .INIT(64'h000000FF00004747)) 
    \sr[4]_i_89 
       (.I0(\badr[3]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\badr[7]_INST_0_i_1 ),
        .I3(\sr[4]_i_30_0 ),
        .I4(\rgf_c1bus_wb_reg[5] ),
        .I5(\rgf_c1bus_wb_reg[5]_1 ),
        .O(\rgf_c1bus_wb[15]_i_14_0 ));
  LUT6 #(
    .INIT(64'hAACCAACC0F0FFF0F)) 
    \sr[4]_i_91 
       (.I0(\badr[10]_INST_0_i_1 ),
        .I1(\badr[6]_INST_0_i_1_0 ),
        .I2(\sr[4]_i_30 ),
        .I3(\rgf_c1bus_wb_reg[7] ),
        .I4(\badr[2]_INST_0_i_1 ),
        .I5(\rgf_c1bus_wb_reg[5]_1 ),
        .O(\rgf_c1bus_wb[15]_i_14 ));
  LUT6 #(
    .INIT(64'h00000000AAAA303F)) 
    \sr[4]_i_94 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(\sr_reg[6]_1 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .I3(\badr[3]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb_reg[5] ),
        .I5(\rgf_c1bus_wb_reg[5]_1 ),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAA0CFC)) 
    \sr[6]_i_12 
       (.I0(\rgf_c0bus_wb[11]_i_8 ),
        .I1(\badr[4]_INST_0_i_2 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\sr[6]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb_reg[10]_0 ),
        .I5(\rgf_c0bus_wb[0]_i_14 ),
        .O(\rgf_c0bus_wb[15]_i_25_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_13 
       (.I0(\badr[8]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb_reg[10] ),
        .I2(\badr[3]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[8]_i_6_0 ));
  LUT6 #(
    .INIT(64'hFCFCFECECCCCFECE)) 
    \sr[6]_i_16 
       (.I0(\sr[6]_i_11_3 ),
        .I1(\sr[6]_i_11_4 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_11_5 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[6]_i_11_6 ),
        .O(\badr[1]_INST_0_i_1 ));
  LUT5 #(
    .INIT(32'hACAC0F00)) 
    \sr[6]_i_17 
       (.I0(\rgf_c0bus_wb[3]_i_7_2 ),
        .I1(\rgf_c0bus_wb[3]_i_7_4 ),
        .I2(\rgf_c0bus_wb[3]_i_7_1 ),
        .I3(\rgf_c0bus_wb[3]_i_7_3 ),
        .I4(\rgf_c0bus_wb[3]_i_7_0 ),
        .O(\sr[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0A0C0C0)) 
    \sr[6]_i_20 
       (.I0(\sr[4]_i_77 ),
        .I1(\sr[4]_i_77_0 ),
        .I2(\sr[6]_i_11_2 ),
        .I3(\sr[6]_i_15 ),
        .I4(\sr[6]_i_11_1 ),
        .I5(\sr[4]_i_77_1 ),
        .O(\stat_reg[2]_1 ));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_1__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[6] ),
        .I2(\sr[6]_i_11 ),
        .O(\badr[6]_INST_0_i_1_3 [1]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_2__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[5] ),
        .I2(\sr[6]_i_11_0 ),
        .O(\badr[6]_INST_0_i_1_3 [0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_5__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[7]_0 ),
        .I2(\sr[4]_i_99 ),
        .I3(\badr[6]_INST_0_i_1_3 [1]),
        .O(tout__1_carry__0_i_1__0_0[1]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_6__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[6] ),
        .I2(\sr[6]_i_11 ),
        .I3(\badr[6]_INST_0_i_1_3 [0]),
        .O(tout__1_carry__0_i_1__0_0[0]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_1__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[10] ),
        .I2(\sr[4]_i_99_2 ),
        .O(\badr[10]_INST_0_i_1_2 [3]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_2__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[9] ),
        .I2(\sr[4]_i_99_1 ),
        .O(\badr[10]_INST_0_i_1_2 [2]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_3__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[8] ),
        .I2(\sr[4]_i_99_0 ),
        .O(\badr[10]_INST_0_i_1_2 [1]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_4__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[7]_0 ),
        .I2(\sr[4]_i_99 ),
        .O(\badr[10]_INST_0_i_1_2 [0]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_5__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[11] ),
        .I2(\sr[4]_i_102 ),
        .I3(\badr[10]_INST_0_i_1_2 [3]),
        .O(tout__1_carry__1_i_1__0_0[3]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_6__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[10] ),
        .I2(\sr[4]_i_99_2 ),
        .I3(\badr[10]_INST_0_i_1_2 [2]),
        .O(tout__1_carry__1_i_1__0_0[2]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_7__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[9] ),
        .I2(\sr[4]_i_99_1 ),
        .I3(\badr[10]_INST_0_i_1_2 [1]),
        .O(tout__1_carry__1_i_1__0_0[1]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_8__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[8] ),
        .I2(\sr[4]_i_99_0 ),
        .I3(\badr[10]_INST_0_i_1_2 [0]),
        .O(tout__1_carry__1_i_1__0_0[0]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_2__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[13]_0 ),
        .I2(\sr[4]_i_77_0 ),
        .O(\badr[13]_INST_0_i_1_0 [2]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_3__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[12] ),
        .I2(\sr[4]_i_77_2 ),
        .O(\badr[13]_INST_0_i_1_0 [1]));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_4__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[11] ),
        .I2(\sr[4]_i_102 ),
        .O(\badr[13]_INST_0_i_1_0 [0]));
  LUT5 #(
    .INIT(32'hC33C5AA5)) 
    tout__1_carry__2_i_5
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[14]_0 ),
        .I2(tout__1_carry__2_0),
        .I3(\sr[4]_i_77_1 ),
        .I4(\sr[4]_i_77 ),
        .O(\badr[14]_INST_0_i_1_1 [3]));
  LUT6 #(
    .INIT(64'hF00F0FF0EE1111EE)) 
    tout__1_carry__2_i_5__0
       (.I0(\rgf_c0bus_wb[14]_i_2 ),
        .I1(tout__1_carry__2_1),
        .I2(\tr_reg[14] ),
        .I3(\tr_reg[15] ),
        .I4(\rgf_c0bus_wb[12]_i_10 ),
        .I5(\rgf_c0bus_wb[14]_i_13_6 ),
        .O(\badr[14]_INST_0_i_2_2 ));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_6
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[14]_0 ),
        .I2(\badr[13]_INST_0_i_1_0 [2]),
        .I3(\sr[4]_i_77 ),
        .O(\badr[14]_INST_0_i_1_1 [2]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_7__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[13]_0 ),
        .I2(\sr[4]_i_77_0 ),
        .I3(\badr[13]_INST_0_i_1_0 [1]),
        .O(\badr[14]_INST_0_i_1_1 [1]));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_8__0
       (.I0(tout__1_carry__2),
        .I1(\tr_reg[12] ),
        .I2(\sr[4]_i_77_2 ),
        .I3(\badr[13]_INST_0_i_1_0 [0]),
        .O(\badr[14]_INST_0_i_1_1 [0]));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank" *) 
module mcss_rgf_bank_5
   (.out({gr20[15],gr20[14],gr20[13],gr20[12],gr20[11],gr20[10],gr20[9],gr20[8],gr20[7],gr20[6],gr20[5],gr20[4],gr20[3],gr20[2],gr20[1],gr20[0]}),
    .\grn_reg[4] ({gr23[4],gr23[3],gr23[2],gr23[1],gr23[0]}),
    .\grn_reg[4]_0 ({gr24[4],gr24[3],gr24[2],gr24[1],gr24[0]}),
    .\grn_reg[15] ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_0 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[4]_1 ({gr27[4],gr27[3],gr27[2],gr27[1],gr27[0]}),
    .\grn_reg[15]_1 ({gr00[15],gr00[14],gr00[13],gr00[12],gr00[11],gr00[10],gr00[9],gr00[8],gr00[7],gr00[6],gr00[5],gr00[4],gr00[3],gr00[2],gr00[1],gr00[0]}),
    .\grn_reg[4]_2 ({gr03[4],gr03[3],gr03[2],gr03[1],gr03[0]}),
    .\grn_reg[4]_3 ({gr04[4],gr04[3],gr04[2],gr04[1],gr04[0]}),
    .\grn_reg[15]_2 ({gr05[15],gr05[14],gr05[13],gr05[12],gr05[11],gr05[10],gr05[9],gr05[8],gr05[7],gr05[6],gr05[5],gr05[4],gr05[3],gr05[2],gr05[1],gr05[0]}),
    .\grn_reg[15]_3 ({gr06[15],gr06[14],gr06[13],gr06[12],gr06[11],gr06[10],gr06[9],gr06[8],gr06[7],gr06[6],gr06[5],gr06[4],gr06[3],gr06[2],gr06[1],gr06[0]}),
    .\grn_reg[4]_4 ({gr07[4],gr07[3],gr07[2],gr07[1],gr07[0]}),
    SR,
    \sr[4]_i_156_0 ,
    \tr_reg[11] ,
    \tr_reg[13] ,
    \sr_reg[6] ,
    \badr[15]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_28 ,
    \sr_reg[6]_0 ,
    \rgf_c1bus_wb[4]_i_28_0 ,
    \tr_reg[12] ,
    \tr_reg[1] ,
    \tr_reg[3] ,
    \tr_reg[13]_0 ,
    \tr_reg[1]_0 ,
    \tr_reg[14] ,
    \sr[4]_i_133_0 ,
    \rgf_c0bus_wb[4]_i_26_0 ,
    \sr[4]_i_200_0 ,
    \sr[4]_i_195_0 ,
    \rgf_c0bus_wb[4]_i_32_0 ,
    \rgf_c0bus_wb[13]_i_27_0 ,
    \sr_reg[6]_1 ,
    \sr_reg[6]_2 ,
    \sp_reg[2] ,
    \rgf_c0bus_wb[13]_i_30_0 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    \sp_reg[13] ,
    \sp_reg[11] ,
    \rgf_c0bus_wb[4]_i_29_0 ,
    \sp_reg[14] ,
    \rgf_c0bus_wb[4]_i_33_0 ,
    \rgf_c0bus_wb[4]_i_31_0 ,
    \sr[4]_i_232_0 ,
    \sp_reg[1] ,
    \sr_reg[6]_5 ,
    \sp_reg[4] ,
    \badr[15]_INST_0_i_2 ,
    \sp_reg[6] ,
    \fdatx[15] ,
    .fdat_12_sp_1(fdat_12_sn_1),
    \fdat[15] ,
    \grn_reg[15]_4 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4]_5 ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_5 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_6 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[15]_7 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_8 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[15]_8 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_9 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_9 ,
    gr6_bus1,
    \grn_reg[15]_10 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_11 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[8]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_11 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_6 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[8]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_12 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_7 ,
    \grn_reg[4]_13 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_8 ,
    p_0_in,
    \grn_reg[15]_12 ,
    \grn_reg[14]_7 ,
    \grn_reg[13]_7 ,
    \grn_reg[12]_7 ,
    \grn_reg[11]_7 ,
    \grn_reg[10]_7 ,
    \grn_reg[9]_7 ,
    \grn_reg[8]_7 ,
    \grn_reg[7]_7 ,
    \grn_reg[6]_7 ,
    \grn_reg[5]_7 ,
    \grn_reg[4]_14 ,
    \grn_reg[3]_8 ,
    \grn_reg[2]_8 ,
    \grn_reg[1]_8 ,
    \grn_reg[0]_9 ,
    \grn_reg[15]_13 ,
    \grn_reg[14]_8 ,
    \grn_reg[13]_8 ,
    \grn_reg[12]_8 ,
    \grn_reg[11]_8 ,
    \grn_reg[10]_8 ,
    \grn_reg[9]_8 ,
    \grn_reg[8]_8 ,
    \grn_reg[7]_8 ,
    \grn_reg[6]_8 ,
    \grn_reg[5]_8 ,
    \grn_reg[4]_15 ,
    \grn_reg[3]_9 ,
    \grn_reg[2]_9 ,
    \grn_reg[1]_9 ,
    \grn_reg[0]_10 ,
    \grn_reg[15]_14 ,
    \grn_reg[14]_9 ,
    \grn_reg[13]_9 ,
    \grn_reg[12]_9 ,
    \grn_reg[11]_9 ,
    \grn_reg[10]_9 ,
    \grn_reg[9]_9 ,
    \grn_reg[8]_9 ,
    \grn_reg[7]_9 ,
    \grn_reg[6]_9 ,
    \grn_reg[5]_9 ,
    \grn_reg[4]_16 ,
    \grn_reg[3]_10 ,
    \grn_reg[2]_10 ,
    \grn_reg[1]_10 ,
    \grn_reg[0]_11 ,
    \grn_reg[15]_15 ,
    \grn_reg[14]_10 ,
    \grn_reg[13]_10 ,
    \grn_reg[12]_10 ,
    \grn_reg[11]_10 ,
    \grn_reg[10]_10 ,
    \grn_reg[9]_10 ,
    \grn_reg[8]_10 ,
    \grn_reg[7]_10 ,
    \grn_reg[6]_10 ,
    \grn_reg[5]_10 ,
    \grn_reg[4]_17 ,
    \grn_reg[3]_11 ,
    \grn_reg[2]_11 ,
    \grn_reg[1]_11 ,
    \grn_reg[0]_12 ,
    \grn_reg[15]_16 ,
    gr6_bus1_0,
    \grn_reg[14]_11 ,
    \grn_reg[13]_11 ,
    \grn_reg[12]_11 ,
    \grn_reg[11]_11 ,
    \grn_reg[10]_11 ,
    \grn_reg[9]_11 ,
    \grn_reg[8]_11 ,
    \grn_reg[7]_11 ,
    \grn_reg[6]_11 ,
    \grn_reg[5]_11 ,
    \grn_reg[4]_18 ,
    \grn_reg[3]_12 ,
    \grn_reg[2]_12 ,
    \grn_reg[1]_12 ,
    \grn_reg[0]_13 ,
    \grn_reg[15]_17 ,
    \grn_reg[14]_12 ,
    \grn_reg[13]_12 ,
    \grn_reg[12]_12 ,
    \grn_reg[11]_12 ,
    \grn_reg[10]_12 ,
    \grn_reg[9]_12 ,
    \grn_reg[8]_12 ,
    \grn_reg[7]_12 ,
    \grn_reg[6]_12 ,
    \grn_reg[5]_12 ,
    \grn_reg[4]_19 ,
    \grn_reg[3]_13 ,
    \grn_reg[2]_13 ,
    \grn_reg[1]_13 ,
    \grn_reg[0]_14 ,
    \grn_reg[15]_18 ,
    \grn_reg[14]_13 ,
    \grn_reg[13]_13 ,
    \grn_reg[12]_13 ,
    \grn_reg[11]_13 ,
    \grn_reg[10]_13 ,
    \grn_reg[9]_13 ,
    \grn_reg[8]_13 ,
    \grn_reg[7]_13 ,
    \grn_reg[6]_13 ,
    \grn_reg[5]_13 ,
    \grn_reg[4]_20 ,
    \grn_reg[3]_14 ,
    \grn_reg[2]_14 ,
    \grn_reg[1]_14 ,
    \grn_reg[0]_15 ,
    \grn_reg[14]_14 ,
    \grn_reg[13]_14 ,
    \grn_reg[12]_14 ,
    \grn_reg[11]_14 ,
    \grn_reg[10]_14 ,
    \grn_reg[9]_14 ,
    \grn_reg[8]_14 ,
    \grn_reg[7]_14 ,
    \grn_reg[6]_14 ,
    \grn_reg[5]_14 ,
    \grn_reg[4]_21 ,
    \grn_reg[3]_15 ,
    \grn_reg[2]_15 ,
    \grn_reg[1]_15 ,
    \grn_reg[0]_16 ,
    a1bus_b13,
    rst_n,
    \sr[4]_i_27 ,
    \sr[4]_i_27_0 ,
    \sr[4]_i_27_1 ,
    \sr[4]_i_80_0 ,
    \sr[4]_i_80_1 ,
    \sr[4]_i_80_2 ,
    \sr[4]_i_83 ,
    \sr[4]_i_90 ,
    \sr[4]_i_164_0 ,
    \rgf_c1bus_wb[4]_i_11 ,
    \sr[4]_i_170 ,
    \sr[4]_i_170_0 ,
    \sr[4]_i_164_1 ,
    \sr[4]_i_170_1 ,
    \sr[4]_i_155_0 ,
    \sr[4]_i_170_2 ,
    \sr[4]_i_155_1 ,
    \sr[4]_i_170_3 ,
    \rgf_c1bus_wb[4]_i_11_0 ,
    \sr[4]_i_168 ,
    \rgf_c1bus_wb[4]_i_11_1 ,
    \sr[4]_i_168_0 ,
    \sr[4]_i_168_1 ,
    \sr[4]_i_168_2 ,
    \sr[4]_i_159_0 ,
    \sr[4]_i_168_3 ,
    \sr[4]_i_159_1 ,
    \sr[4]_i_154_0 ,
    \sr[4]_i_159_2 ,
    \sr[4]_i_154_1 ,
    \rgf_c1bus_wb[4]_i_11_2 ,
    \rgf_c1bus_wb[4]_i_11_3 ,
    \rgf_c1bus_wb[4]_i_11_4 ,
    \sr[4]_i_155_2 ,
    \sr[4]_i_155_3 ,
    \sr[4]_i_155_4 ,
    \sr[4]_i_155_5 ,
    \sr[4]_i_155_6 ,
    \sr[4]_i_155_7 ,
    \sr[4]_i_164_2 ,
    \sr[4]_i_164_3 ,
    \sr[4]_i_159_3 ,
    \sr[4]_i_159_4 ,
    \sr[4]_i_159_5 ,
    \sr[4]_i_155_8 ,
    \sr[4]_i_155_9 ,
    \sr[4]_i_155_10 ,
    \sr[4]_i_155_11 ,
    \rgf_c1bus_wb[4]_i_11_5 ,
    \rgf_c1bus_wb[4]_i_11_6 ,
    \sr[4]_i_159_6 ,
    \sr[4]_i_159_7 ,
    \sr[4]_i_15 ,
    \sr[4]_i_15_0 ,
    \sr[4]_i_15_1 ,
    \sr[4]_i_57_0 ,
    \sr[4]_i_57_1 ,
    \sr[4]_i_57_2 ,
    \sr[4]_i_66 ,
    \sr[4]_i_66_0 ,
    \sr[4]_i_57_3 ,
    \sr[4]_i_67 ,
    \sr[4]_i_67_0 ,
    \sr[4]_i_139 ,
    \sr[4]_i_139_0 ,
    \rgf_c0bus_wb[12]_i_7 ,
    \sr[4]_i_138_0 ,
    \sr[4]_i_138_1 ,
    \rgf_c0bus_wb[13]_i_13 ,
    \sr[4]_i_129 ,
    \sr[4]_i_197_0 ,
    \sr[4]_i_197_1 ,
    \sr[4]_i_197_2 ,
    \sr[4]_i_185 ,
    \sr[4]_i_185_0 ,
    \rgf_c0bus_wb[4]_i_12 ,
    \rgf_c0bus_wb[15]_i_23_0 ,
    \rgf_c0bus_wb[15]_i_23_1 ,
    \sr[4]_i_183_0 ,
    \rgf_c0bus_wb[15]_i_23_2 ,
    \sr[4]_i_183_1 ,
    \sr[4]_i_186_0 ,
    \sr[4]_i_186_1 ,
    \sr[4]_i_183_2 ,
    \rgf_c0bus_wb[15]_i_23_3 ,
    \sr[4]_i_183_3 ,
    \sr[4]_i_197_3 ,
    \sr[4]_i_197_4 ,
    \sr[4]_i_183_4 ,
    \sr[4]_i_197_5 ,
    \rgf_c0bus_wb[15]_i_23_4 ,
    \rgf_c0bus_wb[15]_i_23_5 ,
    \sr[4]_i_183_5 ,
    \rgf_c0bus_wb[15]_i_23_6 ,
    \sr[4]_i_183_6 ,
    \sr[4]_i_183_7 ,
    \sr[4]_i_183_8 ,
    \sr[4]_i_183_9 ,
    \sr[4]_i_183_10 ,
    \sr[4]_i_183_11 ,
    \sr[4]_i_183_12 ,
    \sr[4]_i_183_13 ,
    \sr[4]_i_183_14 ,
    \sr[4]_i_183_15 ,
    \rgf_c0bus_wb[4]_i_8_0 ,
    \rgf_c0bus_wb[4]_i_8_1 ,
    \sr[4]_i_183_16 ,
    \sr[4]_i_183_17 ,
    \sr[4]_i_183_18 ,
    \rgf_c0bus_wb[4]_i_8_2 ,
    \rgf_c0bus_wb[4]_i_8_3 ,
    \rgf_c0bus_wb[4]_i_8_4 ,
    \sr[4]_i_197_6 ,
    \sr[4]_i_197_7 ,
    \rgf_c0bus_wb[4]_i_8_5 ,
    \rgf_c0bus_wb[4]_i_8_6 ,
    \rgf_c0bus_wb[4]_i_8_7 ,
    \rgf_c0bus_wb[4]_i_8_8 ,
    \rgf_c0bus_wb[4]_i_8_9 ,
    \rgf_c0bus_wb[4]_i_12_0 ,
    \rgf_c0bus_wb[4]_i_12_1 ,
    \rgf_c0bus_wb[4]_i_12_2 ,
    \rgf_c0bus_wb[15]_i_23_7 ,
    \sr[4]_i_186_2 ,
    \sr[4]_i_186_3 ,
    \sr[4]_i_186_4 ,
    \sr[4]_i_186_5 ,
    \sr[4]_i_194_0 ,
    \sr[4]_i_194_1 ,
    \sr[4]_i_194_2 ,
    \sr[4]_i_194_3 ,
    \sr[4]_i_194_4 ,
    \sr[4]_i_194_5 ,
    \rgf_c0bus_wb[15]_i_23_8 ,
    \rgf_c0bus_wb[15]_i_23_9 ,
    \sr[4]_i_183_19 ,
    fdatx,
    \ir0_id_fl[20]_i_4 ,
    fdat,
    \nir_id_reg[20] ,
    a0bus_sel_0,
    \i_/badr[15]_INST_0_i_135 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_135_0 ,
    ctl_sela0,
    \i_/badr[15]_INST_0_i_135_1 ,
    \bbus_o[4]_INST_0_i_7 ,
    \bbus_o[4]_INST_0_i_7_0 ,
    \bbus_o[3]_INST_0_i_7 ,
    \bbus_o[3]_INST_0_i_7_0 ,
    \bbus_o[2]_INST_0_i_7 ,
    \bbus_o[2]_INST_0_i_7_0 ,
    \bbus_o[1]_INST_0_i_7 ,
    \bbus_o[1]_INST_0_i_7_0 ,
    \bbus_o[0]_INST_0_i_7 ,
    \bbus_o[0]_INST_0_i_7_0 ,
    \i_/bdatw[15]_INST_0_i_34 ,
    \i_/bbus_o[4]_INST_0_i_20 ,
    \i_/bbus_o[4]_INST_0_i_21 ,
    \i_/bbus_o[4]_INST_0_i_21_0 ,
    ctl_selb0_0,
    \bbus_o[4]_INST_0_i_7_1 ,
    \bbus_o[4]_INST_0_i_7_2 ,
    \bbus_o[3]_INST_0_i_7_1 ,
    \bbus_o[3]_INST_0_i_7_2 ,
    \bbus_o[2]_INST_0_i_7_1 ,
    \bbus_o[2]_INST_0_i_7_2 ,
    \bbus_o[1]_INST_0_i_7_1 ,
    \bbus_o[1]_INST_0_i_7_2 ,
    \bbus_o[0]_INST_0_i_7_1 ,
    \bbus_o[0]_INST_0_i_7_2 ,
    \i_/bdatw[15]_INST_0_i_92 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_34_0 ,
    b0bus_sel_0,
    \i_/bbus_o[4]_INST_0_i_20_0 ,
    \i_/bbus_o[4]_INST_0_i_20_1 ,
    \i_/bdatw[15]_INST_0_i_33 ,
    \i_/bbus_o[4]_INST_0_i_21_1 ,
    \i_/badr[0]_INST_0_i_18 ,
    \i_/badr[0]_INST_0_i_18_0 ,
    \i_/badr[0]_INST_0_i_18_1 ,
    \rgf_c1bus_wb[4]_i_40 ,
    \rgf_c1bus_wb[4]_i_40_0 ,
    \rgf_c1bus_wb[4]_i_42 ,
    \rgf_c1bus_wb[4]_i_42_0 ,
    \rgf_c1bus_wb[4]_i_50 ,
    \rgf_c1bus_wb[4]_i_50_0 ,
    \rgf_c1bus_wb[4]_i_48 ,
    \rgf_c1bus_wb[4]_i_48_0 ,
    \rgf_c1bus_wb[4]_i_64 ,
    \rgf_c1bus_wb[4]_i_64_0 ,
    \rgf_c1bus_wb[4]_i_62 ,
    \rgf_c1bus_wb[4]_i_62_0 ,
    \rgf_c1bus_wb[4]_i_60 ,
    \rgf_c1bus_wb[4]_i_60_0 ,
    \rgf_c1bus_wb[4]_i_58 ,
    \rgf_c1bus_wb[4]_i_58_0 ,
    \rgf_c1bus_wb[4]_i_56 ,
    \rgf_c1bus_wb[4]_i_56_0 ,
    \rgf_c1bus_wb[4]_i_54 ,
    \rgf_c1bus_wb[4]_i_54_0 ,
    \rgf_c1bus_wb[4]_i_52 ,
    \rgf_c1bus_wb[4]_i_52_0 ,
    \rgf_c1bus_wb[4]_i_32 ,
    \rgf_c1bus_wb[4]_i_32_0 ,
    \rgf_c1bus_wb[4]_i_34 ,
    \rgf_c1bus_wb[4]_i_34_0 ,
    \rgf_c1bus_wb[4]_i_36 ,
    \rgf_c1bus_wb[4]_i_36_0 ,
    \rgf_c1bus_wb[4]_i_38 ,
    \rgf_c1bus_wb[4]_i_38_0 ,
    \sr[4]_i_239 ,
    \sr[4]_i_239_0 ,
    a1bus_sel_0,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_212 ,
    \i_/bdatw[15]_INST_0_i_124 ,
    \i_/bdatw[15]_INST_0_i_121 ,
    \i_/bdatw[15]_INST_0_i_121_0 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_121_1 ,
    \i_/badr[15]_INST_0_i_52 ,
    \bbus_o[4]_INST_0_i_7_3 ,
    \bbus_o[4]_INST_0_i_7_4 ,
    \bbus_o[3]_INST_0_i_7_3 ,
    \bbus_o[3]_INST_0_i_7_4 ,
    \bbus_o[2]_INST_0_i_7_3 ,
    \bbus_o[2]_INST_0_i_7_4 ,
    \bbus_o[1]_INST_0_i_7_3 ,
    \bbus_o[1]_INST_0_i_7_4 ,
    \bbus_o[0]_INST_0_i_7_3 ,
    \bbus_o[0]_INST_0_i_7_4 ,
    \bbus_o[4]_INST_0_i_7_5 ,
    \bbus_o[4]_INST_0_i_7_6 ,
    \bbus_o[3]_INST_0_i_7_5 ,
    \bbus_o[3]_INST_0_i_7_6 ,
    \bbus_o[2]_INST_0_i_7_5 ,
    \bbus_o[2]_INST_0_i_7_6 ,
    \bbus_o[1]_INST_0_i_7_5 ,
    \bbus_o[1]_INST_0_i_7_6 ,
    \bbus_o[0]_INST_0_i_7_5 ,
    \bbus_o[0]_INST_0_i_7_6 ,
    \rgf_c1bus_wb[4]_i_45 ,
    \rgf_c1bus_wb[4]_i_45_0 ,
    \rgf_c1bus_wb[4]_i_42_1 ,
    \rgf_c1bus_wb[4]_i_42_2 ,
    \rgf_c1bus_wb[4]_i_50_1 ,
    \rgf_c1bus_wb[4]_i_50_2 ,
    \rgf_c1bus_wb[4]_i_48_1 ,
    \rgf_c1bus_wb[4]_i_48_2 ,
    \rgf_c1bus_wb[4]_i_64_1 ,
    \rgf_c1bus_wb[4]_i_64_2 ,
    \rgf_c1bus_wb[4]_i_62_1 ,
    \rgf_c1bus_wb[4]_i_62_2 ,
    \rgf_c1bus_wb[4]_i_60_1 ,
    \rgf_c1bus_wb[4]_i_60_2 ,
    \rgf_c1bus_wb[4]_i_58_1 ,
    \rgf_c1bus_wb[4]_i_58_2 ,
    \rgf_c1bus_wb[4]_i_56_1 ,
    \rgf_c1bus_wb[4]_i_56_2 ,
    \rgf_c1bus_wb[4]_i_54_1 ,
    \rgf_c1bus_wb[4]_i_54_2 ,
    \rgf_c1bus_wb[4]_i_52_1 ,
    \rgf_c1bus_wb[4]_i_52_2 ,
    \rgf_c1bus_wb[4]_i_32_1 ,
    \rgf_c1bus_wb[4]_i_32_2 ,
    \rgf_c1bus_wb[4]_i_34_1 ,
    \rgf_c1bus_wb[4]_i_34_2 ,
    \rgf_c1bus_wb[4]_i_36_1 ,
    \rgf_c1bus_wb[4]_i_36_2 ,
    \rgf_c1bus_wb[4]_i_38_1 ,
    \rgf_c1bus_wb[4]_i_38_2 ,
    \rgf_c1bus_wb[4]_i_44 ,
    \rgf_c1bus_wb[4]_i_44_0 ,
    \bdatw[12]_INST_0_i_42 ,
    \bdatw[12]_INST_0_i_42_0 ,
    \bdatw[11]_INST_0_i_44 ,
    \bdatw[11]_INST_0_i_44_0 ,
    \bdatw[10]_INST_0_i_43 ,
    \bdatw[10]_INST_0_i_43_0 ,
    \bdatw[9]_INST_0_i_42 ,
    \bdatw[9]_INST_0_i_42_0 ,
    \bdatw[8]_INST_0_i_43 ,
    \bdatw[8]_INST_0_i_43_0 ,
    \badr[15]_INST_0_i_1_0 ,
    \badr[15]_INST_0_i_1_1 ,
    \badr[14]_INST_0_i_1 ,
    \badr[14]_INST_0_i_1_0 ,
    \badr[13]_INST_0_i_1 ,
    \badr[13]_INST_0_i_1_0 ,
    \badr[12]_INST_0_i_1 ,
    \badr[12]_INST_0_i_1_0 ,
    \badr[11]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1_0 ,
    \badr[10]_INST_0_i_1 ,
    \badr[10]_INST_0_i_1_0 ,
    \badr[9]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1_0 ,
    \badr[8]_INST_0_i_1 ,
    \badr[8]_INST_0_i_1_0 ,
    \badr[7]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1_0 ,
    \badr[6]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1_0 ,
    \badr[5]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1_0 ,
    \badr[4]_INST_0_i_1 ,
    \badr[4]_INST_0_i_1_0 ,
    \badr[3]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1_0 ,
    \badr[2]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1_0 ,
    \badr[1]_INST_0_i_1 ,
    \badr[1]_INST_0_i_1_0 ,
    \badr[0]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1_0 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    clk,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 ,
    \grn_reg[15]_25 ,
    \grn_reg[15]_26 ,
    \grn_reg[15]_27 ,
    \grn_reg[15]_28 ,
    \grn_reg[15]_29 ,
    \grn_reg[15]_30 ,
    \grn_reg[15]_31 ,
    \grn_reg[15]_32 ,
    \grn_reg[15]_33 ,
    \grn_reg[15]_34 ,
    \grn_reg[15]_35 ,
    \grn_reg[15]_36 ,
    \grn_reg[15]_37 ,
    \grn_reg[15]_38 ,
    \grn_reg[15]_39 ,
    \grn_reg[15]_40 ,
    \grn_reg[15]_41 ,
    \grn_reg[15]_42 ,
    \grn_reg[15]_43 ,
    \grn_reg[15]_44 ,
    \grn_reg[15]_45 ,
    \grn_reg[15]_46 ,
    \grn_reg[15]_47 ,
    \grn_reg[15]_48 ,
    \grn_reg[15]_49 ,
    \grn_reg[15]_50 );
  output [0:0]SR;
  output \sr[4]_i_156_0 ;
  output \tr_reg[11] ;
  output \tr_reg[13] ;
  output \sr_reg[6] ;
  output \badr[15]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_28 ;
  output \sr_reg[6]_0 ;
  output \rgf_c1bus_wb[4]_i_28_0 ;
  output \tr_reg[12] ;
  output \tr_reg[1] ;
  output \tr_reg[3] ;
  output \tr_reg[13]_0 ;
  output \tr_reg[1]_0 ;
  output \tr_reg[14] ;
  output \sr[4]_i_133_0 ;
  output \rgf_c0bus_wb[4]_i_26_0 ;
  output \sr[4]_i_200_0 ;
  output \sr[4]_i_195_0 ;
  output \rgf_c0bus_wb[4]_i_32_0 ;
  output \rgf_c0bus_wb[13]_i_27_0 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[6]_2 ;
  output \sp_reg[2] ;
  output \rgf_c0bus_wb[13]_i_30_0 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[6]_4 ;
  output \sp_reg[13] ;
  output \sp_reg[11] ;
  output \rgf_c0bus_wb[4]_i_29_0 ;
  output \sp_reg[14] ;
  output \rgf_c0bus_wb[4]_i_33_0 ;
  output \rgf_c0bus_wb[4]_i_31_0 ;
  output \sr[4]_i_232_0 ;
  output \sp_reg[1] ;
  output \sr_reg[6]_5 ;
  output \sp_reg[4] ;
  output \badr[15]_INST_0_i_2 ;
  output \sp_reg[6] ;
  output \fdatx[15] ;
  output [0:0]\fdat[15] ;
  output \grn_reg[15]_4 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_5 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_6 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_8 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_9 ;
  output gr6_bus1;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[8]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_11 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_6 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[8]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_12 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_7 ;
  output \grn_reg[4]_13 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_8 ;
  output [15:0]p_0_in;
  output \grn_reg[15]_12 ;
  output \grn_reg[14]_7 ;
  output \grn_reg[13]_7 ;
  output \grn_reg[12]_7 ;
  output \grn_reg[11]_7 ;
  output \grn_reg[10]_7 ;
  output \grn_reg[9]_7 ;
  output \grn_reg[8]_7 ;
  output \grn_reg[7]_7 ;
  output \grn_reg[6]_7 ;
  output \grn_reg[5]_7 ;
  output \grn_reg[4]_14 ;
  output \grn_reg[3]_8 ;
  output \grn_reg[2]_8 ;
  output \grn_reg[1]_8 ;
  output \grn_reg[0]_9 ;
  output \grn_reg[15]_13 ;
  output \grn_reg[14]_8 ;
  output \grn_reg[13]_8 ;
  output \grn_reg[12]_8 ;
  output \grn_reg[11]_8 ;
  output \grn_reg[10]_8 ;
  output \grn_reg[9]_8 ;
  output \grn_reg[8]_8 ;
  output \grn_reg[7]_8 ;
  output \grn_reg[6]_8 ;
  output \grn_reg[5]_8 ;
  output \grn_reg[4]_15 ;
  output \grn_reg[3]_9 ;
  output \grn_reg[2]_9 ;
  output \grn_reg[1]_9 ;
  output \grn_reg[0]_10 ;
  output \grn_reg[15]_14 ;
  output \grn_reg[14]_9 ;
  output \grn_reg[13]_9 ;
  output \grn_reg[12]_9 ;
  output \grn_reg[11]_9 ;
  output \grn_reg[10]_9 ;
  output \grn_reg[9]_9 ;
  output \grn_reg[8]_9 ;
  output \grn_reg[7]_9 ;
  output \grn_reg[6]_9 ;
  output \grn_reg[5]_9 ;
  output \grn_reg[4]_16 ;
  output \grn_reg[3]_10 ;
  output \grn_reg[2]_10 ;
  output \grn_reg[1]_10 ;
  output \grn_reg[0]_11 ;
  output \grn_reg[15]_15 ;
  output \grn_reg[14]_10 ;
  output \grn_reg[13]_10 ;
  output \grn_reg[12]_10 ;
  output \grn_reg[11]_10 ;
  output \grn_reg[10]_10 ;
  output \grn_reg[9]_10 ;
  output \grn_reg[8]_10 ;
  output \grn_reg[7]_10 ;
  output \grn_reg[6]_10 ;
  output \grn_reg[5]_10 ;
  output \grn_reg[4]_17 ;
  output \grn_reg[3]_11 ;
  output \grn_reg[2]_11 ;
  output \grn_reg[1]_11 ;
  output \grn_reg[0]_12 ;
  output \grn_reg[15]_16 ;
  output gr6_bus1_0;
  output \grn_reg[14]_11 ;
  output \grn_reg[13]_11 ;
  output \grn_reg[12]_11 ;
  output \grn_reg[11]_11 ;
  output \grn_reg[10]_11 ;
  output \grn_reg[9]_11 ;
  output \grn_reg[8]_11 ;
  output \grn_reg[7]_11 ;
  output \grn_reg[6]_11 ;
  output \grn_reg[5]_11 ;
  output \grn_reg[4]_18 ;
  output \grn_reg[3]_12 ;
  output \grn_reg[2]_12 ;
  output \grn_reg[1]_12 ;
  output \grn_reg[0]_13 ;
  output \grn_reg[15]_17 ;
  output \grn_reg[14]_12 ;
  output \grn_reg[13]_12 ;
  output \grn_reg[12]_12 ;
  output \grn_reg[11]_12 ;
  output \grn_reg[10]_12 ;
  output \grn_reg[9]_12 ;
  output \grn_reg[8]_12 ;
  output \grn_reg[7]_12 ;
  output \grn_reg[6]_12 ;
  output \grn_reg[5]_12 ;
  output \grn_reg[4]_19 ;
  output \grn_reg[3]_13 ;
  output \grn_reg[2]_13 ;
  output \grn_reg[1]_13 ;
  output \grn_reg[0]_14 ;
  output \grn_reg[15]_18 ;
  output \grn_reg[14]_13 ;
  output \grn_reg[13]_13 ;
  output \grn_reg[12]_13 ;
  output \grn_reg[11]_13 ;
  output \grn_reg[10]_13 ;
  output \grn_reg[9]_13 ;
  output \grn_reg[8]_13 ;
  output \grn_reg[7]_13 ;
  output \grn_reg[6]_13 ;
  output \grn_reg[5]_13 ;
  output \grn_reg[4]_20 ;
  output \grn_reg[3]_14 ;
  output \grn_reg[2]_14 ;
  output \grn_reg[1]_14 ;
  output \grn_reg[0]_15 ;
  output \grn_reg[14]_14 ;
  output \grn_reg[13]_14 ;
  output \grn_reg[12]_14 ;
  output \grn_reg[11]_14 ;
  output \grn_reg[10]_14 ;
  output \grn_reg[9]_14 ;
  output \grn_reg[8]_14 ;
  output \grn_reg[7]_14 ;
  output \grn_reg[6]_14 ;
  output \grn_reg[5]_14 ;
  output \grn_reg[4]_21 ;
  output \grn_reg[3]_15 ;
  output \grn_reg[2]_15 ;
  output \grn_reg[1]_15 ;
  output \grn_reg[0]_16 ;
  output [15:0]a1bus_b13;
  input rst_n;
  input \sr[4]_i_27 ;
  input \sr[4]_i_27_0 ;
  input \sr[4]_i_27_1 ;
  input \sr[4]_i_80_0 ;
  input \sr[4]_i_80_1 ;
  input \sr[4]_i_80_2 ;
  input \sr[4]_i_83 ;
  input \sr[4]_i_90 ;
  input \sr[4]_i_164_0 ;
  input [12:0]\rgf_c1bus_wb[4]_i_11 ;
  input \sr[4]_i_170 ;
  input \sr[4]_i_170_0 ;
  input \sr[4]_i_164_1 ;
  input \sr[4]_i_170_1 ;
  input \sr[4]_i_155_0 ;
  input \sr[4]_i_170_2 ;
  input \sr[4]_i_155_1 ;
  input \sr[4]_i_170_3 ;
  input \rgf_c1bus_wb[4]_i_11_0 ;
  input \sr[4]_i_168 ;
  input \rgf_c1bus_wb[4]_i_11_1 ;
  input \sr[4]_i_168_0 ;
  input \sr[4]_i_168_1 ;
  input \sr[4]_i_168_2 ;
  input \sr[4]_i_159_0 ;
  input \sr[4]_i_168_3 ;
  input \sr[4]_i_159_1 ;
  input \sr[4]_i_154_0 ;
  input \sr[4]_i_159_2 ;
  input \sr[4]_i_154_1 ;
  input \rgf_c1bus_wb[4]_i_11_2 ;
  input \rgf_c1bus_wb[4]_i_11_3 ;
  input \rgf_c1bus_wb[4]_i_11_4 ;
  input \sr[4]_i_155_2 ;
  input \sr[4]_i_155_3 ;
  input \sr[4]_i_155_4 ;
  input \sr[4]_i_155_5 ;
  input \sr[4]_i_155_6 ;
  input \sr[4]_i_155_7 ;
  input \sr[4]_i_164_2 ;
  input \sr[4]_i_164_3 ;
  input \sr[4]_i_159_3 ;
  input \sr[4]_i_159_4 ;
  input \sr[4]_i_159_5 ;
  input \sr[4]_i_155_8 ;
  input \sr[4]_i_155_9 ;
  input \sr[4]_i_155_10 ;
  input \sr[4]_i_155_11 ;
  input \rgf_c1bus_wb[4]_i_11_5 ;
  input \rgf_c1bus_wb[4]_i_11_6 ;
  input \sr[4]_i_159_6 ;
  input \sr[4]_i_159_7 ;
  input \sr[4]_i_15 ;
  input \sr[4]_i_15_0 ;
  input \sr[4]_i_15_1 ;
  input \sr[4]_i_57_0 ;
  input \sr[4]_i_57_1 ;
  input \sr[4]_i_57_2 ;
  input \sr[4]_i_66 ;
  input \sr[4]_i_66_0 ;
  input \sr[4]_i_57_3 ;
  input \sr[4]_i_67 ;
  input \sr[4]_i_67_0 ;
  input \sr[4]_i_139 ;
  input \sr[4]_i_139_0 ;
  input \rgf_c0bus_wb[12]_i_7 ;
  input \sr[4]_i_138_0 ;
  input \sr[4]_i_138_1 ;
  input \rgf_c0bus_wb[13]_i_13 ;
  input \sr[4]_i_129 ;
  input \sr[4]_i_197_0 ;
  input \sr[4]_i_197_1 ;
  input \sr[4]_i_197_2 ;
  input \sr[4]_i_185 ;
  input \sr[4]_i_185_0 ;
  input \rgf_c0bus_wb[4]_i_12 ;
  input \rgf_c0bus_wb[15]_i_23_0 ;
  input \rgf_c0bus_wb[15]_i_23_1 ;
  input \sr[4]_i_183_0 ;
  input \rgf_c0bus_wb[15]_i_23_2 ;
  input \sr[4]_i_183_1 ;
  input \sr[4]_i_186_0 ;
  input \sr[4]_i_186_1 ;
  input \sr[4]_i_183_2 ;
  input \rgf_c0bus_wb[15]_i_23_3 ;
  input \sr[4]_i_183_3 ;
  input \sr[4]_i_197_3 ;
  input \sr[4]_i_197_4 ;
  input \sr[4]_i_183_4 ;
  input [2:0]\sr[4]_i_197_5 ;
  input \rgf_c0bus_wb[15]_i_23_4 ;
  input \rgf_c0bus_wb[15]_i_23_5 ;
  input \sr[4]_i_183_5 ;
  input \rgf_c0bus_wb[15]_i_23_6 ;
  input \sr[4]_i_183_6 ;
  input \sr[4]_i_183_7 ;
  input \sr[4]_i_183_8 ;
  input \sr[4]_i_183_9 ;
  input \sr[4]_i_183_10 ;
  input \sr[4]_i_183_11 ;
  input \sr[4]_i_183_12 ;
  input \sr[4]_i_183_13 ;
  input \sr[4]_i_183_14 ;
  input \sr[4]_i_183_15 ;
  input \rgf_c0bus_wb[4]_i_8_0 ;
  input \rgf_c0bus_wb[4]_i_8_1 ;
  input \sr[4]_i_183_16 ;
  input \sr[4]_i_183_17 ;
  input \sr[4]_i_183_18 ;
  input \rgf_c0bus_wb[4]_i_8_2 ;
  input \rgf_c0bus_wb[4]_i_8_3 ;
  input \rgf_c0bus_wb[4]_i_8_4 ;
  input \sr[4]_i_197_6 ;
  input \sr[4]_i_197_7 ;
  input \rgf_c0bus_wb[4]_i_8_5 ;
  input \rgf_c0bus_wb[4]_i_8_6 ;
  input \rgf_c0bus_wb[4]_i_8_7 ;
  input \rgf_c0bus_wb[4]_i_8_8 ;
  input \rgf_c0bus_wb[4]_i_8_9 ;
  input \rgf_c0bus_wb[4]_i_12_0 ;
  input \rgf_c0bus_wb[4]_i_12_1 ;
  input \rgf_c0bus_wb[4]_i_12_2 ;
  input \rgf_c0bus_wb[15]_i_23_7 ;
  input \sr[4]_i_186_2 ;
  input \sr[4]_i_186_3 ;
  input \sr[4]_i_186_4 ;
  input \sr[4]_i_186_5 ;
  input \sr[4]_i_194_0 ;
  input \sr[4]_i_194_1 ;
  input \sr[4]_i_194_2 ;
  input \sr[4]_i_194_3 ;
  input \sr[4]_i_194_4 ;
  input \sr[4]_i_194_5 ;
  input \rgf_c0bus_wb[15]_i_23_8 ;
  input \rgf_c0bus_wb[15]_i_23_9 ;
  input \sr[4]_i_183_19 ;
  input [13:0]fdatx;
  input \ir0_id_fl[20]_i_4 ;
  input [13:0]fdat;
  input \nir_id_reg[20] ;
  input [3:0]a0bus_sel_0;
  input \i_/badr[15]_INST_0_i_135 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_135_0 ;
  input [0:0]ctl_sela0;
  input \i_/badr[15]_INST_0_i_135_1 ;
  input \bbus_o[4]_INST_0_i_7 ;
  input \bbus_o[4]_INST_0_i_7_0 ;
  input \bbus_o[3]_INST_0_i_7 ;
  input \bbus_o[3]_INST_0_i_7_0 ;
  input \bbus_o[2]_INST_0_i_7 ;
  input \bbus_o[2]_INST_0_i_7_0 ;
  input \bbus_o[1]_INST_0_i_7 ;
  input \bbus_o[1]_INST_0_i_7_0 ;
  input \bbus_o[0]_INST_0_i_7 ;
  input \bbus_o[0]_INST_0_i_7_0 ;
  input \i_/bdatw[15]_INST_0_i_34 ;
  input \i_/bbus_o[4]_INST_0_i_20 ;
  input \i_/bbus_o[4]_INST_0_i_21 ;
  input \i_/bbus_o[4]_INST_0_i_21_0 ;
  input [0:0]ctl_selb0_0;
  input \bbus_o[4]_INST_0_i_7_1 ;
  input \bbus_o[4]_INST_0_i_7_2 ;
  input \bbus_o[3]_INST_0_i_7_1 ;
  input \bbus_o[3]_INST_0_i_7_2 ;
  input \bbus_o[2]_INST_0_i_7_1 ;
  input \bbus_o[2]_INST_0_i_7_2 ;
  input \bbus_o[1]_INST_0_i_7_1 ;
  input \bbus_o[1]_INST_0_i_7_2 ;
  input \bbus_o[0]_INST_0_i_7_1 ;
  input \bbus_o[0]_INST_0_i_7_2 ;
  input \i_/bdatw[15]_INST_0_i_92 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_34_0 ;
  input [1:0]b0bus_sel_0;
  input \i_/bbus_o[4]_INST_0_i_20_0 ;
  input \i_/bbus_o[4]_INST_0_i_20_1 ;
  input \i_/bdatw[15]_INST_0_i_33 ;
  input \i_/bbus_o[4]_INST_0_i_21_1 ;
  input \i_/badr[0]_INST_0_i_18 ;
  input \i_/badr[0]_INST_0_i_18_0 ;
  input \i_/badr[0]_INST_0_i_18_1 ;
  input \rgf_c1bus_wb[4]_i_40 ;
  input \rgf_c1bus_wb[4]_i_40_0 ;
  input \rgf_c1bus_wb[4]_i_42 ;
  input \rgf_c1bus_wb[4]_i_42_0 ;
  input \rgf_c1bus_wb[4]_i_50 ;
  input \rgf_c1bus_wb[4]_i_50_0 ;
  input \rgf_c1bus_wb[4]_i_48 ;
  input \rgf_c1bus_wb[4]_i_48_0 ;
  input \rgf_c1bus_wb[4]_i_64 ;
  input \rgf_c1bus_wb[4]_i_64_0 ;
  input \rgf_c1bus_wb[4]_i_62 ;
  input \rgf_c1bus_wb[4]_i_62_0 ;
  input \rgf_c1bus_wb[4]_i_60 ;
  input \rgf_c1bus_wb[4]_i_60_0 ;
  input \rgf_c1bus_wb[4]_i_58 ;
  input \rgf_c1bus_wb[4]_i_58_0 ;
  input \rgf_c1bus_wb[4]_i_56 ;
  input \rgf_c1bus_wb[4]_i_56_0 ;
  input \rgf_c1bus_wb[4]_i_54 ;
  input \rgf_c1bus_wb[4]_i_54_0 ;
  input \rgf_c1bus_wb[4]_i_52 ;
  input \rgf_c1bus_wb[4]_i_52_0 ;
  input \rgf_c1bus_wb[4]_i_32 ;
  input \rgf_c1bus_wb[4]_i_32_0 ;
  input \rgf_c1bus_wb[4]_i_34 ;
  input \rgf_c1bus_wb[4]_i_34_0 ;
  input \rgf_c1bus_wb[4]_i_36 ;
  input \rgf_c1bus_wb[4]_i_36_0 ;
  input \rgf_c1bus_wb[4]_i_38 ;
  input \rgf_c1bus_wb[4]_i_38_0 ;
  input \sr[4]_i_239 ;
  input \sr[4]_i_239_0 ;
  input [2:0]a1bus_sel_0;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_212 ;
  input \i_/bdatw[15]_INST_0_i_124 ;
  input \i_/bdatw[15]_INST_0_i_121 ;
  input \i_/bdatw[15]_INST_0_i_121_0 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_121_1 ;
  input \i_/badr[15]_INST_0_i_52 ;
  input \bbus_o[4]_INST_0_i_7_3 ;
  input \bbus_o[4]_INST_0_i_7_4 ;
  input \bbus_o[3]_INST_0_i_7_3 ;
  input \bbus_o[3]_INST_0_i_7_4 ;
  input \bbus_o[2]_INST_0_i_7_3 ;
  input \bbus_o[2]_INST_0_i_7_4 ;
  input \bbus_o[1]_INST_0_i_7_3 ;
  input \bbus_o[1]_INST_0_i_7_4 ;
  input \bbus_o[0]_INST_0_i_7_3 ;
  input \bbus_o[0]_INST_0_i_7_4 ;
  input \bbus_o[4]_INST_0_i_7_5 ;
  input \bbus_o[4]_INST_0_i_7_6 ;
  input \bbus_o[3]_INST_0_i_7_5 ;
  input \bbus_o[3]_INST_0_i_7_6 ;
  input \bbus_o[2]_INST_0_i_7_5 ;
  input \bbus_o[2]_INST_0_i_7_6 ;
  input \bbus_o[1]_INST_0_i_7_5 ;
  input \bbus_o[1]_INST_0_i_7_6 ;
  input \bbus_o[0]_INST_0_i_7_5 ;
  input \bbus_o[0]_INST_0_i_7_6 ;
  input \rgf_c1bus_wb[4]_i_45 ;
  input \rgf_c1bus_wb[4]_i_45_0 ;
  input \rgf_c1bus_wb[4]_i_42_1 ;
  input \rgf_c1bus_wb[4]_i_42_2 ;
  input \rgf_c1bus_wb[4]_i_50_1 ;
  input \rgf_c1bus_wb[4]_i_50_2 ;
  input \rgf_c1bus_wb[4]_i_48_1 ;
  input \rgf_c1bus_wb[4]_i_48_2 ;
  input \rgf_c1bus_wb[4]_i_64_1 ;
  input \rgf_c1bus_wb[4]_i_64_2 ;
  input \rgf_c1bus_wb[4]_i_62_1 ;
  input \rgf_c1bus_wb[4]_i_62_2 ;
  input \rgf_c1bus_wb[4]_i_60_1 ;
  input \rgf_c1bus_wb[4]_i_60_2 ;
  input \rgf_c1bus_wb[4]_i_58_1 ;
  input \rgf_c1bus_wb[4]_i_58_2 ;
  input \rgf_c1bus_wb[4]_i_56_1 ;
  input \rgf_c1bus_wb[4]_i_56_2 ;
  input \rgf_c1bus_wb[4]_i_54_1 ;
  input \rgf_c1bus_wb[4]_i_54_2 ;
  input \rgf_c1bus_wb[4]_i_52_1 ;
  input \rgf_c1bus_wb[4]_i_52_2 ;
  input \rgf_c1bus_wb[4]_i_32_1 ;
  input \rgf_c1bus_wb[4]_i_32_2 ;
  input \rgf_c1bus_wb[4]_i_34_1 ;
  input \rgf_c1bus_wb[4]_i_34_2 ;
  input \rgf_c1bus_wb[4]_i_36_1 ;
  input \rgf_c1bus_wb[4]_i_36_2 ;
  input \rgf_c1bus_wb[4]_i_38_1 ;
  input \rgf_c1bus_wb[4]_i_38_2 ;
  input \rgf_c1bus_wb[4]_i_44 ;
  input \rgf_c1bus_wb[4]_i_44_0 ;
  input \bdatw[12]_INST_0_i_42 ;
  input \bdatw[12]_INST_0_i_42_0 ;
  input \bdatw[11]_INST_0_i_44 ;
  input \bdatw[11]_INST_0_i_44_0 ;
  input \bdatw[10]_INST_0_i_43 ;
  input \bdatw[10]_INST_0_i_43_0 ;
  input \bdatw[9]_INST_0_i_42 ;
  input \bdatw[9]_INST_0_i_42_0 ;
  input \bdatw[8]_INST_0_i_43 ;
  input \bdatw[8]_INST_0_i_43_0 ;
  input \badr[15]_INST_0_i_1_0 ;
  input \badr[15]_INST_0_i_1_1 ;
  input \badr[14]_INST_0_i_1 ;
  input \badr[14]_INST_0_i_1_0 ;
  input \badr[13]_INST_0_i_1 ;
  input \badr[13]_INST_0_i_1_0 ;
  input \badr[12]_INST_0_i_1 ;
  input \badr[12]_INST_0_i_1_0 ;
  input \badr[11]_INST_0_i_1 ;
  input \badr[11]_INST_0_i_1_0 ;
  input \badr[10]_INST_0_i_1 ;
  input \badr[10]_INST_0_i_1_0 ;
  input \badr[9]_INST_0_i_1 ;
  input \badr[9]_INST_0_i_1_0 ;
  input \badr[8]_INST_0_i_1 ;
  input \badr[8]_INST_0_i_1_0 ;
  input \badr[7]_INST_0_i_1 ;
  input \badr[7]_INST_0_i_1_0 ;
  input \badr[6]_INST_0_i_1 ;
  input \badr[6]_INST_0_i_1_0 ;
  input \badr[5]_INST_0_i_1 ;
  input \badr[5]_INST_0_i_1_0 ;
  input \badr[4]_INST_0_i_1 ;
  input \badr[4]_INST_0_i_1_0 ;
  input \badr[3]_INST_0_i_1 ;
  input \badr[3]_INST_0_i_1_0 ;
  input \badr[2]_INST_0_i_1 ;
  input \badr[2]_INST_0_i_1_0 ;
  input \badr[1]_INST_0_i_1 ;
  input \badr[1]_INST_0_i_1_0 ;
  input \badr[0]_INST_0_i_1 ;
  input \badr[0]_INST_0_i_1_0 ;
  input [0:0]\grn_reg[15]_19 ;
  input [15:0]\grn_reg[15]_20 ;
  input clk;
  input [0:0]\grn_reg[15]_21 ;
  input [15:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[15]_23 ;
  input [15:0]\grn_reg[15]_24 ;
  input [0:0]\grn_reg[15]_25 ;
  input [15:0]\grn_reg[15]_26 ;
  input [0:0]\grn_reg[15]_27 ;
  input [15:0]\grn_reg[15]_28 ;
  input [0:0]\grn_reg[15]_29 ;
  input [15:0]\grn_reg[15]_30 ;
  input [0:0]\grn_reg[15]_31 ;
  input [15:0]\grn_reg[15]_32 ;
  input [0:0]\grn_reg[15]_33 ;
  input [15:0]\grn_reg[15]_34 ;
  input [0:0]\grn_reg[15]_35 ;
  input [15:0]\grn_reg[15]_36 ;
  input [0:0]\grn_reg[15]_37 ;
  input [15:0]\grn_reg[15]_38 ;
  input [0:0]\grn_reg[15]_39 ;
  input [15:0]\grn_reg[15]_40 ;
  input [0:0]\grn_reg[15]_41 ;
  input [15:0]\grn_reg[15]_42 ;
  input [0:0]\grn_reg[15]_43 ;
  input [15:0]\grn_reg[15]_44 ;
  input [0:0]\grn_reg[15]_45 ;
  input [15:0]\grn_reg[15]_46 ;
  input [0:0]\grn_reg[15]_47 ;
  input [15:0]\grn_reg[15]_48 ;
  input [0:0]\grn_reg[15]_49 ;
  input [15:0]\grn_reg[15]_50 ;
     output [15:0]gr20;
     output [15:0]gr23;
     output [15:0]gr24;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr27;
     output [15:0]gr00;
     output [15:0]gr03;
     output [15:0]gr04;
     output [15:0]gr05;
     output [15:0]gr06;
     output [15:0]gr07;
  output fdat_12_sn_1;

  wire [0:0]SR;
  wire [3:0]a0bus_sel_0;
  wire [15:0]a1bus_b13;
  wire [2:0]a1bus_sel_0;
  wire a1buso2l_n_10;
  wire a1buso2l_n_12;
  wire a1buso2l_n_14;
  wire a1buso2l_n_16;
  wire a1buso2l_n_18;
  wire a1buso2l_n_2;
  wire a1buso2l_n_20;
  wire a1buso2l_n_22;
  wire a1buso2l_n_24;
  wire a1buso2l_n_26;
  wire a1buso2l_n_28;
  wire a1buso2l_n_30;
  wire a1buso2l_n_32;
  wire a1buso2l_n_4;
  wire a1buso2l_n_6;
  wire a1buso2l_n_8;
  wire a1buso_n_20;
  wire a1buso_n_22;
  wire a1buso_n_24;
  wire a1buso_n_26;
  wire a1buso_n_28;
  wire a1buso_n_30;
  wire a1buso_n_32;
  wire a1buso_n_34;
  wire a1buso_n_36;
  wire a1buso_n_38;
  wire a1buso_n_40;
  wire a1buso_n_42;
  wire a1buso_n_44;
  wire a1buso_n_46;
  wire [1:0]b0bus_sel_0;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[0]_INST_0_i_1_0 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1_0 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_1_0 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_1_0 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_1_0 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_1_1 ;
  wire \badr[15]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1_0 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1_0 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1_0 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[4]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1_0 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1_0 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1_0 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1_0 ;
  wire \badr[9]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1_0 ;
  wire \bbus_o[0]_INST_0_i_7 ;
  wire \bbus_o[0]_INST_0_i_7_0 ;
  wire \bbus_o[0]_INST_0_i_7_1 ;
  wire \bbus_o[0]_INST_0_i_7_2 ;
  wire \bbus_o[0]_INST_0_i_7_3 ;
  wire \bbus_o[0]_INST_0_i_7_4 ;
  wire \bbus_o[0]_INST_0_i_7_5 ;
  wire \bbus_o[0]_INST_0_i_7_6 ;
  wire \bbus_o[1]_INST_0_i_7 ;
  wire \bbus_o[1]_INST_0_i_7_0 ;
  wire \bbus_o[1]_INST_0_i_7_1 ;
  wire \bbus_o[1]_INST_0_i_7_2 ;
  wire \bbus_o[1]_INST_0_i_7_3 ;
  wire \bbus_o[1]_INST_0_i_7_4 ;
  wire \bbus_o[1]_INST_0_i_7_5 ;
  wire \bbus_o[1]_INST_0_i_7_6 ;
  wire \bbus_o[2]_INST_0_i_7 ;
  wire \bbus_o[2]_INST_0_i_7_0 ;
  wire \bbus_o[2]_INST_0_i_7_1 ;
  wire \bbus_o[2]_INST_0_i_7_2 ;
  wire \bbus_o[2]_INST_0_i_7_3 ;
  wire \bbus_o[2]_INST_0_i_7_4 ;
  wire \bbus_o[2]_INST_0_i_7_5 ;
  wire \bbus_o[2]_INST_0_i_7_6 ;
  wire \bbus_o[3]_INST_0_i_7 ;
  wire \bbus_o[3]_INST_0_i_7_0 ;
  wire \bbus_o[3]_INST_0_i_7_1 ;
  wire \bbus_o[3]_INST_0_i_7_2 ;
  wire \bbus_o[3]_INST_0_i_7_3 ;
  wire \bbus_o[3]_INST_0_i_7_4 ;
  wire \bbus_o[3]_INST_0_i_7_5 ;
  wire \bbus_o[3]_INST_0_i_7_6 ;
  wire \bbus_o[4]_INST_0_i_7 ;
  wire \bbus_o[4]_INST_0_i_7_0 ;
  wire \bbus_o[4]_INST_0_i_7_1 ;
  wire \bbus_o[4]_INST_0_i_7_2 ;
  wire \bbus_o[4]_INST_0_i_7_3 ;
  wire \bbus_o[4]_INST_0_i_7_4 ;
  wire \bbus_o[4]_INST_0_i_7_5 ;
  wire \bbus_o[4]_INST_0_i_7_6 ;
  wire \bdatw[10]_INST_0_i_43 ;
  wire \bdatw[10]_INST_0_i_43_0 ;
  wire \bdatw[11]_INST_0_i_44 ;
  wire \bdatw[11]_INST_0_i_44_0 ;
  wire \bdatw[12]_INST_0_i_42 ;
  wire \bdatw[12]_INST_0_i_42_0 ;
  wire \bdatw[8]_INST_0_i_43 ;
  wire \bdatw[8]_INST_0_i_43_0 ;
  wire \bdatw[9]_INST_0_i_42 ;
  wire \bdatw[9]_INST_0_i_42_0 ;
  wire clk;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [13:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_12_sn_1;
  wire [13:0]fdatx;
  wire \fdatx[15] ;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire gr6_bus1;
  wire gr6_bus1_0;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_10 ;
  wire \grn_reg[0]_11 ;
  wire \grn_reg[0]_12 ;
  wire \grn_reg[0]_13 ;
  wire \grn_reg[0]_14 ;
  wire \grn_reg[0]_15 ;
  wire \grn_reg[0]_16 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire \grn_reg[0]_9 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_10 ;
  wire \grn_reg[10]_11 ;
  wire \grn_reg[10]_12 ;
  wire \grn_reg[10]_13 ;
  wire \grn_reg[10]_14 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[10]_7 ;
  wire \grn_reg[10]_8 ;
  wire \grn_reg[10]_9 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_10 ;
  wire \grn_reg[11]_11 ;
  wire \grn_reg[11]_12 ;
  wire \grn_reg[11]_13 ;
  wire \grn_reg[11]_14 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[11]_7 ;
  wire \grn_reg[11]_8 ;
  wire \grn_reg[11]_9 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_10 ;
  wire \grn_reg[12]_11 ;
  wire \grn_reg[12]_12 ;
  wire \grn_reg[12]_13 ;
  wire \grn_reg[12]_14 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[12]_7 ;
  wire \grn_reg[12]_8 ;
  wire \grn_reg[12]_9 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_10 ;
  wire \grn_reg[13]_11 ;
  wire \grn_reg[13]_12 ;
  wire \grn_reg[13]_13 ;
  wire \grn_reg[13]_14 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[13]_7 ;
  wire \grn_reg[13]_8 ;
  wire \grn_reg[13]_9 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_10 ;
  wire \grn_reg[14]_11 ;
  wire \grn_reg[14]_12 ;
  wire \grn_reg[14]_13 ;
  wire \grn_reg[14]_14 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[14]_7 ;
  wire \grn_reg[14]_8 ;
  wire \grn_reg[14]_9 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire \grn_reg[15]_12 ;
  wire \grn_reg[15]_13 ;
  wire \grn_reg[15]_14 ;
  wire \grn_reg[15]_15 ;
  wire \grn_reg[15]_16 ;
  wire \grn_reg[15]_17 ;
  wire \grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [15:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [15:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [15:0]\grn_reg[15]_24 ;
  wire [0:0]\grn_reg[15]_25 ;
  wire [15:0]\grn_reg[15]_26 ;
  wire [0:0]\grn_reg[15]_27 ;
  wire [15:0]\grn_reg[15]_28 ;
  wire [0:0]\grn_reg[15]_29 ;
  wire [15:0]\grn_reg[15]_30 ;
  wire [0:0]\grn_reg[15]_31 ;
  wire [15:0]\grn_reg[15]_32 ;
  wire [0:0]\grn_reg[15]_33 ;
  wire [15:0]\grn_reg[15]_34 ;
  wire [0:0]\grn_reg[15]_35 ;
  wire [15:0]\grn_reg[15]_36 ;
  wire [0:0]\grn_reg[15]_37 ;
  wire [15:0]\grn_reg[15]_38 ;
  wire [0:0]\grn_reg[15]_39 ;
  wire \grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_40 ;
  wire [0:0]\grn_reg[15]_41 ;
  wire [15:0]\grn_reg[15]_42 ;
  wire [0:0]\grn_reg[15]_43 ;
  wire [15:0]\grn_reg[15]_44 ;
  wire [0:0]\grn_reg[15]_45 ;
  wire [15:0]\grn_reg[15]_46 ;
  wire [0:0]\grn_reg[15]_47 ;
  wire [15:0]\grn_reg[15]_48 ;
  wire [0:0]\grn_reg[15]_49 ;
  wire \grn_reg[15]_5 ;
  wire [15:0]\grn_reg[15]_50 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_10 ;
  wire \grn_reg[1]_11 ;
  wire \grn_reg[1]_12 ;
  wire \grn_reg[1]_13 ;
  wire \grn_reg[1]_14 ;
  wire \grn_reg[1]_15 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[1]_8 ;
  wire \grn_reg[1]_9 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_10 ;
  wire \grn_reg[2]_11 ;
  wire \grn_reg[2]_12 ;
  wire \grn_reg[2]_13 ;
  wire \grn_reg[2]_14 ;
  wire \grn_reg[2]_15 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[2]_8 ;
  wire \grn_reg[2]_9 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_10 ;
  wire \grn_reg[3]_11 ;
  wire \grn_reg[3]_12 ;
  wire \grn_reg[3]_13 ;
  wire \grn_reg[3]_14 ;
  wire \grn_reg[3]_15 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[3]_8 ;
  wire \grn_reg[3]_9 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_11 ;
  wire \grn_reg[4]_12 ;
  wire \grn_reg[4]_13 ;
  wire \grn_reg[4]_14 ;
  wire \grn_reg[4]_15 ;
  wire \grn_reg[4]_16 ;
  wire \grn_reg[4]_17 ;
  wire \grn_reg[4]_18 ;
  wire \grn_reg[4]_19 ;
  wire \grn_reg[4]_20 ;
  wire \grn_reg[4]_21 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_10 ;
  wire \grn_reg[5]_11 ;
  wire \grn_reg[5]_12 ;
  wire \grn_reg[5]_13 ;
  wire \grn_reg[5]_14 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[5]_7 ;
  wire \grn_reg[5]_8 ;
  wire \grn_reg[5]_9 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_10 ;
  wire \grn_reg[6]_11 ;
  wire \grn_reg[6]_12 ;
  wire \grn_reg[6]_13 ;
  wire \grn_reg[6]_14 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[6]_7 ;
  wire \grn_reg[6]_8 ;
  wire \grn_reg[6]_9 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_10 ;
  wire \grn_reg[7]_11 ;
  wire \grn_reg[7]_12 ;
  wire \grn_reg[7]_13 ;
  wire \grn_reg[7]_14 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[7]_7 ;
  wire \grn_reg[7]_8 ;
  wire \grn_reg[7]_9 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_10 ;
  wire \grn_reg[8]_11 ;
  wire \grn_reg[8]_12 ;
  wire \grn_reg[8]_13 ;
  wire \grn_reg[8]_14 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[8]_5 ;
  wire \grn_reg[8]_6 ;
  wire \grn_reg[8]_7 ;
  wire \grn_reg[8]_8 ;
  wire \grn_reg[8]_9 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_10 ;
  wire \grn_reg[9]_11 ;
  wire \grn_reg[9]_12 ;
  wire \grn_reg[9]_13 ;
  wire \grn_reg[9]_14 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire \grn_reg[9]_7 ;
  wire \grn_reg[9]_8 ;
  wire \grn_reg[9]_9 ;
  wire \i_/badr[0]_INST_0_i_18 ;
  wire \i_/badr[0]_INST_0_i_18_0 ;
  wire \i_/badr[0]_INST_0_i_18_1 ;
  wire \i_/badr[15]_INST_0_i_135 ;
  wire \i_/badr[15]_INST_0_i_135_0 ;
  wire \i_/badr[15]_INST_0_i_135_1 ;
  wire \i_/badr[15]_INST_0_i_52 ;
  wire \i_/bbus_o[4]_INST_0_i_20 ;
  wire \i_/bbus_o[4]_INST_0_i_20_0 ;
  wire \i_/bbus_o[4]_INST_0_i_20_1 ;
  wire \i_/bbus_o[4]_INST_0_i_21 ;
  wire \i_/bbus_o[4]_INST_0_i_21_0 ;
  wire \i_/bbus_o[4]_INST_0_i_21_1 ;
  wire \i_/bdatw[15]_INST_0_i_121 ;
  wire \i_/bdatw[15]_INST_0_i_121_0 ;
  wire \i_/bdatw[15]_INST_0_i_121_1 ;
  wire \i_/bdatw[15]_INST_0_i_124 ;
  wire \i_/bdatw[15]_INST_0_i_212 ;
  wire \i_/bdatw[15]_INST_0_i_33 ;
  wire \i_/bdatw[15]_INST_0_i_34 ;
  wire \i_/bdatw[15]_INST_0_i_34_0 ;
  wire \i_/bdatw[15]_INST_0_i_92 ;
  wire \ir0_id_fl[20]_i_4 ;
  wire \nir_id_reg[20] ;
  wire [15:0]p_0_in;
  wire \rgf_c0bus_wb[12]_i_7 ;
  wire \rgf_c0bus_wb[13]_i_13 ;
  wire \rgf_c0bus_wb[13]_i_27_0 ;
  wire \rgf_c0bus_wb[13]_i_30_0 ;
  wire \rgf_c0bus_wb[13]_i_30_n_0 ;
  wire \rgf_c0bus_wb[13]_i_31_n_0 ;
  wire \rgf_c0bus_wb[13]_i_32_n_0 ;
  wire \rgf_c0bus_wb[15]_i_23_0 ;
  wire \rgf_c0bus_wb[15]_i_23_1 ;
  wire \rgf_c0bus_wb[15]_i_23_2 ;
  wire \rgf_c0bus_wb[15]_i_23_3 ;
  wire \rgf_c0bus_wb[15]_i_23_4 ;
  wire \rgf_c0bus_wb[15]_i_23_5 ;
  wire \rgf_c0bus_wb[15]_i_23_6 ;
  wire \rgf_c0bus_wb[15]_i_23_7 ;
  wire \rgf_c0bus_wb[15]_i_23_8 ;
  wire \rgf_c0bus_wb[15]_i_23_9 ;
  wire \rgf_c0bus_wb[15]_i_27_n_0 ;
  wire \rgf_c0bus_wb[15]_i_28_n_0 ;
  wire \rgf_c0bus_wb[15]_i_29_n_0 ;
  wire \rgf_c0bus_wb[15]_i_30_n_0 ;
  wire \rgf_c0bus_wb[4]_i_12 ;
  wire \rgf_c0bus_wb[4]_i_12_0 ;
  wire \rgf_c0bus_wb[4]_i_12_1 ;
  wire \rgf_c0bus_wb[4]_i_12_2 ;
  wire \rgf_c0bus_wb[4]_i_22_n_0 ;
  wire \rgf_c0bus_wb[4]_i_23_n_0 ;
  wire \rgf_c0bus_wb[4]_i_24_n_0 ;
  wire \rgf_c0bus_wb[4]_i_25_n_0 ;
  wire \rgf_c0bus_wb[4]_i_26_0 ;
  wire \rgf_c0bus_wb[4]_i_26_n_0 ;
  wire \rgf_c0bus_wb[4]_i_29_0 ;
  wire \rgf_c0bus_wb[4]_i_29_n_0 ;
  wire \rgf_c0bus_wb[4]_i_30_n_0 ;
  wire \rgf_c0bus_wb[4]_i_31_0 ;
  wire \rgf_c0bus_wb[4]_i_31_n_0 ;
  wire \rgf_c0bus_wb[4]_i_32_0 ;
  wire \rgf_c0bus_wb[4]_i_32_n_0 ;
  wire \rgf_c0bus_wb[4]_i_33_0 ;
  wire \rgf_c0bus_wb[4]_i_8_0 ;
  wire \rgf_c0bus_wb[4]_i_8_1 ;
  wire \rgf_c0bus_wb[4]_i_8_2 ;
  wire \rgf_c0bus_wb[4]_i_8_3 ;
  wire \rgf_c0bus_wb[4]_i_8_4 ;
  wire \rgf_c0bus_wb[4]_i_8_5 ;
  wire \rgf_c0bus_wb[4]_i_8_6 ;
  wire \rgf_c0bus_wb[4]_i_8_7 ;
  wire \rgf_c0bus_wb[4]_i_8_8 ;
  wire \rgf_c0bus_wb[4]_i_8_9 ;
  wire \rgf_c1bus_wb[14]_i_28 ;
  wire [12:0]\rgf_c1bus_wb[4]_i_11 ;
  wire \rgf_c1bus_wb[4]_i_11_0 ;
  wire \rgf_c1bus_wb[4]_i_11_1 ;
  wire \rgf_c1bus_wb[4]_i_11_2 ;
  wire \rgf_c1bus_wb[4]_i_11_3 ;
  wire \rgf_c1bus_wb[4]_i_11_4 ;
  wire \rgf_c1bus_wb[4]_i_11_5 ;
  wire \rgf_c1bus_wb[4]_i_11_6 ;
  wire \rgf_c1bus_wb[4]_i_25_n_0 ;
  wire \rgf_c1bus_wb[4]_i_26_n_0 ;
  wire \rgf_c1bus_wb[4]_i_27_n_0 ;
  wire \rgf_c1bus_wb[4]_i_28_0 ;
  wire \rgf_c1bus_wb[4]_i_28_n_0 ;
  wire \rgf_c1bus_wb[4]_i_32 ;
  wire \rgf_c1bus_wb[4]_i_32_0 ;
  wire \rgf_c1bus_wb[4]_i_32_1 ;
  wire \rgf_c1bus_wb[4]_i_32_2 ;
  wire \rgf_c1bus_wb[4]_i_34 ;
  wire \rgf_c1bus_wb[4]_i_34_0 ;
  wire \rgf_c1bus_wb[4]_i_34_1 ;
  wire \rgf_c1bus_wb[4]_i_34_2 ;
  wire \rgf_c1bus_wb[4]_i_36 ;
  wire \rgf_c1bus_wb[4]_i_36_0 ;
  wire \rgf_c1bus_wb[4]_i_36_1 ;
  wire \rgf_c1bus_wb[4]_i_36_2 ;
  wire \rgf_c1bus_wb[4]_i_38 ;
  wire \rgf_c1bus_wb[4]_i_38_0 ;
  wire \rgf_c1bus_wb[4]_i_38_1 ;
  wire \rgf_c1bus_wb[4]_i_38_2 ;
  wire \rgf_c1bus_wb[4]_i_40 ;
  wire \rgf_c1bus_wb[4]_i_40_0 ;
  wire \rgf_c1bus_wb[4]_i_42 ;
  wire \rgf_c1bus_wb[4]_i_42_0 ;
  wire \rgf_c1bus_wb[4]_i_42_1 ;
  wire \rgf_c1bus_wb[4]_i_42_2 ;
  wire \rgf_c1bus_wb[4]_i_44 ;
  wire \rgf_c1bus_wb[4]_i_44_0 ;
  wire \rgf_c1bus_wb[4]_i_45 ;
  wire \rgf_c1bus_wb[4]_i_45_0 ;
  wire \rgf_c1bus_wb[4]_i_48 ;
  wire \rgf_c1bus_wb[4]_i_48_0 ;
  wire \rgf_c1bus_wb[4]_i_48_1 ;
  wire \rgf_c1bus_wb[4]_i_48_2 ;
  wire \rgf_c1bus_wb[4]_i_50 ;
  wire \rgf_c1bus_wb[4]_i_50_0 ;
  wire \rgf_c1bus_wb[4]_i_50_1 ;
  wire \rgf_c1bus_wb[4]_i_50_2 ;
  wire \rgf_c1bus_wb[4]_i_52 ;
  wire \rgf_c1bus_wb[4]_i_52_0 ;
  wire \rgf_c1bus_wb[4]_i_52_1 ;
  wire \rgf_c1bus_wb[4]_i_52_2 ;
  wire \rgf_c1bus_wb[4]_i_54 ;
  wire \rgf_c1bus_wb[4]_i_54_0 ;
  wire \rgf_c1bus_wb[4]_i_54_1 ;
  wire \rgf_c1bus_wb[4]_i_54_2 ;
  wire \rgf_c1bus_wb[4]_i_56 ;
  wire \rgf_c1bus_wb[4]_i_56_0 ;
  wire \rgf_c1bus_wb[4]_i_56_1 ;
  wire \rgf_c1bus_wb[4]_i_56_2 ;
  wire \rgf_c1bus_wb[4]_i_58 ;
  wire \rgf_c1bus_wb[4]_i_58_0 ;
  wire \rgf_c1bus_wb[4]_i_58_1 ;
  wire \rgf_c1bus_wb[4]_i_58_2 ;
  wire \rgf_c1bus_wb[4]_i_60 ;
  wire \rgf_c1bus_wb[4]_i_60_0 ;
  wire \rgf_c1bus_wb[4]_i_60_1 ;
  wire \rgf_c1bus_wb[4]_i_60_2 ;
  wire \rgf_c1bus_wb[4]_i_62 ;
  wire \rgf_c1bus_wb[4]_i_62_0 ;
  wire \rgf_c1bus_wb[4]_i_62_1 ;
  wire \rgf_c1bus_wb[4]_i_62_2 ;
  wire \rgf_c1bus_wb[4]_i_64 ;
  wire \rgf_c1bus_wb[4]_i_64_0 ;
  wire \rgf_c1bus_wb[4]_i_64_1 ;
  wire \rgf_c1bus_wb[4]_i_64_2 ;
  wire rst_n;
  wire \sp_reg[11] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[4] ;
  wire \sp_reg[6] ;
  wire \sr[4]_i_129 ;
  wire \sr[4]_i_130_n_0 ;
  wire \sr[4]_i_131_n_0 ;
  wire \sr[4]_i_133_0 ;
  wire \sr[4]_i_133_n_0 ;
  wire \sr[4]_i_138_0 ;
  wire \sr[4]_i_138_1 ;
  wire \sr[4]_i_139 ;
  wire \sr[4]_i_139_0 ;
  wire \sr[4]_i_15 ;
  wire \sr[4]_i_154_0 ;
  wire \sr[4]_i_154_1 ;
  wire \sr[4]_i_154_n_0 ;
  wire \sr[4]_i_155_0 ;
  wire \sr[4]_i_155_1 ;
  wire \sr[4]_i_155_10 ;
  wire \sr[4]_i_155_11 ;
  wire \sr[4]_i_155_2 ;
  wire \sr[4]_i_155_3 ;
  wire \sr[4]_i_155_4 ;
  wire \sr[4]_i_155_5 ;
  wire \sr[4]_i_155_6 ;
  wire \sr[4]_i_155_7 ;
  wire \sr[4]_i_155_8 ;
  wire \sr[4]_i_155_9 ;
  wire \sr[4]_i_155_n_0 ;
  wire \sr[4]_i_156_0 ;
  wire \sr[4]_i_156_n_0 ;
  wire \sr[4]_i_159_0 ;
  wire \sr[4]_i_159_1 ;
  wire \sr[4]_i_159_2 ;
  wire \sr[4]_i_159_3 ;
  wire \sr[4]_i_159_4 ;
  wire \sr[4]_i_159_5 ;
  wire \sr[4]_i_159_6 ;
  wire \sr[4]_i_159_7 ;
  wire \sr[4]_i_15_0 ;
  wire \sr[4]_i_15_1 ;
  wire \sr[4]_i_164_0 ;
  wire \sr[4]_i_164_1 ;
  wire \sr[4]_i_164_2 ;
  wire \sr[4]_i_164_3 ;
  wire \sr[4]_i_168 ;
  wire \sr[4]_i_168_0 ;
  wire \sr[4]_i_168_1 ;
  wire \sr[4]_i_168_2 ;
  wire \sr[4]_i_168_3 ;
  wire \sr[4]_i_170 ;
  wire \sr[4]_i_170_0 ;
  wire \sr[4]_i_170_1 ;
  wire \sr[4]_i_170_2 ;
  wire \sr[4]_i_170_3 ;
  wire \sr[4]_i_183_0 ;
  wire \sr[4]_i_183_1 ;
  wire \sr[4]_i_183_10 ;
  wire \sr[4]_i_183_11 ;
  wire \sr[4]_i_183_12 ;
  wire \sr[4]_i_183_13 ;
  wire \sr[4]_i_183_14 ;
  wire \sr[4]_i_183_15 ;
  wire \sr[4]_i_183_16 ;
  wire \sr[4]_i_183_17 ;
  wire \sr[4]_i_183_18 ;
  wire \sr[4]_i_183_19 ;
  wire \sr[4]_i_183_2 ;
  wire \sr[4]_i_183_3 ;
  wire \sr[4]_i_183_4 ;
  wire \sr[4]_i_183_5 ;
  wire \sr[4]_i_183_6 ;
  wire \sr[4]_i_183_7 ;
  wire \sr[4]_i_183_8 ;
  wire \sr[4]_i_183_9 ;
  wire \sr[4]_i_185 ;
  wire \sr[4]_i_185_0 ;
  wire \sr[4]_i_186_0 ;
  wire \sr[4]_i_186_1 ;
  wire \sr[4]_i_186_2 ;
  wire \sr[4]_i_186_3 ;
  wire \sr[4]_i_186_4 ;
  wire \sr[4]_i_186_5 ;
  wire \sr[4]_i_190_n_0 ;
  wire \sr[4]_i_191_n_0 ;
  wire \sr[4]_i_193_n_0 ;
  wire \sr[4]_i_194_0 ;
  wire \sr[4]_i_194_1 ;
  wire \sr[4]_i_194_2 ;
  wire \sr[4]_i_194_3 ;
  wire \sr[4]_i_194_4 ;
  wire \sr[4]_i_194_5 ;
  wire \sr[4]_i_194_n_0 ;
  wire \sr[4]_i_195_0 ;
  wire \sr[4]_i_195_n_0 ;
  wire \sr[4]_i_197_0 ;
  wire \sr[4]_i_197_1 ;
  wire \sr[4]_i_197_2 ;
  wire \sr[4]_i_197_3 ;
  wire \sr[4]_i_197_4 ;
  wire [2:0]\sr[4]_i_197_5 ;
  wire \sr[4]_i_197_6 ;
  wire \sr[4]_i_197_7 ;
  wire \sr[4]_i_198_n_0 ;
  wire \sr[4]_i_199_n_0 ;
  wire \sr[4]_i_200_0 ;
  wire \sr[4]_i_200_n_0 ;
  wire \sr[4]_i_208_n_0 ;
  wire \sr[4]_i_210_n_0 ;
  wire \sr[4]_i_211_n_0 ;
  wire \sr[4]_i_229_n_0 ;
  wire \sr[4]_i_230_n_0 ;
  wire \sr[4]_i_231_n_0 ;
  wire \sr[4]_i_232_0 ;
  wire \sr[4]_i_232_n_0 ;
  wire \sr[4]_i_239 ;
  wire \sr[4]_i_239_0 ;
  wire \sr[4]_i_27 ;
  wire \sr[4]_i_27_0 ;
  wire \sr[4]_i_27_1 ;
  wire \sr[4]_i_57_0 ;
  wire \sr[4]_i_57_1 ;
  wire \sr[4]_i_57_2 ;
  wire \sr[4]_i_57_3 ;
  wire \sr[4]_i_66 ;
  wire \sr[4]_i_66_0 ;
  wire \sr[4]_i_67 ;
  wire \sr[4]_i_67_0 ;
  wire \sr[4]_i_80_0 ;
  wire \sr[4]_i_80_1 ;
  wire \sr[4]_i_80_2 ;
  wire \sr[4]_i_83 ;
  wire \sr[4]_i_90 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[14] ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[3] ;

  mcss_rgf_bank_bus a0buso
       (.a0bus_sel_0(a0bus_sel_0),
        .\badr[15]_INST_0_i_12 (gr04),
        .\badr[15]_INST_0_i_12_0 (gr07),
        .\badr[15]_INST_0_i_12_1 (gr00),
        .ctl_sela0(ctl_sela0),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[10]_0 (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[11]_0 (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[12]_0 (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[13]_0 (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[14]_0 (\grn_reg[14]_0 ),
        .\grn_reg[15] (\grn_reg[15]_4 ),
        .\grn_reg[15]_0 (\grn_reg[15]_5 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\grn_reg[5] (\grn_reg[5] ),
        .\grn_reg[5]_0 (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[6]_0 (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[7]_0 (\grn_reg[7]_0 ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[8]_0 (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\grn_reg[9]_0 (\grn_reg[9]_0 ),
        .\i_/badr[15]_INST_0_i_135_0 (\i_/badr[15]_INST_0_i_135 ),
        .\i_/badr[15]_INST_0_i_135_1 (\i_/badr[15]_INST_0_i_135_0 ),
        .\i_/badr[15]_INST_0_i_135_2 (\i_/badr[15]_INST_0_i_135_1 ),
        .\i_/badr[15]_INST_0_i_54_0 (gr06),
        .\i_/badr[15]_INST_0_i_54_1 (gr05),
        .\i_/badr[15]_INST_0_i_55_0 (\sr[4]_i_197_5 [1:0]),
        .\i_/badr[15]_INST_0_i_55_1 (gr02),
        .\i_/badr[15]_INST_0_i_55_2 (gr01),
        .out(gr03));
  mcss_rgf_bank_bus_6 a0buso2l
       (.ctl_sela0(ctl_sela0),
        .ctl_sela0_rn(ctl_sela0_rn),
        .\grn_reg[0] (\grn_reg[0]_9 ),
        .\grn_reg[0]_0 (\grn_reg[0]_10 ),
        .\grn_reg[10] (\grn_reg[10]_7 ),
        .\grn_reg[10]_0 (\grn_reg[10]_8 ),
        .\grn_reg[11] (\grn_reg[11]_7 ),
        .\grn_reg[11]_0 (\grn_reg[11]_8 ),
        .\grn_reg[12] (\grn_reg[12]_7 ),
        .\grn_reg[12]_0 (\grn_reg[12]_8 ),
        .\grn_reg[13] (\grn_reg[13]_7 ),
        .\grn_reg[13]_0 (\grn_reg[13]_8 ),
        .\grn_reg[14] (\grn_reg[14]_7 ),
        .\grn_reg[14]_0 (\grn_reg[14]_8 ),
        .\grn_reg[15] (\grn_reg[15]_12 ),
        .\grn_reg[15]_0 (\grn_reg[15]_13 ),
        .\grn_reg[1] (\grn_reg[1]_8 ),
        .\grn_reg[1]_0 (\grn_reg[1]_9 ),
        .\grn_reg[2] (\grn_reg[2]_8 ),
        .\grn_reg[2]_0 (\grn_reg[2]_9 ),
        .\grn_reg[3] (\grn_reg[3]_8 ),
        .\grn_reg[3]_0 (\grn_reg[3]_9 ),
        .\grn_reg[4] (\grn_reg[4]_14 ),
        .\grn_reg[4]_0 (\grn_reg[4]_15 ),
        .\grn_reg[5] (\grn_reg[5]_7 ),
        .\grn_reg[5]_0 (\grn_reg[5]_8 ),
        .\grn_reg[6] (\grn_reg[6]_7 ),
        .\grn_reg[6]_0 (\grn_reg[6]_8 ),
        .\grn_reg[7] (\grn_reg[7]_7 ),
        .\grn_reg[7]_0 (\grn_reg[7]_8 ),
        .\grn_reg[8] (\grn_reg[8]_7 ),
        .\grn_reg[8]_0 (\grn_reg[8]_8 ),
        .\grn_reg[9] (\grn_reg[9]_7 ),
        .\grn_reg[9]_0 (\grn_reg[9]_8 ),
        .\i_/badr[15]_INST_0_i_52_0 (\i_/badr[15]_INST_0_i_52 ),
        .\i_/badr[15]_INST_0_i_52_1 (\i_/badr[15]_INST_0_i_135_0 ),
        .\i_/badr[15]_INST_0_i_52_2 (\i_/badr[15]_INST_0_i_135_1 ),
        .\i_/rgf_c0bus_wb[4]_i_108_0 (gr20),
        .\i_/rgf_c0bus_wb[4]_i_108_1 (gr26),
        .\i_/rgf_c0bus_wb[4]_i_108_2 (gr25),
        .\i_/rgf_c0bus_wb[4]_i_108_3 (gr23),
        .\i_/rgf_c0bus_wb[4]_i_108_4 (gr24),
        .\i_/rgf_c0bus_wb[4]_i_108_5 (gr22),
        .\i_/rgf_c0bus_wb[4]_i_108_6 (gr21),
        .out(gr27),
        .p_0_in(p_0_in));
  mcss_rgf_bank_bus_7 a1buso
       (.a1bus_sel_0(a1bus_sel_0),
        .\badr[15]_INST_0_i_31 (\sr[4]_i_197_5 [1:0]),
        .\grn_reg[0] (\grn_reg[0]_3 ),
        .\grn_reg[0]_0 (\grn_reg[0]_4 ),
        .\grn_reg[0]_1 (\grn_reg[0]_5 ),
        .\grn_reg[10] (\grn_reg[10]_3 ),
        .\grn_reg[10]_0 (\grn_reg[10]_4 ),
        .\grn_reg[10]_1 (a1buso_n_28),
        .\grn_reg[11] (\grn_reg[11]_3 ),
        .\grn_reg[11]_0 (\grn_reg[11]_4 ),
        .\grn_reg[11]_1 (a1buso_n_26),
        .\grn_reg[12] (\grn_reg[12]_3 ),
        .\grn_reg[12]_0 (\grn_reg[12]_4 ),
        .\grn_reg[12]_1 (a1buso_n_24),
        .\grn_reg[13] (\grn_reg[13]_3 ),
        .\grn_reg[13]_0 (\grn_reg[13]_4 ),
        .\grn_reg[13]_1 (a1buso_n_22),
        .\grn_reg[14] (\grn_reg[14]_3 ),
        .\grn_reg[14]_0 (\grn_reg[14]_4 ),
        .\grn_reg[14]_1 (a1buso_n_20),
        .\grn_reg[15] (\grn_reg[15]_8 ),
        .\grn_reg[15]_0 (\grn_reg[15]_9 ),
        .\grn_reg[15]_1 (\grn_reg[15]_10 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[1]_0 (\grn_reg[1]_4 ),
        .\grn_reg[1]_1 (a1buso_n_46),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[2]_0 (\grn_reg[2]_4 ),
        .\grn_reg[2]_1 (a1buso_n_44),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[3]_1 (a1buso_n_42),
        .\grn_reg[4] (\grn_reg[4]_9 ),
        .\grn_reg[4]_0 (\grn_reg[4]_10 ),
        .\grn_reg[4]_1 (a1buso_n_40),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\grn_reg[5]_1 (a1buso_n_38),
        .\grn_reg[6] (\grn_reg[6]_3 ),
        .\grn_reg[6]_0 (\grn_reg[6]_4 ),
        .\grn_reg[6]_1 (a1buso_n_36),
        .\grn_reg[7] (\grn_reg[7]_3 ),
        .\grn_reg[7]_0 (\grn_reg[7]_4 ),
        .\grn_reg[7]_1 (a1buso_n_34),
        .\grn_reg[8] (\grn_reg[8]_3 ),
        .\grn_reg[8]_0 (\grn_reg[8]_4 ),
        .\grn_reg[8]_1 (a1buso_n_32),
        .\grn_reg[9] (\grn_reg[9]_3 ),
        .\grn_reg[9]_0 (\grn_reg[9]_4 ),
        .\grn_reg[9]_1 (a1buso_n_30),
        .\i_/badr[0]_INST_0_i_18_0 (\i_/badr[0]_INST_0_i_18 ),
        .\i_/badr[0]_INST_0_i_18_1 (\i_/badr[0]_INST_0_i_18_0 ),
        .\i_/badr[0]_INST_0_i_18_2 (\i_/badr[0]_INST_0_i_18_1 ),
        .\i_/badr[0]_INST_0_i_18_3 (\i_/badr[15]_INST_0_i_135 ),
        .\i_/badr[15]_INST_0_i_29_0 (gr02),
        .\i_/badr[15]_INST_0_i_29_1 (gr01),
        .out(gr03),
        .\rgf_c1bus_wb[4]_i_32 (\rgf_c1bus_wb[4]_i_32 ),
        .\rgf_c1bus_wb[4]_i_32_0 (\rgf_c1bus_wb[4]_i_32_0 ),
        .\rgf_c1bus_wb[4]_i_34 (\rgf_c1bus_wb[4]_i_34 ),
        .\rgf_c1bus_wb[4]_i_34_0 (\rgf_c1bus_wb[4]_i_34_0 ),
        .\rgf_c1bus_wb[4]_i_36 (\rgf_c1bus_wb[4]_i_36 ),
        .\rgf_c1bus_wb[4]_i_36_0 (\rgf_c1bus_wb[4]_i_36_0 ),
        .\rgf_c1bus_wb[4]_i_38 (\rgf_c1bus_wb[4]_i_38 ),
        .\rgf_c1bus_wb[4]_i_38_0 (\rgf_c1bus_wb[4]_i_38_0 ),
        .\rgf_c1bus_wb[4]_i_40 (\rgf_c1bus_wb[4]_i_40 ),
        .\rgf_c1bus_wb[4]_i_40_0 (\rgf_c1bus_wb[4]_i_40_0 ),
        .\rgf_c1bus_wb[4]_i_40_1 (gr06),
        .\rgf_c1bus_wb[4]_i_42 (\rgf_c1bus_wb[4]_i_42 ),
        .\rgf_c1bus_wb[4]_i_42_0 (\rgf_c1bus_wb[4]_i_42_0 ),
        .\rgf_c1bus_wb[4]_i_45 (gr04),
        .\rgf_c1bus_wb[4]_i_45_0 (gr07),
        .\rgf_c1bus_wb[4]_i_45_1 (gr00),
        .\rgf_c1bus_wb[4]_i_48 (\rgf_c1bus_wb[4]_i_48 ),
        .\rgf_c1bus_wb[4]_i_48_0 (\rgf_c1bus_wb[4]_i_48_0 ),
        .\rgf_c1bus_wb[4]_i_50 (\rgf_c1bus_wb[4]_i_50 ),
        .\rgf_c1bus_wb[4]_i_50_0 (\rgf_c1bus_wb[4]_i_50_0 ),
        .\rgf_c1bus_wb[4]_i_52 (\rgf_c1bus_wb[4]_i_52 ),
        .\rgf_c1bus_wb[4]_i_52_0 (\rgf_c1bus_wb[4]_i_52_0 ),
        .\rgf_c1bus_wb[4]_i_54 (\rgf_c1bus_wb[4]_i_54 ),
        .\rgf_c1bus_wb[4]_i_54_0 (\rgf_c1bus_wb[4]_i_54_0 ),
        .\rgf_c1bus_wb[4]_i_56 (\rgf_c1bus_wb[4]_i_56 ),
        .\rgf_c1bus_wb[4]_i_56_0 (\rgf_c1bus_wb[4]_i_56_0 ),
        .\rgf_c1bus_wb[4]_i_58 (\rgf_c1bus_wb[4]_i_58 ),
        .\rgf_c1bus_wb[4]_i_58_0 (\rgf_c1bus_wb[4]_i_58_0 ),
        .\rgf_c1bus_wb[4]_i_60 (\rgf_c1bus_wb[4]_i_60 ),
        .\rgf_c1bus_wb[4]_i_60_0 (\rgf_c1bus_wb[4]_i_60_0 ),
        .\rgf_c1bus_wb[4]_i_62 (\rgf_c1bus_wb[4]_i_62 ),
        .\rgf_c1bus_wb[4]_i_62_0 (\rgf_c1bus_wb[4]_i_62_0 ),
        .\rgf_c1bus_wb[4]_i_64 (\rgf_c1bus_wb[4]_i_64 ),
        .\rgf_c1bus_wb[4]_i_64_0 (\rgf_c1bus_wb[4]_i_64_0 ),
        .\sr[4]_i_239 (\sr[4]_i_239 ),
        .\sr[4]_i_239_0 (\sr[4]_i_239_0 ),
        .\sr_reg[1] (gr6_bus1));
  mcss_rgf_bank_bus_8 a1buso2l
       (.a1bus_sel_0(a1bus_sel_0),
        .\badr[15]_INST_0_i_7 (gr20),
        .\grn_reg[0] (\grn_reg[0]_13 ),
        .\grn_reg[0]_0 (a1buso2l_n_32),
        .\grn_reg[0]_1 (\grn_reg[0]_14 ),
        .\grn_reg[10] (\grn_reg[10]_11 ),
        .\grn_reg[10]_0 (a1buso2l_n_12),
        .\grn_reg[10]_1 (\grn_reg[10]_12 ),
        .\grn_reg[11] (\grn_reg[11]_11 ),
        .\grn_reg[11]_0 (a1buso2l_n_10),
        .\grn_reg[11]_1 (\grn_reg[11]_12 ),
        .\grn_reg[12] (\grn_reg[12]_11 ),
        .\grn_reg[12]_0 (a1buso2l_n_8),
        .\grn_reg[12]_1 (\grn_reg[12]_12 ),
        .\grn_reg[13] (\grn_reg[13]_11 ),
        .\grn_reg[13]_0 (a1buso2l_n_6),
        .\grn_reg[13]_1 (\grn_reg[13]_12 ),
        .\grn_reg[14] (\grn_reg[14]_11 ),
        .\grn_reg[14]_0 (a1buso2l_n_4),
        .\grn_reg[14]_1 (\grn_reg[14]_12 ),
        .\grn_reg[15] (\grn_reg[15]_16 ),
        .\grn_reg[15]_0 (a1buso2l_n_2),
        .\grn_reg[15]_1 (\grn_reg[15]_17 ),
        .\grn_reg[1] (\grn_reg[1]_12 ),
        .\grn_reg[1]_0 (a1buso2l_n_30),
        .\grn_reg[1]_1 (\grn_reg[1]_13 ),
        .\grn_reg[2] (\grn_reg[2]_12 ),
        .\grn_reg[2]_0 (a1buso2l_n_28),
        .\grn_reg[2]_1 (\grn_reg[2]_13 ),
        .\grn_reg[3] (\grn_reg[3]_12 ),
        .\grn_reg[3]_0 (a1buso2l_n_26),
        .\grn_reg[3]_1 (\grn_reg[3]_13 ),
        .\grn_reg[4] (\grn_reg[4]_18 ),
        .\grn_reg[4]_0 (a1buso2l_n_24),
        .\grn_reg[4]_1 (\grn_reg[4]_19 ),
        .\grn_reg[5] (\grn_reg[5]_11 ),
        .\grn_reg[5]_0 (a1buso2l_n_22),
        .\grn_reg[5]_1 (\grn_reg[5]_12 ),
        .\grn_reg[6] (\grn_reg[6]_11 ),
        .\grn_reg[6]_0 (a1buso2l_n_20),
        .\grn_reg[6]_1 (\grn_reg[6]_12 ),
        .\grn_reg[7] (\grn_reg[7]_11 ),
        .\grn_reg[7]_0 (a1buso2l_n_18),
        .\grn_reg[7]_1 (\grn_reg[7]_12 ),
        .\grn_reg[8] (\grn_reg[8]_11 ),
        .\grn_reg[8]_0 (a1buso2l_n_16),
        .\grn_reg[8]_1 (\grn_reg[8]_12 ),
        .\grn_reg[9] (\grn_reg[9]_11 ),
        .\grn_reg[9]_0 (a1buso2l_n_14),
        .\grn_reg[9]_1 (\grn_reg[9]_12 ),
        .\i_/badr[0]_INST_0_i_21_0 (\i_/badr[15]_INST_0_i_52 ),
        .\i_/badr[15]_INST_0_i_32_0 (\i_/badr[0]_INST_0_i_18 ),
        .\i_/badr[15]_INST_0_i_32_1 (\i_/badr[0]_INST_0_i_18_0 ),
        .\i_/badr[15]_INST_0_i_32_2 (\i_/badr[0]_INST_0_i_18_1 ),
        .\i_/badr[15]_INST_0_i_32_3 (gr22),
        .\i_/badr[15]_INST_0_i_32_4 (gr21),
        .\i_/rgf_c1bus_wb[4]_i_87_0 (\sr[4]_i_197_5 [1:0]),
        .out(gr27),
        .\rgf_c1bus_wb[4]_i_32 (\rgf_c1bus_wb[4]_i_32_1 ),
        .\rgf_c1bus_wb[4]_i_32_0 (\rgf_c1bus_wb[4]_i_32_2 ),
        .\rgf_c1bus_wb[4]_i_34 (\rgf_c1bus_wb[4]_i_34_1 ),
        .\rgf_c1bus_wb[4]_i_34_0 (\rgf_c1bus_wb[4]_i_34_2 ),
        .\rgf_c1bus_wb[4]_i_36 (\rgf_c1bus_wb[4]_i_36_1 ),
        .\rgf_c1bus_wb[4]_i_36_0 (\rgf_c1bus_wb[4]_i_36_2 ),
        .\rgf_c1bus_wb[4]_i_38 (\rgf_c1bus_wb[4]_i_38_1 ),
        .\rgf_c1bus_wb[4]_i_38_0 (\rgf_c1bus_wb[4]_i_38_2 ),
        .\rgf_c1bus_wb[4]_i_42 (\rgf_c1bus_wb[4]_i_42_1 ),
        .\rgf_c1bus_wb[4]_i_42_0 (\rgf_c1bus_wb[4]_i_42_2 ),
        .\rgf_c1bus_wb[4]_i_44 (\rgf_c1bus_wb[4]_i_44 ),
        .\rgf_c1bus_wb[4]_i_44_0 (\rgf_c1bus_wb[4]_i_44_0 ),
        .\rgf_c1bus_wb[4]_i_45 (\rgf_c1bus_wb[4]_i_45 ),
        .\rgf_c1bus_wb[4]_i_45_0 (\rgf_c1bus_wb[4]_i_45_0 ),
        .\rgf_c1bus_wb[4]_i_45_1 (gr26),
        .\rgf_c1bus_wb[4]_i_45_2 (gr23),
        .\rgf_c1bus_wb[4]_i_45_3 (gr24),
        .\rgf_c1bus_wb[4]_i_48 (\rgf_c1bus_wb[4]_i_48_1 ),
        .\rgf_c1bus_wb[4]_i_48_0 (\rgf_c1bus_wb[4]_i_48_2 ),
        .\rgf_c1bus_wb[4]_i_50 (\rgf_c1bus_wb[4]_i_50_1 ),
        .\rgf_c1bus_wb[4]_i_50_0 (\rgf_c1bus_wb[4]_i_50_2 ),
        .\rgf_c1bus_wb[4]_i_52 (\rgf_c1bus_wb[4]_i_52_1 ),
        .\rgf_c1bus_wb[4]_i_52_0 (\rgf_c1bus_wb[4]_i_52_2 ),
        .\rgf_c1bus_wb[4]_i_54 (\rgf_c1bus_wb[4]_i_54_1 ),
        .\rgf_c1bus_wb[4]_i_54_0 (\rgf_c1bus_wb[4]_i_54_2 ),
        .\rgf_c1bus_wb[4]_i_56 (\rgf_c1bus_wb[4]_i_56_1 ),
        .\rgf_c1bus_wb[4]_i_56_0 (\rgf_c1bus_wb[4]_i_56_2 ),
        .\rgf_c1bus_wb[4]_i_58 (\rgf_c1bus_wb[4]_i_58_1 ),
        .\rgf_c1bus_wb[4]_i_58_0 (\rgf_c1bus_wb[4]_i_58_2 ),
        .\rgf_c1bus_wb[4]_i_60 (\rgf_c1bus_wb[4]_i_60_1 ),
        .\rgf_c1bus_wb[4]_i_60_0 (\rgf_c1bus_wb[4]_i_60_2 ),
        .\rgf_c1bus_wb[4]_i_62 (\rgf_c1bus_wb[4]_i_62_1 ),
        .\rgf_c1bus_wb[4]_i_62_0 (\rgf_c1bus_wb[4]_i_62_2 ),
        .\rgf_c1bus_wb[4]_i_64 (\rgf_c1bus_wb[4]_i_64_1 ),
        .\rgf_c1bus_wb[4]_i_64_0 (\rgf_c1bus_wb[4]_i_64_2 ),
        .\sr_reg[1] (gr6_bus1_0));
  mcss_rgf_bank_bus_9 b0buso
       (.b0bus_sel_0(b0bus_sel_0),
        .\bbus_o[0]_INST_0_i_7 (\bbus_o[0]_INST_0_i_7 ),
        .\bbus_o[0]_INST_0_i_7_0 (\bbus_o[0]_INST_0_i_7_0 ),
        .\bbus_o[0]_INST_0_i_7_1 (\bbus_o[0]_INST_0_i_7_1 ),
        .\bbus_o[0]_INST_0_i_7_2 (\bbus_o[0]_INST_0_i_7_2 ),
        .\bbus_o[1]_INST_0_i_7 (\bbus_o[1]_INST_0_i_7 ),
        .\bbus_o[1]_INST_0_i_7_0 (\bbus_o[1]_INST_0_i_7_0 ),
        .\bbus_o[1]_INST_0_i_7_1 (\bbus_o[1]_INST_0_i_7_1 ),
        .\bbus_o[1]_INST_0_i_7_2 (\bbus_o[1]_INST_0_i_7_2 ),
        .\bbus_o[2]_INST_0_i_7 (\bbus_o[2]_INST_0_i_7 ),
        .\bbus_o[2]_INST_0_i_7_0 (\bbus_o[2]_INST_0_i_7_0 ),
        .\bbus_o[2]_INST_0_i_7_1 (\bbus_o[2]_INST_0_i_7_1 ),
        .\bbus_o[2]_INST_0_i_7_2 (\bbus_o[2]_INST_0_i_7_2 ),
        .\bbus_o[3]_INST_0_i_7 (\bbus_o[3]_INST_0_i_7 ),
        .\bbus_o[3]_INST_0_i_7_0 (\bbus_o[3]_INST_0_i_7_0 ),
        .\bbus_o[3]_INST_0_i_7_1 (\bbus_o[3]_INST_0_i_7_1 ),
        .\bbus_o[3]_INST_0_i_7_2 (\bbus_o[3]_INST_0_i_7_2 ),
        .\bbus_o[4]_INST_0_i_7 (\bbus_o[4]_INST_0_i_7 ),
        .\bbus_o[4]_INST_0_i_7_0 (\bbus_o[4]_INST_0_i_7_0 ),
        .\bbus_o[4]_INST_0_i_7_1 (\bbus_o[4]_INST_0_i_7_1 ),
        .\bbus_o[4]_INST_0_i_7_2 (\bbus_o[4]_INST_0_i_7_2 ),
        .\bdatw[15]_INST_0_i_11 (gr04[15:5]),
        .\bdatw[15]_INST_0_i_11_0 (gr07[15:5]),
        .\bdatw[15]_INST_0_i_11_1 (gr00),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[0] (\grn_reg[0]_1 ),
        .\grn_reg[0]_0 (\grn_reg[0]_2 ),
        .\grn_reg[10] (\grn_reg[10]_1 ),
        .\grn_reg[10]_0 (\grn_reg[10]_2 ),
        .\grn_reg[11] (\grn_reg[11]_1 ),
        .\grn_reg[11]_0 (\grn_reg[11]_2 ),
        .\grn_reg[12] (\grn_reg[12]_1 ),
        .\grn_reg[12]_0 (\grn_reg[12]_2 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[13]_0 (\grn_reg[13]_2 ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[14]_0 (\grn_reg[14]_2 ),
        .\grn_reg[15] (\grn_reg[15]_6 ),
        .\grn_reg[15]_0 (\grn_reg[15]_7 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (\grn_reg[1]_2 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (\grn_reg[2]_2 ),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (\grn_reg[3]_2 ),
        .\grn_reg[4] (\grn_reg[4]_7 ),
        .\grn_reg[4]_0 (\grn_reg[4]_8 ),
        .\grn_reg[5] (\grn_reg[5]_1 ),
        .\grn_reg[5]_0 (\grn_reg[5]_2 ),
        .\grn_reg[6] (\grn_reg[6]_1 ),
        .\grn_reg[6]_0 (\grn_reg[6]_2 ),
        .\grn_reg[7] (\grn_reg[7]_1 ),
        .\grn_reg[7]_0 (\grn_reg[7]_2 ),
        .\grn_reg[8] (\grn_reg[8]_1 ),
        .\grn_reg[8]_0 (\grn_reg[8]_2 ),
        .\grn_reg[9] (\grn_reg[9]_1 ),
        .\grn_reg[9]_0 (\grn_reg[9]_2 ),
        .\i_/bbus_o[4]_INST_0_i_20_0 (\i_/bbus_o[4]_INST_0_i_20 ),
        .\i_/bbus_o[4]_INST_0_i_20_1 (\i_/bbus_o[4]_INST_0_i_20_0 ),
        .\i_/bbus_o[4]_INST_0_i_20_2 (\i_/bbus_o[4]_INST_0_i_20_1 ),
        .\i_/bbus_o[4]_INST_0_i_21_0 (\i_/badr[15]_INST_0_i_135 ),
        .\i_/bbus_o[4]_INST_0_i_21_1 (\i_/bbus_o[4]_INST_0_i_21 ),
        .\i_/bbus_o[4]_INST_0_i_21_2 (\i_/bbus_o[4]_INST_0_i_21_0 ),
        .\i_/bbus_o[4]_INST_0_i_21_3 (\i_/bbus_o[4]_INST_0_i_21_1 ),
        .\i_/bbus_o[5]_INST_0_i_14_0 (\sr[4]_i_197_5 [1:0]),
        .\i_/bdatw[15]_INST_0_i_33_0 (gr01),
        .\i_/bdatw[15]_INST_0_i_33_1 (gr02),
        .\i_/bdatw[15]_INST_0_i_33_2 (\i_/bdatw[15]_INST_0_i_33 ),
        .\i_/bdatw[15]_INST_0_i_34_0 (\i_/bdatw[15]_INST_0_i_34 ),
        .\i_/bdatw[15]_INST_0_i_34_1 (gr06),
        .\i_/bdatw[15]_INST_0_i_34_2 (gr05[15:5]),
        .\i_/bdatw[15]_INST_0_i_34_3 (\i_/bdatw[15]_INST_0_i_34_0 ),
        .\i_/bdatw[15]_INST_0_i_92_0 (\i_/bdatw[15]_INST_0_i_92 ),
        .out(gr03[15:5]));
  mcss_rgf_bank_bus_10 b0buso2l
       (.b0bus_sel_0(b0bus_sel_0),
        .\bbus_o[0]_INST_0_i_7 (\bbus_o[0]_INST_0_i_7_3 ),
        .\bbus_o[0]_INST_0_i_7_0 (\bbus_o[0]_INST_0_i_7_4 ),
        .\bbus_o[0]_INST_0_i_7_1 (\bbus_o[0]_INST_0_i_7_5 ),
        .\bbus_o[0]_INST_0_i_7_2 (\bbus_o[0]_INST_0_i_7_6 ),
        .\bbus_o[1]_INST_0_i_7 (\bbus_o[1]_INST_0_i_7_3 ),
        .\bbus_o[1]_INST_0_i_7_0 (\bbus_o[1]_INST_0_i_7_4 ),
        .\bbus_o[1]_INST_0_i_7_1 (\bbus_o[1]_INST_0_i_7_5 ),
        .\bbus_o[1]_INST_0_i_7_2 (\bbus_o[1]_INST_0_i_7_6 ),
        .\bbus_o[2]_INST_0_i_7 (\bbus_o[2]_INST_0_i_7_3 ),
        .\bbus_o[2]_INST_0_i_7_0 (\bbus_o[2]_INST_0_i_7_4 ),
        .\bbus_o[2]_INST_0_i_7_1 (\bbus_o[2]_INST_0_i_7_5 ),
        .\bbus_o[2]_INST_0_i_7_2 (\bbus_o[2]_INST_0_i_7_6 ),
        .\bbus_o[3]_INST_0_i_7 (\bbus_o[3]_INST_0_i_7_3 ),
        .\bbus_o[3]_INST_0_i_7_0 (\bbus_o[3]_INST_0_i_7_4 ),
        .\bbus_o[3]_INST_0_i_7_1 (\bbus_o[3]_INST_0_i_7_5 ),
        .\bbus_o[3]_INST_0_i_7_2 (\bbus_o[3]_INST_0_i_7_6 ),
        .\bbus_o[4]_INST_0_i_7 (\bbus_o[4]_INST_0_i_7_3 ),
        .\bbus_o[4]_INST_0_i_7_0 (\bbus_o[4]_INST_0_i_7_4 ),
        .\bbus_o[4]_INST_0_i_7_1 (\bbus_o[4]_INST_0_i_7_5 ),
        .\bbus_o[4]_INST_0_i_7_2 (\bbus_o[4]_INST_0_i_7_6 ),
        .\bdatw[15]_INST_0_i_11 (gr20),
        .\bdatw[15]_INST_0_i_11_0 (gr23[15:5]),
        .\bdatw[15]_INST_0_i_11_1 (gr24[15:5]),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .\grn_reg[0] (\grn_reg[0]_11 ),
        .\grn_reg[0]_0 (\grn_reg[0]_12 ),
        .\grn_reg[10] (\grn_reg[10]_9 ),
        .\grn_reg[10]_0 (\grn_reg[10]_10 ),
        .\grn_reg[11] (\grn_reg[11]_9 ),
        .\grn_reg[11]_0 (\grn_reg[11]_10 ),
        .\grn_reg[12] (\grn_reg[12]_9 ),
        .\grn_reg[12]_0 (\grn_reg[12]_10 ),
        .\grn_reg[13] (\grn_reg[13]_9 ),
        .\grn_reg[13]_0 (\grn_reg[13]_10 ),
        .\grn_reg[14] (\grn_reg[14]_9 ),
        .\grn_reg[14]_0 (\grn_reg[14]_10 ),
        .\grn_reg[15] (\grn_reg[15]_14 ),
        .\grn_reg[15]_0 (\grn_reg[15]_15 ),
        .\grn_reg[1] (\grn_reg[1]_10 ),
        .\grn_reg[1]_0 (\grn_reg[1]_11 ),
        .\grn_reg[2] (\grn_reg[2]_10 ),
        .\grn_reg[2]_0 (\grn_reg[2]_11 ),
        .\grn_reg[3] (\grn_reg[3]_10 ),
        .\grn_reg[3]_0 (\grn_reg[3]_11 ),
        .\grn_reg[4] (\grn_reg[4]_16 ),
        .\grn_reg[4]_0 (\grn_reg[4]_17 ),
        .\grn_reg[5] (\grn_reg[5]_9 ),
        .\grn_reg[5]_0 (\grn_reg[5]_10 ),
        .\grn_reg[6] (\grn_reg[6]_9 ),
        .\grn_reg[6]_0 (\grn_reg[6]_10 ),
        .\grn_reg[7] (\grn_reg[7]_9 ),
        .\grn_reg[7]_0 (\grn_reg[7]_10 ),
        .\grn_reg[8] (\grn_reg[8]_9 ),
        .\grn_reg[8]_0 (\grn_reg[8]_10 ),
        .\grn_reg[9] (\grn_reg[9]_9 ),
        .\grn_reg[9]_0 (\grn_reg[9]_10 ),
        .\i_/bbus_o[4]_INST_0_i_22_0 (\i_/bbus_o[4]_INST_0_i_20_1 ),
        .\i_/bbus_o[4]_INST_0_i_22_1 (\i_/bbus_o[4]_INST_0_i_20_0 ),
        .\i_/bbus_o[4]_INST_0_i_23_0 (\i_/bbus_o[4]_INST_0_i_21_1 ),
        .\i_/bbus_o[5]_INST_0_i_16_0 (\sr[4]_i_197_5 [1:0]),
        .\i_/bdatw[15]_INST_0_i_35_0 (gr21),
        .\i_/bdatw[15]_INST_0_i_35_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_35_2 (\i_/bdatw[15]_INST_0_i_33 ),
        .\i_/bdatw[15]_INST_0_i_36_0 (gr26),
        .\i_/bdatw[15]_INST_0_i_36_1 (\i_/badr[15]_INST_0_i_52 ),
        .\i_/bdatw[15]_INST_0_i_36_2 (\i_/bdatw[15]_INST_0_i_34_0 ),
        .\i_/bdatw[15]_INST_0_i_36_3 (\i_/bbus_o[4]_INST_0_i_20 ),
        .\i_/bdatw[15]_INST_0_i_36_4 (\i_/bbus_o[4]_INST_0_i_21 ),
        .\i_/bdatw[15]_INST_0_i_36_5 (\i_/bbus_o[4]_INST_0_i_21_0 ),
        .\i_/bdatw[15]_INST_0_i_36_6 (gr25[15:5]),
        .\i_/bdatw[15]_INST_0_i_36_7 (\i_/bdatw[15]_INST_0_i_34 ),
        .\i_/bdatw[15]_INST_0_i_98_0 (\i_/bdatw[15]_INST_0_i_92 ),
        .out(gr27[15:5]));
  mcss_rgf_bank_bus_11 b1buso
       (.\bdatw[15]_INST_0_i_15 (gr07),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_6 ),
        .\grn_reg[0]_0 (\grn_reg[0]_7 ),
        .\grn_reg[0]_1 (\grn_reg[0]_8 ),
        .\grn_reg[10] (\grn_reg[10]_5 ),
        .\grn_reg[10]_0 (\grn_reg[10]_6 ),
        .\grn_reg[11] (\grn_reg[11]_5 ),
        .\grn_reg[11]_0 (\grn_reg[11]_6 ),
        .\grn_reg[12] (\grn_reg[12]_5 ),
        .\grn_reg[12]_0 (\grn_reg[12]_6 ),
        .\grn_reg[13] (\grn_reg[13]_5 ),
        .\grn_reg[13]_0 (\grn_reg[13]_6 ),
        .\grn_reg[14] (\grn_reg[14]_5 ),
        .\grn_reg[14]_0 (\grn_reg[14]_6 ),
        .\grn_reg[15] (\grn_reg[15]_11 ),
        .\grn_reg[1] (\grn_reg[1]_5 ),
        .\grn_reg[1]_0 (\grn_reg[1]_6 ),
        .\grn_reg[1]_1 (\grn_reg[1]_7 ),
        .\grn_reg[2] (\grn_reg[2]_5 ),
        .\grn_reg[2]_0 (\grn_reg[2]_6 ),
        .\grn_reg[2]_1 (\grn_reg[2]_7 ),
        .\grn_reg[3] (\grn_reg[3]_5 ),
        .\grn_reg[3]_0 (\grn_reg[3]_6 ),
        .\grn_reg[3]_1 (\grn_reg[3]_7 ),
        .\grn_reg[4] (\grn_reg[4]_11 ),
        .\grn_reg[4]_0 (\grn_reg[4]_12 ),
        .\grn_reg[4]_1 (\grn_reg[4]_13 ),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\grn_reg[6] (\grn_reg[6]_5 ),
        .\grn_reg[6]_0 (\grn_reg[6]_6 ),
        .\grn_reg[7] (\grn_reg[7]_5 ),
        .\grn_reg[7]_0 (\grn_reg[7]_6 ),
        .\grn_reg[8] (\grn_reg[8]_5 ),
        .\grn_reg[8]_0 (\grn_reg[8]_6 ),
        .\grn_reg[9] (\grn_reg[9]_5 ),
        .\grn_reg[9]_0 (\grn_reg[9]_6 ),
        .\i_/bdatw[15]_INST_0_i_121_0 (\i_/bdatw[15]_INST_0_i_121 ),
        .\i_/bdatw[15]_INST_0_i_121_1 (\i_/bdatw[15]_INST_0_i_121_0 ),
        .\i_/bdatw[15]_INST_0_i_121_2 (\i_/bdatw[15]_INST_0_i_121_1 ),
        .\i_/bdatw[15]_INST_0_i_124_0 (\i_/bdatw[15]_INST_0_i_124 ),
        .\i_/bdatw[15]_INST_0_i_124_1 (gr02),
        .\i_/bdatw[15]_INST_0_i_124_2 (gr01),
        .\i_/bdatw[15]_INST_0_i_212_0 (\sr[4]_i_197_5 [1:0]),
        .\i_/bdatw[15]_INST_0_i_212_1 (\i_/bdatw[15]_INST_0_i_212 ),
        .\i_/bdatw[15]_INST_0_i_48_0 (gr03),
        .\i_/bdatw[15]_INST_0_i_48_1 (gr04),
        .\i_/bdatw[15]_INST_0_i_48_2 (gr06),
        .\i_/bdatw[15]_INST_0_i_48_3 (gr05),
        .\i_/bdatw[8]_INST_0_i_69_0 (\i_/badr[15]_INST_0_i_135 ),
        .out(gr00));
  mcss_rgf_bank_bus_12 b1buso2l
       (.\bdatw[10]_INST_0_i_43 (\bdatw[10]_INST_0_i_43 ),
        .\bdatw[10]_INST_0_i_43_0 (\bdatw[10]_INST_0_i_43_0 ),
        .\bdatw[11]_INST_0_i_44 (\bdatw[11]_INST_0_i_44 ),
        .\bdatw[11]_INST_0_i_44_0 (\bdatw[11]_INST_0_i_44_0 ),
        .\bdatw[12]_INST_0_i_42 (\bdatw[12]_INST_0_i_42 ),
        .\bdatw[12]_INST_0_i_42_0 (\bdatw[12]_INST_0_i_42_0 ),
        .\bdatw[15]_INST_0_i_15 (gr27),
        .\bdatw[8]_INST_0_i_43 (\bdatw[8]_INST_0_i_43 ),
        .\bdatw[8]_INST_0_i_43_0 (\bdatw[8]_INST_0_i_43_0 ),
        .\bdatw[9]_INST_0_i_42 (\bdatw[9]_INST_0_i_42 ),
        .\bdatw[9]_INST_0_i_42_0 (\bdatw[9]_INST_0_i_42_0 ),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .\grn_reg[0] (\grn_reg[0]_15 ),
        .\grn_reg[0]_0 (\grn_reg[0]_16 ),
        .\grn_reg[10] (\grn_reg[10]_13 ),
        .\grn_reg[10]_0 (\grn_reg[10]_14 ),
        .\grn_reg[11] (\grn_reg[11]_13 ),
        .\grn_reg[11]_0 (\grn_reg[11]_14 ),
        .\grn_reg[12] (\grn_reg[12]_13 ),
        .\grn_reg[12]_0 (\grn_reg[12]_14 ),
        .\grn_reg[13] (\grn_reg[13]_13 ),
        .\grn_reg[13]_0 (\grn_reg[13]_14 ),
        .\grn_reg[14] (\grn_reg[14]_13 ),
        .\grn_reg[14]_0 (\grn_reg[14]_14 ),
        .\grn_reg[15] (\grn_reg[15]_18 ),
        .\grn_reg[1] (\grn_reg[1]_14 ),
        .\grn_reg[1]_0 (\grn_reg[1]_15 ),
        .\grn_reg[2] (\grn_reg[2]_14 ),
        .\grn_reg[2]_0 (\grn_reg[2]_15 ),
        .\grn_reg[3] (\grn_reg[3]_14 ),
        .\grn_reg[3]_0 (\grn_reg[3]_15 ),
        .\grn_reg[4] (\grn_reg[4]_20 ),
        .\grn_reg[4]_0 (\grn_reg[4]_21 ),
        .\grn_reg[5] (\grn_reg[5]_13 ),
        .\grn_reg[5]_0 (\grn_reg[5]_14 ),
        .\grn_reg[6] (\grn_reg[6]_13 ),
        .\grn_reg[6]_0 (\grn_reg[6]_14 ),
        .\grn_reg[7] (\grn_reg[7]_13 ),
        .\grn_reg[7]_0 (\grn_reg[7]_14 ),
        .\grn_reg[8] (\grn_reg[8]_13 ),
        .\grn_reg[8]_0 (\grn_reg[8]_14 ),
        .\grn_reg[9] (\grn_reg[9]_13 ),
        .\grn_reg[9]_0 (\grn_reg[9]_14 ),
        .\i_/bdatw[12]_INST_0_i_64_0 (\i_/badr[15]_INST_0_i_52 ),
        .\i_/bdatw[12]_INST_0_i_64_1 (\i_/bdatw[15]_INST_0_i_121 ),
        .\i_/bdatw[12]_INST_0_i_64_2 (\i_/bdatw[15]_INST_0_i_121_0 ),
        .\i_/bdatw[12]_INST_0_i_64_3 (\i_/bdatw[15]_INST_0_i_121_1 ),
        .\i_/bdatw[15]_INST_0_i_128_0 (\i_/bdatw[15]_INST_0_i_212 ),
        .\i_/bdatw[15]_INST_0_i_128_1 (gr22),
        .\i_/bdatw[15]_INST_0_i_128_2 (gr21),
        .\i_/bdatw[15]_INST_0_i_49_0 (gr25),
        .\i_/bdatw[15]_INST_0_i_49_1 (\sr[4]_i_197_5 [1:0]),
        .\i_/bdatw[15]_INST_0_i_49_2 (gr26[15:5]),
        .\i_/bdatw[15]_INST_0_i_49_3 (\i_/bdatw[15]_INST_0_i_124 ),
        .\i_/bdatw[15]_INST_0_i_49_4 (gr23),
        .\i_/bdatw[15]_INST_0_i_49_5 (gr24),
        .out(gr20[15:5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_7 
       (.I0(\grn_reg[0]_3 ),
        .I1(\grn_reg[0]_5 ),
        .I2(\badr[0]_INST_0_i_1 ),
        .I3(\grn_reg[0]_14 ),
        .I4(a1buso2l_n_32),
        .I5(\badr[0]_INST_0_i_1_0 ),
        .O(a1bus_b13[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_7 
       (.I0(\grn_reg[10]_3 ),
        .I1(a1buso_n_28),
        .I2(\badr[10]_INST_0_i_1 ),
        .I3(\grn_reg[10]_12 ),
        .I4(a1buso2l_n_12),
        .I5(\badr[10]_INST_0_i_1_0 ),
        .O(a1bus_b13[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_7 
       (.I0(\grn_reg[11]_3 ),
        .I1(a1buso_n_26),
        .I2(\badr[11]_INST_0_i_1 ),
        .I3(\grn_reg[11]_12 ),
        .I4(a1buso2l_n_10),
        .I5(\badr[11]_INST_0_i_1_0 ),
        .O(a1bus_b13[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_7 
       (.I0(\grn_reg[12]_3 ),
        .I1(a1buso_n_24),
        .I2(\badr[12]_INST_0_i_1 ),
        .I3(\grn_reg[12]_12 ),
        .I4(a1buso2l_n_8),
        .I5(\badr[12]_INST_0_i_1_0 ),
        .O(a1bus_b13[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_7 
       (.I0(\grn_reg[13]_3 ),
        .I1(a1buso_n_22),
        .I2(\badr[13]_INST_0_i_1 ),
        .I3(\grn_reg[13]_12 ),
        .I4(a1buso2l_n_6),
        .I5(\badr[13]_INST_0_i_1_0 ),
        .O(a1bus_b13[13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_7 
       (.I0(\grn_reg[14]_3 ),
        .I1(a1buso_n_20),
        .I2(\badr[14]_INST_0_i_1 ),
        .I3(\grn_reg[14]_12 ),
        .I4(a1buso2l_n_4),
        .I5(\badr[14]_INST_0_i_1_0 ),
        .O(a1bus_b13[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_7 
       (.I0(\grn_reg[15]_8 ),
        .I1(\grn_reg[15]_10 ),
        .I2(\badr[15]_INST_0_i_1_0 ),
        .I3(\grn_reg[15]_17 ),
        .I4(a1buso2l_n_2),
        .I5(\badr[15]_INST_0_i_1_1 ),
        .O(a1bus_b13[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_7 
       (.I0(\grn_reg[1]_3 ),
        .I1(a1buso_n_46),
        .I2(\badr[1]_INST_0_i_1 ),
        .I3(\grn_reg[1]_13 ),
        .I4(a1buso2l_n_30),
        .I5(\badr[1]_INST_0_i_1_0 ),
        .O(a1bus_b13[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_7 
       (.I0(\grn_reg[2]_3 ),
        .I1(a1buso_n_44),
        .I2(\badr[2]_INST_0_i_1 ),
        .I3(\grn_reg[2]_13 ),
        .I4(a1buso2l_n_28),
        .I5(\badr[2]_INST_0_i_1_0 ),
        .O(a1bus_b13[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_7 
       (.I0(\grn_reg[3]_3 ),
        .I1(a1buso_n_42),
        .I2(\badr[3]_INST_0_i_1 ),
        .I3(\grn_reg[3]_13 ),
        .I4(a1buso2l_n_26),
        .I5(\badr[3]_INST_0_i_1_0 ),
        .O(a1bus_b13[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_7 
       (.I0(\grn_reg[4]_9 ),
        .I1(a1buso_n_40),
        .I2(\badr[4]_INST_0_i_1 ),
        .I3(\grn_reg[4]_19 ),
        .I4(a1buso2l_n_24),
        .I5(\badr[4]_INST_0_i_1_0 ),
        .O(a1bus_b13[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_7 
       (.I0(\grn_reg[5]_3 ),
        .I1(a1buso_n_38),
        .I2(\badr[5]_INST_0_i_1 ),
        .I3(\grn_reg[5]_12 ),
        .I4(a1buso2l_n_22),
        .I5(\badr[5]_INST_0_i_1_0 ),
        .O(a1bus_b13[5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_7 
       (.I0(\grn_reg[6]_3 ),
        .I1(a1buso_n_36),
        .I2(\badr[6]_INST_0_i_1 ),
        .I3(\grn_reg[6]_12 ),
        .I4(a1buso2l_n_20),
        .I5(\badr[6]_INST_0_i_1_0 ),
        .O(a1bus_b13[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_7 
       (.I0(\grn_reg[7]_3 ),
        .I1(a1buso_n_34),
        .I2(\badr[7]_INST_0_i_1 ),
        .I3(\grn_reg[7]_12 ),
        .I4(a1buso2l_n_18),
        .I5(\badr[7]_INST_0_i_1_0 ),
        .O(a1bus_b13[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_7 
       (.I0(\grn_reg[8]_3 ),
        .I1(a1buso_n_32),
        .I2(\badr[8]_INST_0_i_1 ),
        .I3(\grn_reg[8]_12 ),
        .I4(a1buso2l_n_16),
        .I5(\badr[8]_INST_0_i_1_0 ),
        .O(a1bus_b13[8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_7 
       (.I0(\grn_reg[9]_3 ),
        .I1(a1buso_n_30),
        .I2(\badr[9]_INST_0_i_1 ),
        .I3(\grn_reg[9]_12 ),
        .I4(a1buso2l_n_14),
        .I5(\badr[9]_INST_0_i_1_0 ),
        .O(a1bus_b13[9]));
  mcss_rgf_grn grn00
       (.Q(gr00),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_19 ),
        .\grn_reg[15]_1 (\grn_reg[15]_20 ));
  mcss_rgf_grn_13 grn01
       (.Q(gr01),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_21 ),
        .\grn_reg[15]_1 (\grn_reg[15]_22 ));
  mcss_rgf_grn_14 grn02
       (.Q(gr02),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_23 ),
        .\grn_reg[15]_1 (\grn_reg[15]_24 ));
  mcss_rgf_grn_15 grn03
       (.Q(gr03),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_25 ),
        .\grn_reg[15]_1 (\grn_reg[15]_26 ));
  mcss_rgf_grn_16 grn04
       (.Q(gr04),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_27 ),
        .\grn_reg[15]_1 (\grn_reg[15]_28 ));
  mcss_rgf_grn_17 grn05
       (.Q(gr05),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_29 ),
        .\grn_reg[15]_1 (\grn_reg[15]_30 ));
  mcss_rgf_grn_18 grn06
       (.Q(gr06),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_31 ),
        .\grn_reg[15]_1 (\grn_reg[15]_32 ));
  mcss_rgf_grn_19 grn07
       (.Q(gr07),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_33 ),
        .\grn_reg[15]_1 (\grn_reg[15]_34 ));
  mcss_rgf_grn_20 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_35 ),
        .\grn_reg[15]_1 (\grn_reg[15]_36 ));
  mcss_rgf_grn_21 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_37 ),
        .\grn_reg[15]_1 (\grn_reg[15]_38 ));
  mcss_rgf_grn_22 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_39 ),
        .\grn_reg[15]_1 (\grn_reg[15]_40 ));
  mcss_rgf_grn_23 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_41 ),
        .\grn_reg[15]_1 (\grn_reg[15]_42 ));
  mcss_rgf_grn_24 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_43 ),
        .\grn_reg[15]_1 (\grn_reg[15]_44 ));
  mcss_rgf_grn_25 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_45 ),
        .\grn_reg[15]_1 (\grn_reg[15]_46 ));
  mcss_rgf_grn_26 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_47 ),
        .\grn_reg[15]_1 (\grn_reg[15]_48 ));
  mcss_rgf_grn_27 grn27
       (.Q(gr27),
        .SR(SR),
        .clk(clk),
        .fdat(fdat),
        .\fdat[15] (\fdat[15] ),
        .fdat_12_sp_1(fdat_12_sn_1),
        .fdatx(fdatx),
        .\fdatx[15] (\fdatx[15] ),
        .\grn_reg[15]_0 (\grn_reg[15]_49 ),
        .\grn_reg[15]_1 (\grn_reg[15]_50 ),
        .\ir0_id_fl[20]_i_4_0 (\ir0_id_fl[20]_i_4 ),
        .\nir_id_reg[20] (\nir_id_reg[20] ),
        .\rgf_c1bus_wb[14]_i_28 (\rgf_c1bus_wb[14]_i_28 ),
        .\rgf_c1bus_wb[4]_i_11 ({\rgf_c1bus_wb[4]_i_11 [12],\rgf_c1bus_wb[4]_i_11 [1]}),
        .\rgf_c1bus_wb[4]_i_11_0 (\sr[4]_i_170_0 ),
        .\rgf_c1bus_wb[4]_i_11_1 (\sr[4]_i_168_1 ),
        .\rgf_c1bus_wb[4]_i_11_2 (\rgf_c1bus_wb[4]_i_11_2 ),
        .\rgf_c1bus_wb[4]_i_11_3 (\rgf_c1bus_wb[4]_i_11_3 ),
        .\rgf_c1bus_wb[4]_i_11_4 (\rgf_c1bus_wb[4]_i_11_4 ),
        .\rgf_c1bus_wb[4]_i_13 (\sr[4]_i_164_0 ),
        .\rgf_c1bus_wb[4]_i_13_0 (\sr[4]_i_170 ),
        .\rgf_c1bus_wb[4]_i_13_1 (\sr[4]_i_155_1 ),
        .\rgf_c1bus_wb[4]_i_13_2 (\sr[4]_i_170_3 ),
        .\rgf_c1bus_wb[4]_i_4 (\rgf_c1bus_wb[4]_i_25_n_0 ),
        .\rgf_c1bus_wb[4]_i_4_0 (\rgf_c1bus_wb[4]_i_26_n_0 ),
        .\rgf_c1bus_wb[4]_i_4_1 (\sr[4]_i_80_2 ),
        .\rgf_c1bus_wb[4]_i_4_2 (\rgf_c1bus_wb[4]_i_27_n_0 ),
        .\rgf_c1bus_wb[4]_i_4_3 (\rgf_c1bus_wb[4]_i_28_n_0 ),
        .\rgf_c1bus_wb[4]_i_4_4 (\sr[4]_i_80_0 ),
        .rst_n(rst_n),
        .\tr_reg[14] (\tr_reg[14] ),
        .\tr_reg[1] (\tr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[12]_i_24 
       (.I0(\sr[4]_i_186_0 ),
        .I1(\sr[4]_i_186_1 ),
        .I2(\sr[4]_i_183_2 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[15]_i_23_3 ),
        .I5(\sr[4]_i_183_3 ),
        .O(\sp_reg[6] ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c0bus_wb[13]_i_27 
       (.I0(\rgf_c0bus_wb[13]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_31_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[13]_i_32_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[13]_i_13 ),
        .O(\sr_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[13]_i_30 
       (.I0(\sr[4]_i_183_7 ),
        .I1(\sr[4]_i_183_8 ),
        .I2(\sr[4]_i_183_1 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_183_12 ),
        .I5(\sr[4]_i_183_5 ),
        .O(\rgf_c0bus_wb[13]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[13]_i_31 
       (.I0(\sr[4]_i_183_16 ),
        .I1(\sr[4]_i_183_17 ),
        .I2(\sr[4]_i_183_3 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_183_9 ),
        .I5(\sr[4]_i_183_0 ),
        .O(\rgf_c0bus_wb[13]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[13]_i_32 
       (.I0(\sr[4]_i_183_10 ),
        .I1(\sr[4]_i_183_11 ),
        .I2(\sr[4]_i_183_6 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_183_19 ),
        .I5(\sr[4]_i_183_4 ),
        .O(\rgf_c0bus_wb[13]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[15]_i_21 
       (.I0(\rgf_c0bus_wb[4]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_29_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[4]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_31_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[15]_i_23 
       (.I0(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[4]_i_30_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .O(\sr_reg[6]_3 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[15]_i_27 
       (.I0(\sr[4]_i_194_0 ),
        .I1(\sr[4]_i_194_1 ),
        .I2(\sr[4]_i_197_7 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_194_2 ),
        .I5(\sr[4]_i_197_2 ),
        .O(\rgf_c0bus_wb[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[15]_i_28 
       (.I0(\sr[4]_i_197_3 ),
        .I1(\sr[4]_i_197_4 ),
        .I2(\sr[4]_i_183_4 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[15]_i_23_6 ),
        .I5(\sr[4]_i_183_6 ),
        .O(\rgf_c0bus_wb[15]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h010001FF)) 
    \rgf_c0bus_wb[15]_i_29 
       (.I0(\rgf_c0bus_wb[15]_i_23_8 ),
        .I1(\rgf_c0bus_wb[15]_i_23_9 ),
        .I2(\rgf_c0bus_wb[15]_i_23_7 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_197_5 [2]),
        .O(\rgf_c0bus_wb[15]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[15]_i_30 
       (.I0(\rgf_c0bus_wb[15]_i_23_4 ),
        .I1(\rgf_c0bus_wb[15]_i_23_5 ),
        .I2(\sr[4]_i_183_5 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[15]_i_23_2 ),
        .I5(\sr[4]_i_183_1 ),
        .O(\rgf_c0bus_wb[15]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[4]_i_11 
       (.I0(\rgf_c0bus_wb[4]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_30_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[4]_i_31_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[4]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_32_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_23_4 ),
        .I1(\rgf_c0bus_wb[15]_i_23_5 ),
        .I2(\sr[4]_i_183_5 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[15]_i_23_6 ),
        .I5(\sr[4]_i_183_6 ),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_19 
       (.I0(\rgf_c0bus_wb[15]_i_23_0 ),
        .I1(\rgf_c0bus_wb[15]_i_23_1 ),
        .I2(\sr[4]_i_183_0 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[15]_i_23_2 ),
        .I5(\sr[4]_i_183_1 ),
        .O(\sp_reg[4] ));
  LUT5 #(
    .INIT(32'h010001FF)) 
    \rgf_c0bus_wb[4]_i_22 
       (.I0(\sr[4]_i_197_3 ),
        .I1(\sr[4]_i_197_4 ),
        .I2(\sr[4]_i_183_4 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_197_5 [2]),
        .O(\rgf_c0bus_wb[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_23 
       (.I0(\rgf_c0bus_wb[4]_i_8_2 ),
        .I1(\rgf_c0bus_wb[4]_i_8_3 ),
        .I2(\rgf_c0bus_wb[4]_i_8_4 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[4]_i_8_8 ),
        .I5(\rgf_c0bus_wb[4]_i_8_9 ),
        .O(\rgf_c0bus_wb[4]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_24 
       (.I0(\sr[4]_i_197_0 ),
        .I1(\sr[4]_i_197_1 ),
        .I2(\sr[4]_i_197_2 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_197_6 ),
        .I5(\sr[4]_i_197_7 ),
        .O(\rgf_c0bus_wb[4]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_25 
       (.I0(\sr[4]_i_183_13 ),
        .I1(\sr[4]_i_183_14 ),
        .I2(\sr[4]_i_183_15 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_183_18 ),
        .I5(\sr[4]_i_183_2 ),
        .O(\rgf_c0bus_wb[4]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_26 
       (.I0(\rgf_c0bus_wb[4]_i_8_5 ),
        .I1(\rgf_c0bus_wb[4]_i_8_6 ),
        .I2(\rgf_c0bus_wb[4]_i_8_7 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[4]_i_8_0 ),
        .I5(\rgf_c0bus_wb[4]_i_8_1 ),
        .O(\rgf_c0bus_wb[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_27 
       (.I0(\sr[4]_i_183_10 ),
        .I1(\sr[4]_i_183_11 ),
        .I2(\sr[4]_i_183_6 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_183_12 ),
        .I5(\sr[4]_i_183_5 ),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_29 
       (.I0(\sr[4]_i_186_0 ),
        .I1(\sr[4]_i_186_1 ),
        .I2(\sr[4]_i_183_2 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_186_5 ),
        .I5(\sr[4]_i_183_15 ),
        .O(\rgf_c0bus_wb[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_30 
       (.I0(\rgf_c0bus_wb[15]_i_23_0 ),
        .I1(\rgf_c0bus_wb[15]_i_23_1 ),
        .I2(\sr[4]_i_183_0 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[15]_i_23_3 ),
        .I5(\sr[4]_i_183_3 ),
        .O(\rgf_c0bus_wb[4]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_31 
       (.I0(\sr[4]_i_194_3 ),
        .I1(\sr[4]_i_194_4 ),
        .I2(\rgf_c0bus_wb[4]_i_8_9 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_194_5 ),
        .I5(\rgf_c0bus_wb[4]_i_8_4 ),
        .O(\rgf_c0bus_wb[4]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_32 
       (.I0(\sr[4]_i_186_2 ),
        .I1(\sr[4]_i_186_3 ),
        .I2(\rgf_c0bus_wb[4]_i_8_1 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_186_4 ),
        .I5(\rgf_c0bus_wb[4]_i_8_7 ),
        .O(\rgf_c0bus_wb[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c0bus_wb[4]_i_33 
       (.I0(\rgf_c0bus_wb[4]_i_12_0 ),
        .I1(\rgf_c0bus_wb[4]_i_12_1 ),
        .I2(\rgf_c0bus_wb[4]_i_12 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[4]_i_12_2 ),
        .I5(\rgf_c0bus_wb[15]_i_23_7 ),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[4]_i_7 
       (.I0(\sp_reg[2] ),
        .I1(\sp_reg[4] ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[12]_i_7 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[4]_i_22_n_0 ),
        .O(\sr_reg[6]_5 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[4]_i_8 
       (.I0(\rgf_c0bus_wb[4]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_24_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[4]_i_25_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[4]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_26_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_24 
       (.I0(\rgf_c1bus_wb[4]_i_11_1 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [10]),
        .I2(\rgf_c1bus_wb[4]_i_11_5 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\rgf_c1bus_wb[4]_i_11_0 ),
        .I5(\rgf_c1bus_wb[4]_i_11_6 ),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_25 
       (.I0(\sr[4]_i_155_2 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [4]),
        .I2(\sr[4]_i_155_3 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_155_4 ),
        .I5(\sr[4]_i_155_5 ),
        .O(\rgf_c1bus_wb[4]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_26 
       (.I0(\sr[4]_i_155_8 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [5]),
        .I2(\sr[4]_i_155_9 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_155_10 ),
        .I5(\sr[4]_i_155_11 ),
        .O(\rgf_c1bus_wb[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_27 
       (.I0(\sr[4]_i_159_3 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [6]),
        .I2(\sr[4]_i_159_4 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_159_1 ),
        .I5(\sr[4]_i_159_5 ),
        .O(\rgf_c1bus_wb[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_28 
       (.I0(\sr[4]_i_159_2 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [8]),
        .I2(\sr[4]_i_159_6 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_159_0 ),
        .I5(\sr[4]_i_159_7 ),
        .O(\rgf_c1bus_wb[4]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h1100030311330303)) 
    \sr[4]_i_130 
       (.I0(\sr[4]_i_190_n_0 ),
        .I1(\sr[4]_i_57_2 ),
        .I2(\rgf_c0bus_wb[4]_i_26_0 ),
        .I3(\sr[4]_i_66_0 ),
        .I4(\sr[4]_i_57_1 ),
        .I5(\sr_reg[6]_1 ),
        .O(\sr[4]_i_130_n_0 ));
  LUT6 #(
    .INIT(64'h3030505F0F0F0F0F)) 
    \sr[4]_i_131 
       (.I0(\rgf_c0bus_wb[4]_i_26_0 ),
        .I1(\sr[4]_i_190_n_0 ),
        .I2(\sr[4]_i_15_0 ),
        .I3(\sr[4]_i_57_0 ),
        .I4(\sr[4]_i_57_1 ),
        .I5(\sr[4]_i_57_2 ),
        .O(\sr[4]_i_131_n_0 ));
  LUT6 #(
    .INIT(64'hCCECCFECCCEFCFEF)) 
    \sr[4]_i_133 
       (.I0(\sr[4]_i_57_3 ),
        .I1(\sr[4]_i_66 ),
        .I2(\sr[4]_i_66_0 ),
        .I3(\sr[4]_i_57_1 ),
        .I4(\rgf_c0bus_wb[4]_i_32_0 ),
        .I5(\sr[4]_i_191_n_0 ),
        .O(\sr[4]_i_133_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCEECFCCFFEECF)) 
    \sr[4]_i_138 
       (.I0(\sr[4]_i_193_n_0 ),
        .I1(\sr[4]_i_66 ),
        .I2(\sr[4]_i_194_n_0 ),
        .I3(\sr[4]_i_66_0 ),
        .I4(\sr[4]_i_57_1 ),
        .I5(\sr[4]_i_195_n_0 ),
        .O(\sr[4]_i_195_0 ));
  LUT6 #(
    .INIT(64'hCCFCEECCCCFCEEFF)) 
    \sr[4]_i_142 
       (.I0(\sr[4]_i_198_n_0 ),
        .I1(\sr[4]_i_66 ),
        .I2(\sr[4]_i_199_n_0 ),
        .I3(\sr[4]_i_66_0 ),
        .I4(\sr[4]_i_57_1 ),
        .I5(\sr[4]_i_200_n_0 ),
        .O(\sr[4]_i_200_0 ));
  LUT5 #(
    .INIT(32'hC005CF05)) 
    \sr[4]_i_148 
       (.I0(\sr[4]_i_190_n_0 ),
        .I1(\sr[4]_i_67 ),
        .I2(\sr[4]_i_57_1 ),
        .I3(\sr[4]_i_67_0 ),
        .I4(\sr_reg[6]_1 ),
        .O(\rgf_c0bus_wb[13]_i_27_0 ));
  LUT6 #(
    .INIT(64'h55335533FF0F000F)) 
    \sr[4]_i_154 
       (.I0(\tr_reg[11] ),
        .I1(\sr[4]_i_208_n_0 ),
        .I2(\tr_reg[13] ),
        .I3(\sr[4]_i_80_0 ),
        .I4(\sr[4]_i_80_1 ),
        .I5(\sr[4]_i_80_2 ),
        .O(\sr[4]_i_154_n_0 ));
  LUT6 #(
    .INIT(64'h000FFF0F33553355)) 
    \sr[4]_i_155 
       (.I0(\rgf_c1bus_wb[4]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_26_n_0 ),
        .I2(\sr[4]_i_210_n_0 ),
        .I3(\sr[4]_i_80_0 ),
        .I4(\sr[4]_i_211_n_0 ),
        .I5(\sr[4]_i_80_2 ),
        .O(\sr[4]_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_156 
       (.I0(\tr_reg[11] ),
        .I1(\sr[4]_i_208_n_0 ),
        .I2(\sr[4]_i_80_2 ),
        .I3(\sr[4]_i_83 ),
        .I4(\sr[4]_i_80_0 ),
        .I5(\tr_reg[13] ),
        .O(\sr[4]_i_156_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_159 
       (.I0(\rgf_c1bus_wb[4]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_26_n_0 ),
        .I2(\sr[4]_i_80_2 ),
        .I3(\tr_reg[12] ),
        .I4(\sr[4]_i_80_0 ),
        .I5(\rgf_c1bus_wb[4]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_28_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \sr[4]_i_160 
       (.I0(\rgf_c1bus_wb[4]_i_25_n_0 ),
        .I1(\sr[4]_i_211_n_0 ),
        .I2(\sr[4]_i_210_n_0 ),
        .I3(\sr[4]_i_80_0 ),
        .I4(\sr[4]_i_83 ),
        .I5(\sr[4]_i_80_2 ),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \sr[4]_i_164 
       (.I0(\tr_reg[11] ),
        .I1(\tr_reg[13] ),
        .I2(\sr[4]_i_80_2 ),
        .I3(\sr[4]_i_210_n_0 ),
        .I4(\sr[4]_i_80_0 ),
        .I5(\sr[4]_i_83 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hE2FFE200E2FFE2FF)) 
    \sr[4]_i_166 
       (.I0(\tr_reg[11] ),
        .I1(\sr[4]_i_80_0 ),
        .I2(\tr_reg[13] ),
        .I3(\sr[4]_i_80_2 ),
        .I4(\sr[4]_i_90 ),
        .I5(\sr[4]_i_80_1 ),
        .O(\badr[15]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_183 
       (.I0(\rgf_c0bus_wb[13]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_25_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[13]_i_32_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[13]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_30_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_186 
       (.I0(\rgf_c0bus_wb[4]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[4]_i_32_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[4]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_29_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_187 
       (.I0(\sp_reg[13] ),
        .I1(\sp_reg[11] ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .O(\sr_reg[6]_4 ));
  LUT6 #(
    .INIT(64'hB8FFB800B8FFB8FF)) 
    \sr[4]_i_189 
       (.I0(\sp_reg[13] ),
        .I1(\sr[4]_i_139_0 ),
        .I2(\sp_reg[11] ),
        .I3(\sr[4]_i_139 ),
        .I4(\sr[4]_i_129 ),
        .I5(\sr[4]_i_138_1 ),
        .O(\badr[15]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \sr[4]_i_190 
       (.I0(\rgf_c0bus_wb[13]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_31_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\sr[4]_i_139_0 ),
        .I4(\rgf_c0bus_wb[13]_i_32_n_0 ),
        .O(\sr[4]_i_190_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_191 
       (.I0(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I1(\sp_reg[13] ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .O(\sr[4]_i_191_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \sr[4]_i_192 
       (.I0(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_31_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\sr[4]_i_139_0 ),
        .I4(\sp_reg[14] ),
        .O(\rgf_c0bus_wb[4]_i_33_0 ));
  LUT6 #(
    .INIT(64'h00A30FA3F0A3FFA3)) 
    \sr[4]_i_193 
       (.I0(\sr[4]_i_138_1 ),
        .I1(\sp_reg[14] ),
        .I2(\sr[4]_i_139_0 ),
        .I3(\sr[4]_i_139 ),
        .I4(\rgf_c0bus_wb[4]_i_31_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .O(\sr[4]_i_193_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_194 
       (.I0(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_31_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\sr[4]_i_138_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\sp_reg[14] ),
        .O(\sr[4]_i_194_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_195 
       (.I0(\sr[4]_i_229_n_0 ),
        .I1(\sp_reg[1] ),
        .I2(\sr[4]_i_139 ),
        .I3(\sr[4]_i_230_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\sr[4]_i_231_n_0 ),
        .O(\sr[4]_i_195_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_197 
       (.I0(\rgf_c0bus_wb[4]_i_22_n_0 ),
        .I1(\sp_reg[2] ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[4]_i_24_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\rgf_c0bus_wb[12]_i_7 ),
        .O(\sr_reg[6]_2 ));
  LUT6 #(
    .INIT(64'h5F5030305F503F3F)) 
    \sr[4]_i_198 
       (.I0(\sp_reg[11] ),
        .I1(\sr[4]_i_232_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\sr[4]_i_138_1 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\sp_reg[13] ),
        .O(\sr[4]_i_198_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \sr[4]_i_199 
       (.I0(\rgf_c0bus_wb[4]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I3(\sr[4]_i_139_0 ),
        .I4(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I5(\sr[4]_i_139 ),
        .O(\sr[4]_i_199_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_200 
       (.I0(\sp_reg[11] ),
        .I1(\sr[4]_i_232_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\sp_reg[13] ),
        .O(\sr[4]_i_200_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_202 
       (.I0(\sr[4]_i_230_n_0 ),
        .I1(\sr[4]_i_231_n_0 ),
        .I2(\sr[4]_i_139 ),
        .I3(\sp_reg[11] ),
        .I4(\sr[4]_i_139_0 ),
        .I5(\sr[4]_i_232_n_0 ),
        .O(\sr[4]_i_232_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_207 
       (.I0(\sr[4]_i_159_0 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [9]),
        .I2(\sr[4]_i_168_3 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\rgf_c1bus_wb[4]_i_11_1 ),
        .I5(\sr[4]_i_168_0 ),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_208 
       (.I0(\sr[4]_i_159_1 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [7]),
        .I2(\sr[4]_i_154_0 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_159_2 ),
        .I5(\sr[4]_i_154_1 ),
        .O(\sr[4]_i_208_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_209 
       (.I0(\rgf_c1bus_wb[4]_i_11_0 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [11]),
        .I2(\sr[4]_i_168 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_168_1 ),
        .I5(\sr[4]_i_168_2 ),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_210 
       (.I0(\sr[4]_i_164_1 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [0]),
        .I2(\sr[4]_i_164_2 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_164_0 ),
        .I5(\sr[4]_i_164_3 ),
        .O(\sr[4]_i_210_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_211 
       (.I0(\sr[4]_i_155_1 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [2]),
        .I2(\sr[4]_i_155_6 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_155_0 ),
        .I5(\sr[4]_i_155_7 ),
        .O(\sr[4]_i_211_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_213 
       (.I0(\sr[4]_i_164_0 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [1]),
        .I2(\sr[4]_i_170 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_164_1 ),
        .I5(\sr[4]_i_170_1 ),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_220 
       (.I0(\sr[4]_i_155_0 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [3]),
        .I2(\sr[4]_i_170_2 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\sr[4]_i_155_1 ),
        .I5(\sr[4]_i_170_3 ),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_223 
       (.I0(\rgf_c1bus_wb[4]_i_11_0 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [11]),
        .I2(\sr[4]_i_168 ),
        .I3(\sr[4]_i_170_0 ),
        .I4(\rgf_c1bus_wb[4]_i_11_1 ),
        .I5(\sr[4]_i_168_0 ),
        .O(\tr_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_227 
       (.I0(\sr[4]_i_197_0 ),
        .I1(\sr[4]_i_197_1 ),
        .I2(\sr[4]_i_197_2 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_185_0 ),
        .I5(\rgf_c0bus_wb[4]_i_12 ),
        .O(\sp_reg[13] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_228 
       (.I0(\rgf_c0bus_wb[4]_i_8_2 ),
        .I1(\rgf_c0bus_wb[4]_i_8_3 ),
        .I2(\rgf_c0bus_wb[4]_i_8_4 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_197_6 ),
        .I5(\sr[4]_i_197_7 ),
        .O(\sp_reg[11] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_229 
       (.I0(\sr[4]_i_183_7 ),
        .I1(\sr[4]_i_183_8 ),
        .I2(\sr[4]_i_183_1 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_183_9 ),
        .I5(\sr[4]_i_183_0 ),
        .O(\sr[4]_i_229_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_230 
       (.I0(\sr[4]_i_183_13 ),
        .I1(\sr[4]_i_183_14 ),
        .I2(\sr[4]_i_183_15 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[4]_i_8_0 ),
        .I5(\rgf_c0bus_wb[4]_i_8_1 ),
        .O(\sr[4]_i_230_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_231 
       (.I0(\sr[4]_i_183_16 ),
        .I1(\sr[4]_i_183_17 ),
        .I2(\sr[4]_i_183_3 ),
        .I3(\sr[4]_i_185 ),
        .I4(\sr[4]_i_183_18 ),
        .I5(\sr[4]_i_183_2 ),
        .O(\sr[4]_i_231_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \sr[4]_i_232 
       (.I0(\rgf_c0bus_wb[4]_i_8_5 ),
        .I1(\rgf_c0bus_wb[4]_i_8_6 ),
        .I2(\rgf_c0bus_wb[4]_i_8_7 ),
        .I3(\sr[4]_i_185 ),
        .I4(\rgf_c0bus_wb[4]_i_8_8 ),
        .I5(\rgf_c0bus_wb[4]_i_8_9 ),
        .O(\sr[4]_i_232_n_0 ));
  LUT6 #(
    .INIT(64'hE000E0E0E000E000)) 
    \sr[4]_i_57 
       (.I0(\sr[4]_i_130_n_0 ),
        .I1(\sr[4]_i_131_n_0 ),
        .I2(\sr[4]_i_15 ),
        .I3(\sr[4]_i_15_0 ),
        .I4(\sr[4]_i_15_1 ),
        .I5(\sr[4]_i_133_n_0 ),
        .O(\sr[4]_i_133_0 ));
  LUT6 #(
    .INIT(64'hEECCCCFCEECCFFFC)) 
    \sr[4]_i_80 
       (.I0(\sr[4]_i_154_n_0 ),
        .I1(\sr[4]_i_27 ),
        .I2(\sr[4]_i_155_n_0 ),
        .I3(\sr[4]_i_27_0 ),
        .I4(\sr[4]_i_27_1 ),
        .I5(\sr[4]_i_156_n_0 ),
        .O(\sr[4]_i_156_0 ));
endmodule

module mcss_rgf_bank_bus
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[15]_INST_0_i_12 ,
    \i_/badr[15]_INST_0_i_55_0 ,
    a0bus_sel_0,
    \badr[15]_INST_0_i_12_0 ,
    \badr[15]_INST_0_i_12_1 ,
    \i_/badr[15]_INST_0_i_54_0 ,
    \i_/badr[15]_INST_0_i_54_1 ,
    \i_/badr[15]_INST_0_i_135_0 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_135_1 ,
    ctl_sela0,
    \i_/badr[15]_INST_0_i_135_2 ,
    \i_/badr[15]_INST_0_i_55_1 ,
    \i_/badr[15]_INST_0_i_55_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_12 ;
  input [1:0]\i_/badr[15]_INST_0_i_55_0 ;
  input [3:0]a0bus_sel_0;
  input [15:0]\badr[15]_INST_0_i_12_0 ;
  input [15:0]\badr[15]_INST_0_i_12_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_54_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_54_1 ;
  input \i_/badr[15]_INST_0_i_135_0 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_135_1 ;
  input [0:0]ctl_sela0;
  input \i_/badr[15]_INST_0_i_135_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_55_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_55_2 ;

  wire [3:0]a0bus_sel_0;
  wire [15:0]\badr[15]_INST_0_i_12 ;
  wire [15:0]\badr[15]_INST_0_i_12_0 ;
  wire [15:0]\badr[15]_INST_0_i_12_1 ;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_42_n_0 ;
  wire \i_/badr[0]_INST_0_i_43_n_0 ;
  wire \i_/badr[10]_INST_0_i_40_n_0 ;
  wire \i_/badr[10]_INST_0_i_41_n_0 ;
  wire \i_/badr[11]_INST_0_i_45_n_0 ;
  wire \i_/badr[11]_INST_0_i_46_n_0 ;
  wire \i_/badr[12]_INST_0_i_40_n_0 ;
  wire \i_/badr[12]_INST_0_i_41_n_0 ;
  wire \i_/badr[13]_INST_0_i_40_n_0 ;
  wire \i_/badr[13]_INST_0_i_41_n_0 ;
  wire \i_/badr[14]_INST_0_i_40_n_0 ;
  wire \i_/badr[14]_INST_0_i_41_n_0 ;
  wire \i_/badr[15]_INST_0_i_135_0 ;
  wire \i_/badr[15]_INST_0_i_135_1 ;
  wire \i_/badr[15]_INST_0_i_135_2 ;
  wire \i_/badr[15]_INST_0_i_135_n_0 ;
  wire \i_/badr[15]_INST_0_i_138_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_54_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_54_1 ;
  wire [1:0]\i_/badr[15]_INST_0_i_55_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_55_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_55_2 ;
  wire \i_/badr[1]_INST_0_i_40_n_0 ;
  wire \i_/badr[1]_INST_0_i_41_n_0 ;
  wire \i_/badr[2]_INST_0_i_40_n_0 ;
  wire \i_/badr[2]_INST_0_i_41_n_0 ;
  wire \i_/badr[3]_INST_0_i_44_n_0 ;
  wire \i_/badr[3]_INST_0_i_45_n_0 ;
  wire \i_/badr[4]_INST_0_i_40_n_0 ;
  wire \i_/badr[4]_INST_0_i_41_n_0 ;
  wire \i_/badr[5]_INST_0_i_40_n_0 ;
  wire \i_/badr[5]_INST_0_i_41_n_0 ;
  wire \i_/badr[6]_INST_0_i_40_n_0 ;
  wire \i_/badr[6]_INST_0_i_41_n_0 ;
  wire \i_/badr[7]_INST_0_i_45_n_0 ;
  wire \i_/badr[7]_INST_0_i_46_n_0 ;
  wire \i_/badr[8]_INST_0_i_40_n_0 ;
  wire \i_/badr[8]_INST_0_i_41_n_0 ;
  wire \i_/badr[9]_INST_0_i_40_n_0 ;
  wire \i_/badr[9]_INST_0_i_41_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [0]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_42_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [0]),
        .I4(\i_/badr[0]_INST_0_i_43_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [10]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_40_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [10]),
        .I4(\i_/badr[10]_INST_0_i_41_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [11]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_45_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [11]),
        .I4(\i_/badr[11]_INST_0_i_46_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_46 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [12]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_40_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [12]),
        .I4(\i_/badr[12]_INST_0_i_41_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [13]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_40_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [13]),
        .I4(\i_/badr[13]_INST_0_i_41_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [14]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_40_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [14]),
        .I4(\i_/badr[14]_INST_0_i_41_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_133 
       (.I0(\i_/badr[15]_INST_0_i_55_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_55_0 [0]),
        .I2(a0bus_sel_0[3]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_134 
       (.I0(\i_/badr[15]_INST_0_i_55_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_55_0 [0]),
        .I2(a0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_135 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_135_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_136 
       (.I0(\i_/badr[15]_INST_0_i_55_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_55_0 [0]),
        .I2(a0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_137 
       (.I0(\i_/badr[15]_INST_0_i_55_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_55_0 [0]),
        .I2(a0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_138 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_138_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_220 
       (.I0(\i_/badr[15]_INST_0_i_135_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\i_/badr[15]_INST_0_i_135_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_135_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_221 
       (.I0(\i_/badr[15]_INST_0_i_135_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\i_/badr[15]_INST_0_i_135_1 ),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_135_2 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_222 
       (.I0(\i_/badr[15]_INST_0_i_135_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\i_/badr[15]_INST_0_i_135_1 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_135_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_223 
       (.I0(\i_/badr[15]_INST_0_i_135_0 ),
        .I1(\i_/badr[15]_INST_0_i_135_1 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_135_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_54 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [15]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_135_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_55 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [15]),
        .I4(\i_/badr[15]_INST_0_i_138_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [1]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_40_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [1]),
        .I4(\i_/badr[1]_INST_0_i_41_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [2]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_40_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [2]),
        .I4(\i_/badr[2]_INST_0_i_41_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [3]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_44_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [3]),
        .I4(\i_/badr[3]_INST_0_i_45_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [4]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_40_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [4]),
        .I4(\i_/badr[4]_INST_0_i_41_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [5]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_40_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [5]),
        .I4(\i_/badr[5]_INST_0_i_41_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [6]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_40_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [6]),
        .I4(\i_/badr[6]_INST_0_i_41_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_31 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [7]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_45_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [7]),
        .I4(\i_/badr[7]_INST_0_i_46_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_46 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [8]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_40_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [8]),
        .I4(\i_/badr[8]_INST_0_i_41_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_12_0 [9]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_12_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_40_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_12 [9]),
        .I4(\i_/badr[9]_INST_0_i_41_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_54_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_54_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_55_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_55_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_41_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_10
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_11 ,
    \bbus_o[4]_INST_0_i_7 ,
    \bbus_o[4]_INST_0_i_7_0 ,
    \i_/bdatw[15]_INST_0_i_36_0 ,
    \bbus_o[3]_INST_0_i_7 ,
    \bbus_o[3]_INST_0_i_7_0 ,
    \bbus_o[2]_INST_0_i_7 ,
    \bbus_o[2]_INST_0_i_7_0 ,
    \bbus_o[1]_INST_0_i_7 ,
    \bbus_o[1]_INST_0_i_7_0 ,
    \bbus_o[0]_INST_0_i_7 ,
    \bbus_o[0]_INST_0_i_7_0 ,
    \i_/bdatw[15]_INST_0_i_36_1 ,
    \i_/bdatw[15]_INST_0_i_36_2 ,
    \i_/bdatw[15]_INST_0_i_36_3 ,
    \i_/bdatw[15]_INST_0_i_36_4 ,
    \i_/bdatw[15]_INST_0_i_36_5 ,
    ctl_selb0_0,
    \i_/bdatw[15]_INST_0_i_36_6 ,
    \i_/bbus_o[4]_INST_0_i_23_0 ,
    ctl_selb0_rn,
    \bdatw[15]_INST_0_i_11_0 ,
    \bdatw[15]_INST_0_i_11_1 ,
    \bbus_o[4]_INST_0_i_7_1 ,
    \bbus_o[4]_INST_0_i_7_2 ,
    \i_/bdatw[15]_INST_0_i_35_0 ,
    \i_/bdatw[15]_INST_0_i_35_1 ,
    \bbus_o[3]_INST_0_i_7_1 ,
    \bbus_o[3]_INST_0_i_7_2 ,
    \bbus_o[2]_INST_0_i_7_1 ,
    \bbus_o[2]_INST_0_i_7_2 ,
    \bbus_o[1]_INST_0_i_7_1 ,
    \bbus_o[1]_INST_0_i_7_2 ,
    \bbus_o[0]_INST_0_i_7_1 ,
    \bbus_o[0]_INST_0_i_7_2 ,
    \i_/bdatw[15]_INST_0_i_35_2 ,
    b0bus_sel_0,
    \i_/bbus_o[5]_INST_0_i_16_0 ,
    \i_/bbus_o[4]_INST_0_i_22_0 ,
    \i_/bbus_o[4]_INST_0_i_22_1 ,
    \i_/bdatw[15]_INST_0_i_36_7 ,
    \i_/bdatw[15]_INST_0_i_98_0 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [10:0]out;
  input [15:0]\bdatw[15]_INST_0_i_11 ;
  input \bbus_o[4]_INST_0_i_7 ;
  input \bbus_o[4]_INST_0_i_7_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_36_0 ;
  input \bbus_o[3]_INST_0_i_7 ;
  input \bbus_o[3]_INST_0_i_7_0 ;
  input \bbus_o[2]_INST_0_i_7 ;
  input \bbus_o[2]_INST_0_i_7_0 ;
  input \bbus_o[1]_INST_0_i_7 ;
  input \bbus_o[1]_INST_0_i_7_0 ;
  input \bbus_o[0]_INST_0_i_7 ;
  input \bbus_o[0]_INST_0_i_7_0 ;
  input \i_/bdatw[15]_INST_0_i_36_1 ;
  input \i_/bdatw[15]_INST_0_i_36_2 ;
  input \i_/bdatw[15]_INST_0_i_36_3 ;
  input \i_/bdatw[15]_INST_0_i_36_4 ;
  input \i_/bdatw[15]_INST_0_i_36_5 ;
  input [0:0]ctl_selb0_0;
  input [10:0]\i_/bdatw[15]_INST_0_i_36_6 ;
  input \i_/bbus_o[4]_INST_0_i_23_0 ;
  input [1:0]ctl_selb0_rn;
  input [10:0]\bdatw[15]_INST_0_i_11_0 ;
  input [10:0]\bdatw[15]_INST_0_i_11_1 ;
  input \bbus_o[4]_INST_0_i_7_1 ;
  input \bbus_o[4]_INST_0_i_7_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_35_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_35_1 ;
  input \bbus_o[3]_INST_0_i_7_1 ;
  input \bbus_o[3]_INST_0_i_7_2 ;
  input \bbus_o[2]_INST_0_i_7_1 ;
  input \bbus_o[2]_INST_0_i_7_2 ;
  input \bbus_o[1]_INST_0_i_7_1 ;
  input \bbus_o[1]_INST_0_i_7_2 ;
  input \bbus_o[0]_INST_0_i_7_1 ;
  input \bbus_o[0]_INST_0_i_7_2 ;
  input \i_/bdatw[15]_INST_0_i_35_2 ;
  input [1:0]b0bus_sel_0;
  input [1:0]\i_/bbus_o[5]_INST_0_i_16_0 ;
  input \i_/bbus_o[4]_INST_0_i_22_0 ;
  input \i_/bbus_o[4]_INST_0_i_22_1 ;
  input \i_/bdatw[15]_INST_0_i_36_7 ;
  input \i_/bdatw[15]_INST_0_i_98_0 ;

  wire [1:0]b0bus_sel_0;
  wire \bbus_o[0]_INST_0_i_7 ;
  wire \bbus_o[0]_INST_0_i_7_0 ;
  wire \bbus_o[0]_INST_0_i_7_1 ;
  wire \bbus_o[0]_INST_0_i_7_2 ;
  wire \bbus_o[1]_INST_0_i_7 ;
  wire \bbus_o[1]_INST_0_i_7_0 ;
  wire \bbus_o[1]_INST_0_i_7_1 ;
  wire \bbus_o[1]_INST_0_i_7_2 ;
  wire \bbus_o[2]_INST_0_i_7 ;
  wire \bbus_o[2]_INST_0_i_7_0 ;
  wire \bbus_o[2]_INST_0_i_7_1 ;
  wire \bbus_o[2]_INST_0_i_7_2 ;
  wire \bbus_o[3]_INST_0_i_7 ;
  wire \bbus_o[3]_INST_0_i_7_0 ;
  wire \bbus_o[3]_INST_0_i_7_1 ;
  wire \bbus_o[3]_INST_0_i_7_2 ;
  wire \bbus_o[4]_INST_0_i_7 ;
  wire \bbus_o[4]_INST_0_i_7_0 ;
  wire \bbus_o[4]_INST_0_i_7_1 ;
  wire \bbus_o[4]_INST_0_i_7_2 ;
  wire [15:0]\bdatw[15]_INST_0_i_11 ;
  wire [10:0]\bdatw[15]_INST_0_i_11_0 ;
  wire [10:0]\bdatw[15]_INST_0_i_11_1 ;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bbus_o[4]_INST_0_i_22_0 ;
  wire \i_/bbus_o[4]_INST_0_i_22_1 ;
  wire \i_/bbus_o[4]_INST_0_i_23_0 ;
  wire [1:0]\i_/bbus_o[5]_INST_0_i_16_0 ;
  wire \i_/bbus_o[5]_INST_0_i_23_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_24_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_23_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_24_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_23_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_56_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_35_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_35_1 ;
  wire \i_/bdatw[15]_INST_0_i_35_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_36_0 ;
  wire \i_/bdatw[15]_INST_0_i_36_1 ;
  wire \i_/bdatw[15]_INST_0_i_36_2 ;
  wire \i_/bdatw[15]_INST_0_i_36_3 ;
  wire \i_/bdatw[15]_INST_0_i_36_4 ;
  wire \i_/bdatw[15]_INST_0_i_36_5 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_36_6 ;
  wire \i_/bdatw[15]_INST_0_i_36_7 ;
  wire \i_/bdatw[15]_INST_0_i_95_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_98_0 ;
  wire \i_/bdatw[15]_INST_0_i_98_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_50_n_0 ;
  wire [10:0]out;

  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[0]_INST_0_i_20 
       (.I0(\bbus_o[0]_INST_0_i_7_1 ),
        .I1(\bbus_o[0]_INST_0_i_7_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_35_0 [0]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_35_1 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[0]_INST_0_i_21 
       (.I0(\bbus_o[0]_INST_0_i_7 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11 [0]),
        .I3(\bbus_o[0]_INST_0_i_7_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[1]_INST_0_i_19 
       (.I0(\bbus_o[1]_INST_0_i_7_1 ),
        .I1(\bbus_o[1]_INST_0_i_7_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_35_0 [1]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_35_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[1]_INST_0_i_20 
       (.I0(\bbus_o[1]_INST_0_i_7 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11 [1]),
        .I3(\bbus_o[1]_INST_0_i_7_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[2]_INST_0_i_20 
       (.I0(\bbus_o[2]_INST_0_i_7_1 ),
        .I1(\bbus_o[2]_INST_0_i_7_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_35_0 [2]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_35_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[2]_INST_0_i_21 
       (.I0(\bbus_o[2]_INST_0_i_7 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11 [2]),
        .I3(\bbus_o[2]_INST_0_i_7_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[3]_INST_0_i_20 
       (.I0(\bbus_o[3]_INST_0_i_7_1 ),
        .I1(\bbus_o[3]_INST_0_i_7_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_35_0 [3]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_35_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[3]_INST_0_i_21 
       (.I0(\bbus_o[3]_INST_0_i_7 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11 [3]),
        .I3(\bbus_o[3]_INST_0_i_7_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[4]_INST_0_i_22 
       (.I0(\bbus_o[4]_INST_0_i_7_1 ),
        .I1(\bbus_o[4]_INST_0_i_7_2 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_35_0 [4]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_35_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[4]_INST_0_i_23 
       (.I0(\bbus_o[4]_INST_0_i_7 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11 [4]),
        .I3(\bbus_o[4]_INST_0_i_7_0 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_36_0 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bbus_o[4]_INST_0_i_22_1 ),
        .I2(\i_/bdatw[15]_INST_0_i_36_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I5(ctl_selb0_0),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bbus_o[4]_INST_0_i_22_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_36_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I5(ctl_selb0_0),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bbus_o[4]_INST_0_i_23_0 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I5(ctl_selb0_0),
        .O(gr6_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [0]),
        .I4(\i_/bbus_o[5]_INST_0_i_23_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [5]),
        .I4(\i_/bbus_o[5]_INST_0_i_24_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bbus_o[5]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [5]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [5]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bbus_o[5]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [0]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [1]),
        .I4(\i_/bbus_o[6]_INST_0_i_23_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [6]),
        .I4(\i_/bbus_o[6]_INST_0_i_24_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bbus_o[6]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [6]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [6]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bbus_o[6]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [1]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [2]),
        .I4(\i_/bbus_o[7]_INST_0_i_23_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [7]),
        .I4(\i_/bbus_o[7]_INST_0_i_24_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bbus_o[7]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [7]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [7]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bbus_o[7]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [2]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [5]),
        .I4(\i_/bdatw[10]_INST_0_i_50_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_27 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_51_n_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[10]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [10]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [10]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[10]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [6]),
        .I4(\i_/bdatw[11]_INST_0_i_50_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_51_n_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[11]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [11]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [11]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[11]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [7]),
        .I4(\i_/bdatw[12]_INST_0_i_48_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_49_n_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[12]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [12]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [12]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[12]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [8]),
        .I4(\i_/bdatw[13]_INST_0_i_50_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_51_n_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[13]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [13]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [13]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[13]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [9]),
        .I4(\i_/bdatw[14]_INST_0_i_55_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_27 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_56_n_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[14]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [14]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [14]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[14]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_176 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_98_0 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I5(ctl_selb0_0),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [10]),
        .I4(\i_/bdatw[15]_INST_0_i_95_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_98_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_93 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_36_7 ),
        .I2(\i_/bdatw[15]_INST_0_i_36_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I5(ctl_selb0_0),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_94 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_35_2 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I5(ctl_selb0_0),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[15]_INST_0_i_95 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [15]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [15]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[15]_INST_0_i_95_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/bdatw[15]_INST_0_i_96 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_36_7 ),
        .I2(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I3(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I4(ctl_selb0_0),
        .I5(\i_/bdatw[15]_INST_0_i_36_3 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_97 
       (.I0(\i_/bdatw[15]_INST_0_i_36_1 ),
        .I1(\i_/bdatw[15]_INST_0_i_36_2 ),
        .I2(\i_/bdatw[15]_INST_0_i_36_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_36_4 ),
        .I4(\i_/bdatw[15]_INST_0_i_36_5 ),
        .I5(ctl_selb0_0),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_98 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_98_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [3]),
        .I4(\i_/bdatw[8]_INST_0_i_49_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_50_n_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[8]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [8]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [8]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[8]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [4]),
        .I4(\i_/bdatw[9]_INST_0_i_49_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_26 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_50_n_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hF800000088000000)) 
    \i_/bdatw[9]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_35_1 [9]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_35_0 [9]),
        .I3(\i_/bbus_o[5]_INST_0_i_16_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_16_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[9]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_36_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_36_6 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_50_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_11
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_15 ,
    \i_/bdatw[15]_INST_0_i_48_0 ,
    \i_/bdatw[15]_INST_0_i_48_1 ,
    \i_/bdatw[15]_INST_0_i_212_0 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_212_1 ,
    \i_/bdatw[15]_INST_0_i_124_0 ,
    \i_/bdatw[15]_INST_0_i_48_2 ,
    \i_/bdatw[15]_INST_0_i_48_3 ,
    \i_/bdatw[8]_INST_0_i_69_0 ,
    \i_/bdatw[15]_INST_0_i_121_0 ,
    \i_/bdatw[15]_INST_0_i_121_1 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_121_2 ,
    \i_/bdatw[15]_INST_0_i_124_1 ,
    \i_/bdatw[15]_INST_0_i_124_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_15 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_1 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_212_0 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_212_1 ;
  input \i_/bdatw[15]_INST_0_i_124_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_3 ;
  input \i_/bdatw[8]_INST_0_i_69_0 ;
  input \i_/bdatw[15]_INST_0_i_121_0 ;
  input \i_/bdatw[15]_INST_0_i_121_1 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_121_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_124_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_124_2 ;

  wire [15:0]\bdatw[15]_INST_0_i_15 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[10]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_76_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_76_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_74_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_72_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_101_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_102_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_72_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_121_0 ;
  wire \i_/bdatw[15]_INST_0_i_121_1 ;
  wire \i_/bdatw[15]_INST_0_i_121_2 ;
  wire \i_/bdatw[15]_INST_0_i_121_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_124_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_124_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_124_2 ;
  wire \i_/bdatw[15]_INST_0_i_124_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_212_0 ;
  wire \i_/bdatw[15]_INST_0_i_212_1 ;
  wire \i_/bdatw[15]_INST_0_i_212_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_218_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_219_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_3 ;
  wire \i_/bdatw[8]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_69_0 ;
  wire \i_/bdatw[8]_INST_0_i_75_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_75_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_54_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [10]),
        .I2(gr0_bus1),
        .I3(out[10]),
        .I4(\i_/bdatw[10]_INST_0_i_55_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_68 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_15 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_69 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [2]),
        .I4(\i_/bdatw[10]_INST_0_i_76_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[10]_INST_0_i_76 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_124_2 [2]),
        .I2(\i_/bdatw[8]_INST_0_i_69_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(\i_/bdatw[10]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_54_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [11]),
        .I2(gr0_bus1),
        .I3(out[11]),
        .I4(\i_/bdatw[11]_INST_0_i_55_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_68 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_69 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_15 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_70 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [3]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [3]),
        .I4(\i_/bdatw[11]_INST_0_i_76_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[11]_INST_0_i_76 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_124_2 [3]),
        .I2(\i_/bdatw[8]_INST_0_i_69_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(\i_/bdatw[11]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_52_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [12]),
        .I2(gr0_bus1),
        .I3(out[12]),
        .I4(\i_/bdatw[12]_INST_0_i_53_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_67 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_15 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_68 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [4]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [4]),
        .I4(\i_/bdatw[12]_INST_0_i_74_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[12]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_124_2 [4]),
        .I2(\i_/bdatw[8]_INST_0_i_69_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(\i_/bdatw[12]_INST_0_i_74_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_54_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [13]),
        .I2(gr0_bus1),
        .I3(out[13]),
        .I4(\i_/bdatw[13]_INST_0_i_55_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_55_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_64 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_71_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_65 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[13]_INST_0_i_72_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_71_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_72 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_72_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_101 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_101_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_102 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_102_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_40 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_71_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_41 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [14]),
        .I2(gr0_bus1),
        .I3(out[14]),
        .I4(\i_/bdatw[14]_INST_0_i_72_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \i_/bdatw[14]_INST_0_i_69 
       (.I0(\i_/bdatw[15]_INST_0_i_212_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_212_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/bdatw[14]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_212_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_212_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_124_0 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_71_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_72 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_72_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_83 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_101_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_84 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [6]),
        .I2(gr0_bus1),
        .I3(out[6]),
        .I4(\i_/bdatw[14]_INST_0_i_102_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[14]_INST_0_i_95 
       (.I0(\i_/bdatw[15]_INST_0_i_212_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_212_0 [0]),
        .I2(ctl_selb1_rn[0]),
        .I3(ctl_selb1_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[14]_INST_0_i_96 
       (.I0(\i_/bdatw[15]_INST_0_i_212_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_212_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_121 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_121_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \i_/bdatw[15]_INST_0_i_122 
       (.I0(\i_/bdatw[15]_INST_0_i_212_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_212_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/bdatw[15]_INST_0_i_123 
       (.I0(\i_/bdatw[15]_INST_0_i_212_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_212_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_124_0 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_124 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_212_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_124_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_135 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_218_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_136 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [7]),
        .I2(gr0_bus1),
        .I3(out[7]),
        .I4(\i_/bdatw[15]_INST_0_i_219_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/bdatw[15]_INST_0_i_210 
       (.I0(\i_/bdatw[15]_INST_0_i_212_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_212_0 [0]),
        .I2(ctl_selb1_rn[2]),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_124_0 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_211 
       (.I0(\i_/bdatw[8]_INST_0_i_69_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_121_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_121_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_121_2 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_212 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_212_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_218 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_218_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_219 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_121_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_15 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_124_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_53_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [8]),
        .I2(gr0_bus1),
        .I3(out[8]),
        .I4(\i_/bdatw[8]_INST_0_i_54_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_68 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_15 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_69 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [0]),
        .I4(\i_/bdatw[8]_INST_0_i_75_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[8]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_124_2 [0]),
        .I2(\i_/bdatw[8]_INST_0_i_69_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(\i_/bdatw[8]_INST_0_i_75_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_53_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [9]),
        .I2(gr0_bus1),
        .I3(out[9]),
        .I4(\i_/bdatw[9]_INST_0_i_54_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_124_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_48_2 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_3 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_67 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_15 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_68 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_48_1 [1]),
        .I4(\i_/bdatw[9]_INST_0_i_75_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[9]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_124_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_124_2 [1]),
        .I2(\i_/bdatw[8]_INST_0_i_69_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_212_1 ),
        .O(\i_/bdatw[9]_INST_0_i_75_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_12
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_15 ,
    \bdatw[12]_INST_0_i_42 ,
    \i_/bdatw[15]_INST_0_i_49_0 ,
    \bdatw[12]_INST_0_i_42_0 ,
    \bdatw[11]_INST_0_i_44 ,
    \bdatw[11]_INST_0_i_44_0 ,
    \bdatw[10]_INST_0_i_43 ,
    \bdatw[10]_INST_0_i_43_0 ,
    \bdatw[9]_INST_0_i_42 ,
    \bdatw[9]_INST_0_i_42_0 ,
    \bdatw[8]_INST_0_i_43 ,
    \bdatw[8]_INST_0_i_43_0 ,
    \i_/bdatw[15]_INST_0_i_49_1 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_128_0 ,
    \i_/bdatw[15]_INST_0_i_49_2 ,
    \i_/bdatw[15]_INST_0_i_49_3 ,
    \i_/bdatw[15]_INST_0_i_49_4 ,
    \i_/bdatw[15]_INST_0_i_49_5 ,
    \i_/bdatw[15]_INST_0_i_128_1 ,
    \i_/bdatw[15]_INST_0_i_128_2 ,
    \i_/bdatw[12]_INST_0_i_64_0 ,
    \i_/bdatw[12]_INST_0_i_64_1 ,
    \i_/bdatw[12]_INST_0_i_64_2 ,
    ctl_selb1_0,
    \i_/bdatw[12]_INST_0_i_64_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [10:0]out;
  input [15:0]\bdatw[15]_INST_0_i_15 ;
  input \bdatw[12]_INST_0_i_42 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_49_0 ;
  input \bdatw[12]_INST_0_i_42_0 ;
  input \bdatw[11]_INST_0_i_44 ;
  input \bdatw[11]_INST_0_i_44_0 ;
  input \bdatw[10]_INST_0_i_43 ;
  input \bdatw[10]_INST_0_i_43_0 ;
  input \bdatw[9]_INST_0_i_42 ;
  input \bdatw[9]_INST_0_i_42_0 ;
  input \bdatw[8]_INST_0_i_43 ;
  input \bdatw[8]_INST_0_i_43_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_49_1 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_128_0 ;
  input [10:0]\i_/bdatw[15]_INST_0_i_49_2 ;
  input \i_/bdatw[15]_INST_0_i_49_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_49_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_49_5 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_128_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_128_2 ;
  input \i_/bdatw[12]_INST_0_i_64_0 ;
  input \i_/bdatw[12]_INST_0_i_64_1 ;
  input \i_/bdatw[12]_INST_0_i_64_2 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[12]_INST_0_i_64_3 ;

  wire \bdatw[10]_INST_0_i_43 ;
  wire \bdatw[10]_INST_0_i_43_0 ;
  wire \bdatw[11]_INST_0_i_44 ;
  wire \bdatw[11]_INST_0_i_44_0 ;
  wire \bdatw[12]_INST_0_i_42 ;
  wire \bdatw[12]_INST_0_i_42_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_15 ;
  wire \bdatw[8]_INST_0_i_43 ;
  wire \bdatw[8]_INST_0_i_43_0 ;
  wire \bdatw[9]_INST_0_i_42 ;
  wire \bdatw[9]_INST_0_i_42_0 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bdatw[10]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_75_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_75_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_64_0 ;
  wire \i_/bdatw[12]_INST_0_i_64_1 ;
  wire \i_/bdatw[12]_INST_0_i_64_2 ;
  wire \i_/bdatw[12]_INST_0_i_64_3 ;
  wire \i_/bdatw[12]_INST_0_i_73_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_57_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_73_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_74_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_103_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_104_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_75_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_76_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_125_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_128_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_128_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_128_2 ;
  wire \i_/bdatw[15]_INST_0_i_128_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_215_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_220_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_221_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_49_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_49_1 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_49_2 ;
  wire \i_/bdatw[15]_INST_0_i_49_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_49_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_49_5 ;
  wire \i_/bdatw[8]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_74_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_74_n_0 ;
  wire [10:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_56_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [10]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[10]_INST_0_i_57_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bdatw[10]_INST_0_i_65 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [2]),
        .I2(\bdatw[10]_INST_0_i_43 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_0 [2]),
        .I5(\bdatw[10]_INST_0_i_43_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_66 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [2]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [2]),
        .I4(\i_/bdatw[10]_INST_0_i_75_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[10]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_128_2 [2]),
        .I2(\i_/bdatw[12]_INST_0_i_64_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(\i_/bdatw[10]_INST_0_i_75_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_56_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [11]),
        .I2(gr0_bus1),
        .I3(out[6]),
        .I4(\i_/bdatw[11]_INST_0_i_57_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bdatw[11]_INST_0_i_66 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [3]),
        .I2(\bdatw[11]_INST_0_i_44 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_0 [3]),
        .I5(\bdatw[11]_INST_0_i_44_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_67 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [3]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [3]),
        .I4(\i_/bdatw[11]_INST_0_i_75_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[11]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_128_2 [3]),
        .I2(\i_/bdatw[12]_INST_0_i_64_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(\i_/bdatw[11]_INST_0_i_75_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_35 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_54_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [12]),
        .I2(gr0_bus1),
        .I3(out[7]),
        .I4(\i_/bdatw[12]_INST_0_i_55_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bdatw[12]_INST_0_i_64 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [4]),
        .I2(\bdatw[12]_INST_0_i_42 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_0 [4]),
        .I5(\bdatw[12]_INST_0_i_42_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_65 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [4]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [4]),
        .I4(\i_/bdatw[12]_INST_0_i_73_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[12]_INST_0_i_73 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_128_2 [4]),
        .I2(\i_/bdatw[12]_INST_0_i_64_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(\i_/bdatw[12]_INST_0_i_73_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_37 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_56_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [13]),
        .I2(gr0_bus1),
        .I3(out[8]),
        .I4(\i_/bdatw[13]_INST_0_i_57_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_66 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_73_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_67 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [5]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/bdatw[13]_INST_0_i_74_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_73 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_73_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_74_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_103 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_103_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_104 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_104_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_42 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_75_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_43 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [14]),
        .I2(gr0_bus1),
        .I3(out[9]),
        .I4(\i_/bdatw[14]_INST_0_i_76_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \i_/bdatw[14]_INST_0_i_73 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \i_/bdatw[14]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_49_3 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_75 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_75_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_76 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_85 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_103_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_86 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [6]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[14]_INST_0_i_104_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[14]_INST_0_i_97 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I2(ctl_selb1_rn[0]),
        .I3(ctl_selb1_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000800)) 
    \i_/bdatw[14]_INST_0_i_98 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_125 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_125_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \i_/bdatw[15]_INST_0_i_126 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \i_/bdatw[15]_INST_0_i_127 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_49_3 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_128 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_215_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_128_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_137 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_220_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_138 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [7]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[15]_INST_0_i_221_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \i_/bdatw[15]_INST_0_i_213 
       (.I0(\i_/bdatw[15]_INST_0_i_49_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_49_1 [0]),
        .I2(ctl_selb1_rn[2]),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_49_3 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[15]_INST_0_i_214 
       (.I0(\i_/bdatw[12]_INST_0_i_64_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_64_1 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[12]_INST_0_i_64_2 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[12]_INST_0_i_64_3 ),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_215 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_215_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_220 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_220_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_221 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_221_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_125_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_15 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_128_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_55_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [8]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[8]_INST_0_i_56_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bdatw[8]_INST_0_i_65 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [0]),
        .I2(\bdatw[8]_INST_0_i_43 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_0 [0]),
        .I5(\bdatw[8]_INST_0_i_43_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_66 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [0]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [0]),
        .I4(\i_/bdatw[8]_INST_0_i_74_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[8]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_128_2 [0]),
        .I2(\i_/bdatw[12]_INST_0_i_64_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(\i_/bdatw[8]_INST_0_i_74_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_36 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_55_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [9]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[9]_INST_0_i_56_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_128_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_49_2 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_49_0 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \i_/bdatw[9]_INST_0_i_64 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_15 [1]),
        .I2(\bdatw[9]_INST_0_i_42 ),
        .I3(gr5_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_49_0 [1]),
        .I5(\bdatw[9]_INST_0_i_42_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_65 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_49_4 [1]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_49_5 [1]),
        .I4(\i_/bdatw[9]_INST_0_i_74_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[9]_INST_0_i_74 
       (.I0(\i_/bdatw[15]_INST_0_i_128_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_128_2 [1]),
        .I2(\i_/bdatw[12]_INST_0_i_64_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_128_0 ),
        .O(\i_/bdatw[9]_INST_0_i_74_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_28
   (p_1_in,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[14] ,
    \grn_reg[14]_0 ,
    \grn_reg[13] ,
    \grn_reg[13]_0 ,
    \grn_reg[12] ,
    \grn_reg[12]_0 ,
    \grn_reg[11] ,
    \grn_reg[11]_0 ,
    \grn_reg[10] ,
    \grn_reg[10]_0 ,
    \grn_reg[9] ,
    \grn_reg[9]_0 ,
    \grn_reg[8] ,
    \grn_reg[8]_0 ,
    \grn_reg[7] ,
    \grn_reg[7]_0 ,
    \grn_reg[6] ,
    \grn_reg[6]_0 ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[3] ,
    \grn_reg[3]_0 ,
    \grn_reg[2] ,
    \grn_reg[2]_0 ,
    \grn_reg[1] ,
    \grn_reg[1]_0 ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[0]_1 ,
    out,
    \rgf_c0bus_wb[4]_i_41 ,
    \i_/badr[15]_INST_0_i_10_0 ,
    a0bus_sel_0,
    \i_/badr[15]_INST_0_i_10_1 ,
    \i_/badr[15]_INST_0_i_10_2 ,
    bank_sel,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_43_0 ,
    ctl_sela0,
    \i_/badr[15]_INST_0_i_43_1 ,
    \rgf_c0bus_wb[4]_i_41_0 ,
    \rgf_c0bus_wb[4]_i_41_1 ,
    \i_/badr[15]_INST_0_i_46_0 ,
    \i_/badr[15]_INST_0_i_46_1 );
  output [14:0]p_1_in;
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14] ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13] ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12] ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11] ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10] ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9] ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8] ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7] ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6] ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3] ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2] ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1] ;
  output \grn_reg[1]_0 ;
  output [0:0]\grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\rgf_c0bus_wb[4]_i_41 ;
  input [1:0]\i_/badr[15]_INST_0_i_10_0 ;
  input [3:0]a0bus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_10_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_10_2 ;
  input [0:0]bank_sel;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_43_0 ;
  input [0:0]ctl_sela0;
  input \i_/badr[15]_INST_0_i_43_1 ;
  input [15:0]\rgf_c0bus_wb[4]_i_41_0 ;
  input [15:0]\rgf_c0bus_wb[4]_i_41_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_46_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_46_1 ;

  wire [3:0]a0bus_sel_0;
  wire [0:0]bank_sel;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [0:0]\grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_25_n_0 ;
  wire \i_/badr[0]_INST_0_i_38_n_0 ;
  wire \i_/badr[10]_INST_0_i_24_n_0 ;
  wire \i_/badr[10]_INST_0_i_36_n_0 ;
  wire \i_/badr[11]_INST_0_i_25_n_0 ;
  wire \i_/badr[11]_INST_0_i_41_n_0 ;
  wire \i_/badr[12]_INST_0_i_24_n_0 ;
  wire \i_/badr[12]_INST_0_i_36_n_0 ;
  wire \i_/badr[13]_INST_0_i_24_n_0 ;
  wire \i_/badr[13]_INST_0_i_36_n_0 ;
  wire \i_/badr[14]_INST_0_i_24_n_0 ;
  wire \i_/badr[14]_INST_0_i_36_n_0 ;
  wire [1:0]\i_/badr[15]_INST_0_i_10_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_10_2 ;
  wire \i_/badr[15]_INST_0_i_121_n_0 ;
  wire \i_/badr[15]_INST_0_i_43_0 ;
  wire \i_/badr[15]_INST_0_i_43_1 ;
  wire \i_/badr[15]_INST_0_i_43_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_46_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_46_1 ;
  wire \i_/badr[1]_INST_0_i_24_n_0 ;
  wire \i_/badr[1]_INST_0_i_36_n_0 ;
  wire \i_/badr[2]_INST_0_i_24_n_0 ;
  wire \i_/badr[2]_INST_0_i_36_n_0 ;
  wire \i_/badr[3]_INST_0_i_25_n_0 ;
  wire \i_/badr[3]_INST_0_i_40_n_0 ;
  wire \i_/badr[4]_INST_0_i_24_n_0 ;
  wire \i_/badr[4]_INST_0_i_36_n_0 ;
  wire \i_/badr[5]_INST_0_i_24_n_0 ;
  wire \i_/badr[5]_INST_0_i_36_n_0 ;
  wire \i_/badr[6]_INST_0_i_24_n_0 ;
  wire \i_/badr[6]_INST_0_i_36_n_0 ;
  wire \i_/badr[7]_INST_0_i_25_n_0 ;
  wire \i_/badr[7]_INST_0_i_41_n_0 ;
  wire \i_/badr[8]_INST_0_i_24_n_0 ;
  wire \i_/badr[8]_INST_0_i_36_n_0 ;
  wire \i_/badr[9]_INST_0_i_24_n_0 ;
  wire \i_/badr[9]_INST_0_i_36_n_0 ;
  wire [15:0]out;
  wire [14:0]p_1_in;
  wire [15:0]\rgf_c0bus_wb[4]_i_41 ;
  wire [15:0]\rgf_c0bus_wb[4]_i_41_0 ;
  wire [15:0]\rgf_c0bus_wb[4]_i_41_1 ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[0]_INST_0_i_10 
       (.I0(\i_/badr[0]_INST_0_i_25_n_0 ),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [0]),
        .I4(gr7_bus1),
        .I5(\grn_reg[0]_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_38_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_38 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[10]_INST_0_i_10 
       (.I0(\i_/badr[10]_INST_0_i_24_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [10]),
        .I4(gr7_bus1),
        .I5(\grn_reg[10] ),
        .O(p_1_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_36_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[11]_INST_0_i_10 
       (.I0(\i_/badr[11]_INST_0_i_25_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [11]),
        .I4(gr7_bus1),
        .I5(\grn_reg[11] ),
        .O(p_1_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_41_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[12]_INST_0_i_10 
       (.I0(\i_/badr[12]_INST_0_i_24_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [12]),
        .I4(gr7_bus1),
        .I5(\grn_reg[12] ),
        .O(p_1_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_36_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[13]_INST_0_i_10 
       (.I0(\i_/badr[13]_INST_0_i_24_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [13]),
        .I4(gr7_bus1),
        .I5(\grn_reg[13] ),
        .O(p_1_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_36_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[14]_INST_0_i_10 
       (.I0(\i_/badr[14]_INST_0_i_24_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [14]),
        .I4(gr7_bus1),
        .I5(\grn_reg[14] ),
        .O(p_1_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_36_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[15]_INST_0_i_10 
       (.I0(\i_/badr[15]_INST_0_i_43_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [15]),
        .I4(gr7_bus1),
        .I5(\grn_reg[15] ),
        .O(p_1_in[14]));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_115 
       (.I0(bank_sel),
        .I1(ctl_sela0_rn[1]),
        .I2(\i_/badr[15]_INST_0_i_43_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_43_1 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_116 
       (.I0(bank_sel),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\i_/badr[15]_INST_0_i_43_0 ),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_43_1 ),
        .O(gr5_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_119 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I2(a0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_120 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I2(a0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_121 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_121_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_212 
       (.I0(bank_sel),
        .I1(ctl_sela0_rn[0]),
        .I2(\i_/badr[15]_INST_0_i_43_0 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_43_1 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_213 
       (.I0(bank_sel),
        .I1(\i_/badr[15]_INST_0_i_43_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_43_1 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_44 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I2(a0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_45 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I2(a0bus_sel_0[3]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_46 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_121_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[1]_INST_0_i_10 
       (.I0(\i_/badr[1]_INST_0_i_24_n_0 ),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [1]),
        .I4(gr7_bus1),
        .I5(\grn_reg[1] ),
        .O(p_1_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_36_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[2]_INST_0_i_10 
       (.I0(\i_/badr[2]_INST_0_i_24_n_0 ),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [2]),
        .I4(gr7_bus1),
        .I5(\grn_reg[2] ),
        .O(p_1_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_36_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[3]_INST_0_i_10 
       (.I0(\i_/badr[3]_INST_0_i_25_n_0 ),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [3]),
        .I4(gr7_bus1),
        .I5(\grn_reg[3] ),
        .O(p_1_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_40_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[4]_INST_0_i_10 
       (.I0(\i_/badr[4]_INST_0_i_24_n_0 ),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [4]),
        .I4(gr7_bus1),
        .I5(\grn_reg[4] ),
        .O(p_1_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_36_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[5]_INST_0_i_10 
       (.I0(\i_/badr[5]_INST_0_i_24_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [5]),
        .I4(gr7_bus1),
        .I5(\grn_reg[5] ),
        .O(p_1_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_36_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[6]_INST_0_i_10 
       (.I0(\i_/badr[6]_INST_0_i_24_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [6]),
        .I4(gr7_bus1),
        .I5(\grn_reg[6] ),
        .O(p_1_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_36_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[7]_INST_0_i_10 
       (.I0(\i_/badr[7]_INST_0_i_25_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [7]),
        .I4(gr7_bus1),
        .I5(\grn_reg[7] ),
        .O(p_1_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_26 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_41_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[8]_INST_0_i_10 
       (.I0(\i_/badr[8]_INST_0_i_24_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [8]),
        .I4(gr7_bus1),
        .I5(\grn_reg[8] ),
        .O(p_1_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_36_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[9]_INST_0_i_10 
       (.I0(\i_/badr[9]_INST_0_i_24_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [9]),
        .I4(gr7_bus1),
        .I5(\grn_reg[9] ),
        .O(p_1_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_10_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_25 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_36_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_46_0 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_46_1 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_100 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [8]),
        .I2(gr0_bus1),
        .I3(out[8]),
        .I4(\i_/badr[8]_INST_0_i_24_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_105 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/badr[5]_INST_0_i_24_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_65 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [2]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/badr[2]_INST_0_i_24_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_68 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [1]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/badr[1]_INST_0_i_24_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_70 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [4]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/badr[4]_INST_0_i_24_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_73 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [3]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/badr[3]_INST_0_i_25_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_75 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [15]),
        .I2(gr0_bus1),
        .I3(out[15]),
        .I4(\i_/badr[15]_INST_0_i_43_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_77 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [14]),
        .I2(gr0_bus1),
        .I3(out[14]),
        .I4(\i_/badr[14]_INST_0_i_24_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_80 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [0]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/badr[0]_INST_0_i_25_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_82 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [11]),
        .I2(gr0_bus1),
        .I3(out[11]),
        .I4(\i_/badr[11]_INST_0_i_25_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_85 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [10]),
        .I2(gr0_bus1),
        .I3(out[10]),
        .I4(\i_/badr[10]_INST_0_i_24_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_87 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [13]),
        .I2(gr0_bus1),
        .I3(out[13]),
        .I4(\i_/badr[13]_INST_0_i_24_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_90 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [12]),
        .I2(gr0_bus1),
        .I3(out[12]),
        .I4(\i_/badr[12]_INST_0_i_24_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_92 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [7]),
        .I2(gr0_bus1),
        .I3(out[7]),
        .I4(\i_/badr[7]_INST_0_i_25_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_95 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [6]),
        .I2(gr0_bus1),
        .I3(out[6]),
        .I4(\i_/badr[6]_INST_0_i_24_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_97 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [9]),
        .I2(gr0_bus1),
        .I3(out[9]),
        .I4(\i_/badr[9]_INST_0_i_24_n_0 ),
        .O(\grn_reg[9]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_29
   (p_0_in,
    \grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_1 ,
    out,
    \rgf_c0bus_wb[4]_i_41 ,
    \rgf_c0bus_wb[4]_i_41_0 ,
    \rgf_c0bus_wb[4]_i_41_1 ,
    \i_/badr[15]_INST_0_i_50_0 ,
    a0bus_sel_0,
    \i_/badr[15]_INST_0_i_11_0 ,
    \i_/badr[15]_INST_0_i_11_1 ,
    \i_/badr[15]_INST_0_i_47_0 ,
    ctl_sela0_rn,
    \i_/badr[15]_INST_0_i_47_1 ,
    ctl_sela0,
    \i_/badr[15]_INST_0_i_47_2 ,
    \i_/badr[15]_INST_0_i_50_1 ,
    \i_/badr[15]_INST_0_i_50_2 );
  output [14:0]p_0_in;
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output [0:0]\grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\rgf_c0bus_wb[4]_i_41 ;
  input [15:0]\rgf_c0bus_wb[4]_i_41_0 ;
  input [15:0]\rgf_c0bus_wb[4]_i_41_1 ;
  input [1:0]\i_/badr[15]_INST_0_i_50_0 ;
  input [3:0]a0bus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_11_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_1 ;
  input \i_/badr[15]_INST_0_i_47_0 ;
  input [1:0]ctl_sela0_rn;
  input \i_/badr[15]_INST_0_i_47_1 ;
  input [0:0]ctl_sela0;
  input \i_/badr[15]_INST_0_i_47_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_50_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_50_2 ;

  wire [3:0]a0bus_sel_0;
  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [0:0]\grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_27_n_0 ;
  wire \i_/badr[0]_INST_0_i_39_n_0 ;
  wire \i_/badr[10]_INST_0_i_26_n_0 ;
  wire \i_/badr[10]_INST_0_i_37_n_0 ;
  wire \i_/badr[11]_INST_0_i_27_n_0 ;
  wire \i_/badr[11]_INST_0_i_42_n_0 ;
  wire \i_/badr[12]_INST_0_i_26_n_0 ;
  wire \i_/badr[12]_INST_0_i_37_n_0 ;
  wire \i_/badr[13]_INST_0_i_26_n_0 ;
  wire \i_/badr[13]_INST_0_i_37_n_0 ;
  wire \i_/badr[14]_INST_0_i_26_n_0 ;
  wire \i_/badr[14]_INST_0_i_37_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_1 ;
  wire \i_/badr[15]_INST_0_i_126_n_0 ;
  wire \i_/badr[15]_INST_0_i_47_0 ;
  wire \i_/badr[15]_INST_0_i_47_1 ;
  wire \i_/badr[15]_INST_0_i_47_2 ;
  wire \i_/badr[15]_INST_0_i_47_n_0 ;
  wire [1:0]\i_/badr[15]_INST_0_i_50_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_50_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_50_2 ;
  wire \i_/badr[1]_INST_0_i_26_n_0 ;
  wire \i_/badr[1]_INST_0_i_37_n_0 ;
  wire \i_/badr[2]_INST_0_i_26_n_0 ;
  wire \i_/badr[2]_INST_0_i_37_n_0 ;
  wire \i_/badr[3]_INST_0_i_27_n_0 ;
  wire \i_/badr[3]_INST_0_i_41_n_0 ;
  wire \i_/badr[4]_INST_0_i_26_n_0 ;
  wire \i_/badr[4]_INST_0_i_37_n_0 ;
  wire \i_/badr[5]_INST_0_i_26_n_0 ;
  wire \i_/badr[5]_INST_0_i_37_n_0 ;
  wire \i_/badr[6]_INST_0_i_26_n_0 ;
  wire \i_/badr[6]_INST_0_i_37_n_0 ;
  wire \i_/badr[7]_INST_0_i_27_n_0 ;
  wire \i_/badr[7]_INST_0_i_42_n_0 ;
  wire \i_/badr[8]_INST_0_i_26_n_0 ;
  wire \i_/badr[8]_INST_0_i_37_n_0 ;
  wire \i_/badr[9]_INST_0_i_26_n_0 ;
  wire \i_/badr[9]_INST_0_i_37_n_0 ;
  wire [15:0]out;
  wire [14:0]p_0_in;
  wire [15:0]\rgf_c0bus_wb[4]_i_41 ;
  wire [15:0]\rgf_c0bus_wb[4]_i_41_0 ;
  wire [15:0]\rgf_c0bus_wb[4]_i_41_1 ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[0]_INST_0_i_11 
       (.I0(\i_/badr[0]_INST_0_i_27_n_0 ),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [0]),
        .I4(gr7_bus1),
        .I5(\grn_reg[0]_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_39_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [0]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[10]_INST_0_i_11 
       (.I0(\i_/badr[10]_INST_0_i_26_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [10]),
        .I4(gr7_bus1),
        .I5(\grn_reg[10] ),
        .O(p_0_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_37_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[11]_INST_0_i_11 
       (.I0(\i_/badr[11]_INST_0_i_27_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [11]),
        .I4(gr7_bus1),
        .I5(\grn_reg[11] ),
        .O(p_0_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_42_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[12]_INST_0_i_11 
       (.I0(\i_/badr[12]_INST_0_i_26_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [12]),
        .I4(gr7_bus1),
        .I5(\grn_reg[12] ),
        .O(p_0_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_37_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[13]_INST_0_i_11 
       (.I0(\i_/badr[13]_INST_0_i_26_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [13]),
        .I4(gr7_bus1),
        .I5(\grn_reg[13] ),
        .O(p_0_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_37_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[14]_INST_0_i_11 
       (.I0(\i_/badr[14]_INST_0_i_26_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [14]),
        .I4(gr7_bus1),
        .I5(\grn_reg[14] ),
        .O(p_0_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_37_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[15]_INST_0_i_11 
       (.I0(\i_/badr[15]_INST_0_i_47_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [15]),
        .I4(gr7_bus1),
        .I5(\grn_reg[15] ),
        .O(p_0_in[14]));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_122 
       (.I0(\i_/badr[15]_INST_0_i_47_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\i_/badr[15]_INST_0_i_47_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_47_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_123 
       (.I0(\i_/badr[15]_INST_0_i_47_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\i_/badr[15]_INST_0_i_47_1 ),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_47_2 ),
        .O(gr5_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_124 
       (.I0(\i_/badr[15]_INST_0_i_50_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_50_0 [1]),
        .I2(a0bus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_125 
       (.I0(\i_/badr[15]_INST_0_i_50_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_50_0 [1]),
        .I2(a0bus_sel_0[2]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_126 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_126_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_214 
       (.I0(\i_/badr[15]_INST_0_i_47_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\i_/badr[15]_INST_0_i_47_1 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_47_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_215 
       (.I0(\i_/badr[15]_INST_0_i_47_0 ),
        .I1(\i_/badr[15]_INST_0_i_47_1 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_47_2 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_47 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_48 
       (.I0(\i_/badr[15]_INST_0_i_50_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_50_0 [1]),
        .I2(a0bus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_49 
       (.I0(\i_/badr[15]_INST_0_i_50_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_50_0 [1]),
        .I2(a0bus_sel_0[3]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_50 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_126_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[1]_INST_0_i_11 
       (.I0(\i_/badr[1]_INST_0_i_26_n_0 ),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [1]),
        .I4(gr7_bus1),
        .I5(\grn_reg[1] ),
        .O(p_0_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [1]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_37_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [1]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[2]_INST_0_i_11 
       (.I0(\i_/badr[2]_INST_0_i_26_n_0 ),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [2]),
        .I4(gr7_bus1),
        .I5(\grn_reg[2] ),
        .O(p_0_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [2]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_37_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [2]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[3]_INST_0_i_11 
       (.I0(\i_/badr[3]_INST_0_i_27_n_0 ),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [3]),
        .I4(gr7_bus1),
        .I5(\grn_reg[3] ),
        .O(p_0_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [3]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_41_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [3]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[4]_INST_0_i_11 
       (.I0(\i_/badr[4]_INST_0_i_26_n_0 ),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [4]),
        .I4(gr7_bus1),
        .I5(\grn_reg[4] ),
        .O(p_0_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [4]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_37_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [4]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[5]_INST_0_i_11 
       (.I0(\i_/badr[5]_INST_0_i_26_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [5]),
        .I4(gr7_bus1),
        .I5(\grn_reg[5] ),
        .O(p_0_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [5]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_37_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[6]_INST_0_i_11 
       (.I0(\i_/badr[6]_INST_0_i_26_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [6]),
        .I4(gr7_bus1),
        .I5(\grn_reg[6] ),
        .O(p_0_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_37_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[7]_INST_0_i_11 
       (.I0(\i_/badr[7]_INST_0_i_27_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [7]),
        .I4(gr7_bus1),
        .I5(\grn_reg[7] ),
        .O(p_0_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_28 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_42_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[8]_INST_0_i_11 
       (.I0(\i_/badr[8]_INST_0_i_26_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [8]),
        .I4(gr7_bus1),
        .I5(\grn_reg[8] ),
        .O(p_0_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_37_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[9]_INST_0_i_11 
       (.I0(\i_/badr[9]_INST_0_i_26_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41 [9]),
        .I4(gr7_bus1),
        .I5(\grn_reg[9] ),
        .O(p_0_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/badr[15]_INST_0_i_11_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_27 
       (.I0(gr3_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41_0 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c0bus_wb[4]_i_41_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_37_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_50_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/badr[15]_INST_0_i_50_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_104 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/badr[5]_INST_0_i_26_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_64 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [2]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/badr[2]_INST_0_i_26_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_67 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [1]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/badr[1]_INST_0_i_26_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_69 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [4]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/badr[4]_INST_0_i_26_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_72 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [3]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/badr[3]_INST_0_i_27_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_74 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [15]),
        .I2(gr0_bus1),
        .I3(out[15]),
        .I4(\i_/badr[15]_INST_0_i_47_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_76 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [14]),
        .I2(gr0_bus1),
        .I3(out[14]),
        .I4(\i_/badr[14]_INST_0_i_26_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_79 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [0]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/badr[0]_INST_0_i_27_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_81 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [11]),
        .I2(gr0_bus1),
        .I3(out[11]),
        .I4(\i_/badr[11]_INST_0_i_27_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_84 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [10]),
        .I2(gr0_bus1),
        .I3(out[10]),
        .I4(\i_/badr[10]_INST_0_i_26_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_86 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [13]),
        .I2(gr0_bus1),
        .I3(out[13]),
        .I4(\i_/badr[13]_INST_0_i_26_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_89 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [12]),
        .I2(gr0_bus1),
        .I3(out[12]),
        .I4(\i_/badr[12]_INST_0_i_26_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_91 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [7]),
        .I2(gr0_bus1),
        .I3(out[7]),
        .I4(\i_/badr[7]_INST_0_i_27_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_94 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [6]),
        .I2(gr0_bus1),
        .I3(out[6]),
        .I4(\i_/badr[6]_INST_0_i_26_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_96 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [9]),
        .I2(gr0_bus1),
        .I3(out[9]),
        .I4(\i_/badr[9]_INST_0_i_26_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/rgf_c0bus_wb[4]_i_99 
       (.I0(gr7_bus1),
        .I1(\rgf_c0bus_wb[4]_i_41 [8]),
        .I2(gr0_bus1),
        .I3(out[8]),
        .I4(\i_/badr[8]_INST_0_i_26_n_0 ),
        .O(\grn_reg[8]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_30
   (p_1_in1_in,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[14] ,
    \grn_reg[14]_0 ,
    \grn_reg[13] ,
    \grn_reg[13]_0 ,
    \grn_reg[12] ,
    \grn_reg[12]_0 ,
    \grn_reg[11] ,
    \grn_reg[11]_0 ,
    \grn_reg[10] ,
    \grn_reg[10]_0 ,
    \grn_reg[9] ,
    \grn_reg[9]_0 ,
    \grn_reg[8] ,
    \grn_reg[8]_0 ,
    \grn_reg[7] ,
    \grn_reg[7]_0 ,
    \grn_reg[6] ,
    \grn_reg[6]_0 ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[3] ,
    \grn_reg[3]_0 ,
    \grn_reg[2] ,
    \grn_reg[2]_0 ,
    \grn_reg[1] ,
    \grn_reg[1]_0 ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \badr[15]_INST_0_i_1 ,
    out,
    \rgf_c1bus_wb[4]_i_47 ,
    \badr[14]_INST_0_i_1 ,
    \badr[13]_INST_0_i_1 ,
    \badr[12]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1 ,
    \badr[10]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1 ,
    \badr[8]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1 ,
    \badr[4]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \badr[1]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1 ,
    \i_/badr[15]_INST_0_i_4_0 ,
    \i_/badr[15]_INST_0_i_19_0 ,
    \i_/badr[15]_INST_0_i_19_1 ,
    \i_/badr[15]_INST_0_i_19_2 ,
    \rgf_c1bus_wb[4]_i_47_0 ,
    \rgf_c1bus_wb[4]_i_47_1 ,
    a1bus_sel_0,
    \i_/badr[15]_INST_0_i_19_3 ,
    \i_/badr[15]_INST_0_i_19_4 ,
    bank_sel);
  output [15:0]p_1_in1_in;
  output \grn_reg[15] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14] ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13] ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12] ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11] ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10] ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9] ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8] ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7] ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6] ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3] ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2] ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1] ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0] ;
  output \grn_reg[0]_0 ;
  input \badr[15]_INST_0_i_1 ;
  input [15:0]out;
  input [15:0]\rgf_c1bus_wb[4]_i_47 ;
  input \badr[14]_INST_0_i_1 ;
  input \badr[13]_INST_0_i_1 ;
  input \badr[12]_INST_0_i_1 ;
  input \badr[11]_INST_0_i_1 ;
  input \badr[10]_INST_0_i_1 ;
  input \badr[9]_INST_0_i_1 ;
  input \badr[8]_INST_0_i_1 ;
  input \badr[7]_INST_0_i_1 ;
  input \badr[6]_INST_0_i_1 ;
  input \badr[5]_INST_0_i_1 ;
  input \badr[4]_INST_0_i_1 ;
  input \badr[3]_INST_0_i_1 ;
  input \badr[2]_INST_0_i_1 ;
  input \badr[1]_INST_0_i_1 ;
  input \badr[0]_INST_0_i_1 ;
  input [1:0]\i_/badr[15]_INST_0_i_4_0 ;
  input \i_/badr[15]_INST_0_i_19_0 ;
  input \i_/badr[15]_INST_0_i_19_1 ;
  input \i_/badr[15]_INST_0_i_19_2 ;
  input [15:0]\rgf_c1bus_wb[4]_i_47_0 ;
  input [15:0]\rgf_c1bus_wb[4]_i_47_1 ;
  input [1:0]a1bus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_19_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_19_4 ;
  input [0:0]bank_sel;

  wire [1:0]a1bus_sel_0;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1 ;
  wire [0:0]bank_sel;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_33_n_0 ;
  wire \i_/badr[10]_INST_0_i_32_n_0 ;
  wire \i_/badr[11]_INST_0_i_33_n_0 ;
  wire \i_/badr[12]_INST_0_i_32_n_0 ;
  wire \i_/badr[13]_INST_0_i_32_n_0 ;
  wire \i_/badr[14]_INST_0_i_32_n_0 ;
  wire \i_/badr[15]_INST_0_i_19_0 ;
  wire \i_/badr[15]_INST_0_i_19_1 ;
  wire \i_/badr[15]_INST_0_i_19_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_19_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_19_4 ;
  wire [1:0]\i_/badr[15]_INST_0_i_4_0 ;
  wire \i_/badr[15]_INST_0_i_65_n_0 ;
  wire \i_/badr[1]_INST_0_i_32_n_0 ;
  wire \i_/badr[2]_INST_0_i_32_n_0 ;
  wire \i_/badr[3]_INST_0_i_33_n_0 ;
  wire \i_/badr[4]_INST_0_i_32_n_0 ;
  wire \i_/badr[5]_INST_0_i_32_n_0 ;
  wire \i_/badr[6]_INST_0_i_32_n_0 ;
  wire \i_/badr[7]_INST_0_i_33_n_0 ;
  wire \i_/badr[8]_INST_0_i_32_n_0 ;
  wire \i_/badr[9]_INST_0_i_32_n_0 ;
  wire [15:0]out;
  wire [15:0]p_1_in1_in;
  wire [15:0]\rgf_c1bus_wb[4]_i_47 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_47_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_47_1 ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_33_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [0]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [0]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[0]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[0]_INST_0_i_4 
       (.I0(\badr[0]_INST_0_i_1 ),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [0]),
        .I4(gr7_bus1),
        .I5(\grn_reg[0] ),
        .O(p_1_in1_in[0]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_32_n_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [10]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [10]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[10]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[10]_INST_0_i_4 
       (.I0(\badr[10]_INST_0_i_1 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [10]),
        .I4(gr7_bus1),
        .I5(\grn_reg[10] ),
        .O(p_1_in1_in[10]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_33_n_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [11]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [11]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[11]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[11]_INST_0_i_4 
       (.I0(\badr[11]_INST_0_i_1 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [11]),
        .I4(gr7_bus1),
        .I5(\grn_reg[11] ),
        .O(p_1_in1_in[11]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_32_n_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [12]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [12]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[12]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[12]_INST_0_i_4 
       (.I0(\badr[12]_INST_0_i_1 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [12]),
        .I4(gr7_bus1),
        .I5(\grn_reg[12] ),
        .O(p_1_in1_in[12]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_32_n_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [13]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [13]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[13]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[13]_INST_0_i_4 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [13]),
        .I4(gr7_bus1),
        .I5(\grn_reg[13] ),
        .O(p_1_in1_in[13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_32_n_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [14]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [14]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[14]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[14]_INST_0_i_4 
       (.I0(\badr[14]_INST_0_i_1 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [14]),
        .I4(gr7_bus1),
        .I5(\grn_reg[14] ),
        .O(p_1_in1_in[14]));
  LUT5 #(
    .INIT(32'h00000001)) 
    \i_/badr[15]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_4_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_4_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_19_0 ),
        .I3(\i_/badr[15]_INST_0_i_19_1 ),
        .I4(\i_/badr[15]_INST_0_i_19_2 ),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_4_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_4_0 [0]),
        .I2(a1bus_sel_0[1]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_65_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[15]_INST_0_i_4 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [15]),
        .I4(gr7_bus1),
        .I5(\grn_reg[15] ),
        .O(p_1_in1_in[15]));
  LUT5 #(
    .INIT(32'h00001000)) 
    \i_/badr[15]_INST_0_i_63 
       (.I0(\i_/badr[15]_INST_0_i_4_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_4_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_19_0 ),
        .I3(\i_/badr[15]_INST_0_i_19_1 ),
        .I4(\i_/badr[15]_INST_0_i_19_2 ),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/badr[15]_INST_0_i_64 
       (.I0(\i_/badr[15]_INST_0_i_4_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_4_0 [0]),
        .I2(a1bus_sel_0[0]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_65 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [15]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [15]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[15]_INST_0_i_65_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_32_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [1]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [1]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[1]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[1]_INST_0_i_4 
       (.I0(\badr[1]_INST_0_i_1 ),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [1]),
        .I4(gr7_bus1),
        .I5(\grn_reg[1] ),
        .O(p_1_in1_in[1]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_32_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [2]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [2]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[2]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[2]_INST_0_i_4 
       (.I0(\badr[2]_INST_0_i_1 ),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [2]),
        .I4(gr7_bus1),
        .I5(\grn_reg[2] ),
        .O(p_1_in1_in[2]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_33_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [3]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [3]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[3]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[3]_INST_0_i_4 
       (.I0(\badr[3]_INST_0_i_1 ),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [3]),
        .I4(gr7_bus1),
        .I5(\grn_reg[3] ),
        .O(p_1_in1_in[3]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_32_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [4]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [4]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[4]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[4]_INST_0_i_4 
       (.I0(\badr[4]_INST_0_i_1 ),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [4]),
        .I4(gr7_bus1),
        .I5(\grn_reg[4] ),
        .O(p_1_in1_in[4]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_32_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [5]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [5]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[5]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[5]_INST_0_i_4 
       (.I0(\badr[5]_INST_0_i_1 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [5]),
        .I4(gr7_bus1),
        .I5(\grn_reg[5] ),
        .O(p_1_in1_in[5]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_32_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [6]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [6]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[6]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[6]_INST_0_i_4 
       (.I0(\badr[6]_INST_0_i_1 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [6]),
        .I4(gr7_bus1),
        .I5(\grn_reg[6] ),
        .O(p_1_in1_in[6]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_33_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [7]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [7]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[7]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[7]_INST_0_i_4 
       (.I0(\badr[7]_INST_0_i_1 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [7]),
        .I4(gr7_bus1),
        .I5(\grn_reg[7] ),
        .O(p_1_in1_in[7]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_32_n_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [8]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [8]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[8]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[8]_INST_0_i_4 
       (.I0(\badr[8]_INST_0_i_1 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [8]),
        .I4(gr7_bus1),
        .I5(\grn_reg[8] ),
        .O(p_1_in1_in[8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47_0 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_32_n_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_19_3 [9]),
        .I1(\i_/badr[15]_INST_0_i_19_4 [9]),
        .I2(bank_sel),
        .I3(\i_/badr[15]_INST_0_i_19_0 ),
        .I4(\i_/badr[15]_INST_0_i_19_1 ),
        .I5(\i_/badr[15]_INST_0_i_19_2 ),
        .O(\i_/badr[9]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[9]_INST_0_i_4 
       (.I0(\badr[9]_INST_0_i_1 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47 [9]),
        .I4(gr7_bus1),
        .I5(\grn_reg[9] ),
        .O(p_1_in1_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_104 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_108 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_111 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_116 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_119 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_124 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_127 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_132 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_68 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_73 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_76 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_81 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_84 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_89 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_92 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_99 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_47 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_31
   (p_0_in0_in,
    \grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \sr_reg[0] ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_0 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_0 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_0 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_0 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_0 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_0 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_0 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_0 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_0 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_0 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_0 ,
    \grn_reg[0]_1 ,
    \badr[15]_INST_0_i_1 ,
    out,
    \rgf_c1bus_wb[4]_i_39 ,
    \rgf_c1bus_wb[4]_i_47 ,
    \rgf_c1bus_wb[4]_i_47_0 ,
    \badr[14]_INST_0_i_1 ,
    \badr[13]_INST_0_i_1 ,
    \badr[12]_INST_0_i_1 ,
    \badr[11]_INST_0_i_1 ,
    \badr[10]_INST_0_i_1 ,
    \badr[9]_INST_0_i_1 ,
    \badr[8]_INST_0_i_1 ,
    \badr[7]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1 ,
    \badr[4]_INST_0_i_1 ,
    \badr[3]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \badr[1]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1 ,
    \badr[15]_INST_0_i_20 ,
    \i_/badr[0]_INST_0_i_17_0 ,
    \i_/badr[0]_INST_0_i_17_1 ,
    \i_/badr[0]_INST_0_i_17_2 ,
    \rgf_c1bus_wb[4]_i_47_1 ,
    \rgf_c1bus_wb[4]_i_47_2 ,
    \rgf_c1bus_wb[4]_i_47_3 ,
    \rgf_c1bus_wb[4]_i_41 ,
    \rgf_c1bus_wb[4]_i_41_0 ,
    \rgf_c1bus_wb[4]_i_51 ,
    \rgf_c1bus_wb[4]_i_51_0 ,
    \sr[4]_i_235 ,
    \sr[4]_i_235_0 ,
    \rgf_c1bus_wb[4]_i_65 ,
    \rgf_c1bus_wb[4]_i_65_0 ,
    \sr[4]_i_237 ,
    \sr[4]_i_237_0 ,
    \rgf_c1bus_wb[4]_i_61 ,
    \rgf_c1bus_wb[4]_i_61_0 ,
    \rgf_c1bus_wb[4]_i_57 ,
    \rgf_c1bus_wb[4]_i_57_0 ,
    \sr[4]_i_245 ,
    \sr[4]_i_245_0 ,
    \rgf_c1bus_wb[4]_i_53 ,
    \rgf_c1bus_wb[4]_i_53_0 ,
    \sr[4]_i_243 ,
    \sr[4]_i_243_0 ,
    \rgf_c1bus_wb[4]_i_33 ,
    \rgf_c1bus_wb[4]_i_33_0 ,
    \rgf_c1bus_wb[4]_i_67 ,
    \rgf_c1bus_wb[4]_i_67_0 ,
    \rgf_c1bus_wb[4]_i_37 ,
    \rgf_c1bus_wb[4]_i_37_0 ,
    \sr[4]_i_240 ,
    \sr[4]_i_240_0 ,
    a1bus_sel_0,
    \i_/badr[15]_INST_0_i_23_0 ,
    \i_/badr[15]_INST_0_i_23_1 ,
    \i_/badr[15]_INST_0_i_23_2 );
  output [15:0]p_0_in0_in;
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \sr_reg[0] ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[0]_1 ;
  input \badr[15]_INST_0_i_1 ;
  input [15:0]out;
  input [15:0]\rgf_c1bus_wb[4]_i_39 ;
  input [15:0]\rgf_c1bus_wb[4]_i_47 ;
  input [15:0]\rgf_c1bus_wb[4]_i_47_0 ;
  input \badr[14]_INST_0_i_1 ;
  input \badr[13]_INST_0_i_1 ;
  input \badr[12]_INST_0_i_1 ;
  input \badr[11]_INST_0_i_1 ;
  input \badr[10]_INST_0_i_1 ;
  input \badr[9]_INST_0_i_1 ;
  input \badr[8]_INST_0_i_1 ;
  input \badr[7]_INST_0_i_1 ;
  input \badr[6]_INST_0_i_1 ;
  input \badr[5]_INST_0_i_1 ;
  input \badr[4]_INST_0_i_1 ;
  input \badr[3]_INST_0_i_1 ;
  input \badr[2]_INST_0_i_1 ;
  input \badr[1]_INST_0_i_1 ;
  input \badr[0]_INST_0_i_1 ;
  input [1:0]\badr[15]_INST_0_i_20 ;
  input \i_/badr[0]_INST_0_i_17_0 ;
  input \i_/badr[0]_INST_0_i_17_1 ;
  input \i_/badr[0]_INST_0_i_17_2 ;
  input \rgf_c1bus_wb[4]_i_47_1 ;
  input \rgf_c1bus_wb[4]_i_47_2 ;
  input [14:0]\rgf_c1bus_wb[4]_i_47_3 ;
  input \rgf_c1bus_wb[4]_i_41 ;
  input \rgf_c1bus_wb[4]_i_41_0 ;
  input \rgf_c1bus_wb[4]_i_51 ;
  input \rgf_c1bus_wb[4]_i_51_0 ;
  input \sr[4]_i_235 ;
  input \sr[4]_i_235_0 ;
  input \rgf_c1bus_wb[4]_i_65 ;
  input \rgf_c1bus_wb[4]_i_65_0 ;
  input \sr[4]_i_237 ;
  input \sr[4]_i_237_0 ;
  input \rgf_c1bus_wb[4]_i_61 ;
  input \rgf_c1bus_wb[4]_i_61_0 ;
  input \rgf_c1bus_wb[4]_i_57 ;
  input \rgf_c1bus_wb[4]_i_57_0 ;
  input \sr[4]_i_245 ;
  input \sr[4]_i_245_0 ;
  input \rgf_c1bus_wb[4]_i_53 ;
  input \rgf_c1bus_wb[4]_i_53_0 ;
  input \sr[4]_i_243 ;
  input \sr[4]_i_243_0 ;
  input \rgf_c1bus_wb[4]_i_33 ;
  input \rgf_c1bus_wb[4]_i_33_0 ;
  input \rgf_c1bus_wb[4]_i_67 ;
  input \rgf_c1bus_wb[4]_i_67_0 ;
  input \rgf_c1bus_wb[4]_i_37 ;
  input \rgf_c1bus_wb[4]_i_37_0 ;
  input \sr[4]_i_240 ;
  input \sr[4]_i_240_0 ;
  input [2:0]a1bus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_23_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_23_1 ;
  input \i_/badr[15]_INST_0_i_23_2 ;

  wire [2:0]a1bus_sel_0;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1 ;
  wire [1:0]\badr[15]_INST_0_i_20 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[7]_INST_0_i_1 ;
  wire \badr[8]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \i_/badr[0]_INST_0_i_17_0 ;
  wire \i_/badr[0]_INST_0_i_17_1 ;
  wire \i_/badr[0]_INST_0_i_17_2 ;
  wire \i_/badr[0]_INST_0_i_34_n_0 ;
  wire \i_/badr[10]_INST_0_i_33_n_0 ;
  wire \i_/badr[11]_INST_0_i_34_n_0 ;
  wire \i_/badr[12]_INST_0_i_33_n_0 ;
  wire \i_/badr[13]_INST_0_i_33_n_0 ;
  wire \i_/badr[14]_INST_0_i_33_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_23_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_23_1 ;
  wire \i_/badr[15]_INST_0_i_23_2 ;
  wire \i_/badr[15]_INST_0_i_69_n_0 ;
  wire \i_/badr[1]_INST_0_i_33_n_0 ;
  wire \i_/badr[2]_INST_0_i_33_n_0 ;
  wire \i_/badr[3]_INST_0_i_34_n_0 ;
  wire \i_/badr[4]_INST_0_i_33_n_0 ;
  wire \i_/badr[5]_INST_0_i_33_n_0 ;
  wire \i_/badr[6]_INST_0_i_33_n_0 ;
  wire \i_/badr[7]_INST_0_i_34_n_0 ;
  wire \i_/badr[8]_INST_0_i_33_n_0 ;
  wire \i_/badr[9]_INST_0_i_33_n_0 ;
  wire [15:0]out;
  wire [15:0]p_0_in0_in;
  wire \rgf_c1bus_wb[4]_i_33 ;
  wire \rgf_c1bus_wb[4]_i_33_0 ;
  wire \rgf_c1bus_wb[4]_i_37 ;
  wire \rgf_c1bus_wb[4]_i_37_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_39 ;
  wire \rgf_c1bus_wb[4]_i_41 ;
  wire \rgf_c1bus_wb[4]_i_41_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_47 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_47_0 ;
  wire \rgf_c1bus_wb[4]_i_47_1 ;
  wire \rgf_c1bus_wb[4]_i_47_2 ;
  wire [14:0]\rgf_c1bus_wb[4]_i_47_3 ;
  wire \rgf_c1bus_wb[4]_i_51 ;
  wire \rgf_c1bus_wb[4]_i_51_0 ;
  wire \rgf_c1bus_wb[4]_i_53 ;
  wire \rgf_c1bus_wb[4]_i_53_0 ;
  wire \rgf_c1bus_wb[4]_i_57 ;
  wire \rgf_c1bus_wb[4]_i_57_0 ;
  wire \rgf_c1bus_wb[4]_i_61 ;
  wire \rgf_c1bus_wb[4]_i_61_0 ;
  wire \rgf_c1bus_wb[4]_i_65 ;
  wire \rgf_c1bus_wb[4]_i_65_0 ;
  wire \rgf_c1bus_wb[4]_i_67 ;
  wire \rgf_c1bus_wb[4]_i_67_0 ;
  wire \sr[4]_i_235 ;
  wire \sr[4]_i_235_0 ;
  wire \sr[4]_i_237 ;
  wire \sr[4]_i_237_0 ;
  wire \sr[4]_i_240 ;
  wire \sr[4]_i_240_0 ;
  wire \sr[4]_i_243 ;
  wire \sr[4]_i_243_0 ;
  wire \sr[4]_i_245 ;
  wire \sr[4]_i_245_0 ;
  wire \sr_reg[0] ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [0]),
        .I4(\i_/badr[0]_INST_0_i_34_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [0]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[0]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[0]_INST_0_i_5 
       (.I0(\badr[0]_INST_0_i_1 ),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [0]),
        .I4(gr7_bus1),
        .I5(\grn_reg[0] ),
        .O(p_0_in0_in[0]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [10]),
        .I4(\i_/badr[10]_INST_0_i_33_n_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [10]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[10]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[10]_INST_0_i_5 
       (.I0(\badr[10]_INST_0_i_1 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [10]),
        .I4(gr7_bus1),
        .I5(\grn_reg[10] ),
        .O(p_0_in0_in[10]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [11]),
        .I4(\i_/badr[11]_INST_0_i_34_n_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [11]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[11]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[11]_INST_0_i_5 
       (.I0(\badr[11]_INST_0_i_1 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [11]),
        .I4(gr7_bus1),
        .I5(\grn_reg[11] ),
        .O(p_0_in0_in[11]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [12]),
        .I4(\i_/badr[12]_INST_0_i_33_n_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [12]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[12]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[12]_INST_0_i_5 
       (.I0(\badr[12]_INST_0_i_1 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [12]),
        .I4(gr7_bus1),
        .I5(\grn_reg[12] ),
        .O(p_0_in0_in[12]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [13]),
        .I4(\i_/badr[13]_INST_0_i_33_n_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [13]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[13]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[13]_INST_0_i_5 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [13]),
        .I4(gr7_bus1),
        .I5(\grn_reg[13] ),
        .O(p_0_in0_in[13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [14]),
        .I4(\i_/badr[14]_INST_0_i_33_n_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [14]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[14]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[14]_INST_0_i_5 
       (.I0(\badr[14]_INST_0_i_1 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [14]),
        .I4(gr7_bus1),
        .I5(\grn_reg[14] ),
        .O(p_0_in0_in[14]));
  LUT5 #(
    .INIT(32'h00000004)) 
    \i_/badr[15]_INST_0_i_21 
       (.I0(\badr[15]_INST_0_i_20 [0]),
        .I1(\badr[15]_INST_0_i_20 [1]),
        .I2(\i_/badr[0]_INST_0_i_17_0 ),
        .I3(\i_/badr[0]_INST_0_i_17_1 ),
        .I4(\i_/badr[0]_INST_0_i_17_2 ),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_20 [0]),
        .I1(\badr[15]_INST_0_i_20 [1]),
        .I2(a1bus_sel_0[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [15]),
        .I4(\i_/badr[15]_INST_0_i_69_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[15]_INST_0_i_5 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [15]),
        .I4(gr7_bus1),
        .I5(\grn_reg[15] ),
        .O(p_0_in0_in[15]));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_66 
       (.I0(\badr[15]_INST_0_i_20 [0]),
        .I1(\badr[15]_INST_0_i_20 [1]),
        .I2(a1bus_sel_0[1]),
        .O(\sr_reg[0] ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \i_/badr[15]_INST_0_i_67 
       (.I0(\badr[15]_INST_0_i_20 [0]),
        .I1(\badr[15]_INST_0_i_20 [1]),
        .I2(\i_/badr[0]_INST_0_i_17_0 ),
        .I3(\i_/badr[0]_INST_0_i_17_1 ),
        .I4(\i_/badr[0]_INST_0_i_17_2 ),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_68 
       (.I0(\badr[15]_INST_0_i_20 [0]),
        .I1(\badr[15]_INST_0_i_20 [1]),
        .I2(a1bus_sel_0[0]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_69 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [15]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[15]_INST_0_i_69_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [1]),
        .I4(\i_/badr[1]_INST_0_i_33_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [1]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[1]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[1]_INST_0_i_5 
       (.I0(\badr[1]_INST_0_i_1 ),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [1]),
        .I4(gr7_bus1),
        .I5(\grn_reg[1] ),
        .O(p_0_in0_in[1]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [2]),
        .I4(\i_/badr[2]_INST_0_i_33_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [2]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[2]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[2]_INST_0_i_5 
       (.I0(\badr[2]_INST_0_i_1 ),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [2]),
        .I4(gr7_bus1),
        .I5(\grn_reg[2] ),
        .O(p_0_in0_in[2]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [3]),
        .I4(\i_/badr[3]_INST_0_i_34_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [3]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[3]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[3]_INST_0_i_5 
       (.I0(\badr[3]_INST_0_i_1 ),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [3]),
        .I4(gr7_bus1),
        .I5(\grn_reg[3] ),
        .O(p_0_in0_in[3]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [4]),
        .I4(\i_/badr[4]_INST_0_i_33_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [4]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[4]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[4]_INST_0_i_5 
       (.I0(\badr[4]_INST_0_i_1 ),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [4]),
        .I4(gr7_bus1),
        .I5(\grn_reg[4] ),
        .O(p_0_in0_in[4]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [5]),
        .I4(\i_/badr[5]_INST_0_i_33_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [5]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[5]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[5]_INST_0_i_5 
       (.I0(\badr[5]_INST_0_i_1 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [5]),
        .I4(gr7_bus1),
        .I5(\grn_reg[5] ),
        .O(p_0_in0_in[5]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [6]),
        .I4(\i_/badr[6]_INST_0_i_33_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [6]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[6]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[6]_INST_0_i_5 
       (.I0(\badr[6]_INST_0_i_1 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [6]),
        .I4(gr7_bus1),
        .I5(\grn_reg[6] ),
        .O(p_0_in0_in[6]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [7]),
        .I4(\i_/badr[7]_INST_0_i_34_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [7]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[7]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[7]_INST_0_i_5 
       (.I0(\badr[7]_INST_0_i_1 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [7]),
        .I4(gr7_bus1),
        .I5(\grn_reg[7] ),
        .O(p_0_in0_in[7]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [8]),
        .I4(\i_/badr[8]_INST_0_i_33_n_0 ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [8]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[8]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[8]_INST_0_i_5 
       (.I0(\badr[8]_INST_0_i_1 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [8]),
        .I4(gr7_bus1),
        .I5(\grn_reg[8] ),
        .O(p_0_in0_in[8]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_47 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_47_0 [9]),
        .I4(\i_/badr[9]_INST_0_i_33_n_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_23_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_23_1 [9]),
        .I2(\i_/badr[15]_INST_0_i_23_2 ),
        .I3(\i_/badr[0]_INST_0_i_17_0 ),
        .I4(\i_/badr[0]_INST_0_i_17_1 ),
        .I5(\i_/badr[0]_INST_0_i_17_2 ),
        .O(\i_/badr[9]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/badr[9]_INST_0_i_5 
       (.I0(\badr[9]_INST_0_i_1 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\rgf_c1bus_wb[4]_i_39 [9]),
        .I4(gr7_bus1),
        .I5(\grn_reg[9] ),
        .O(p_0_in0_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_100 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_103 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [13]),
        .I2(\rgf_c1bus_wb[4]_i_51 ),
        .I3(\rgf_c1bus_wb[4]_i_51_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [12]),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_107 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [5]),
        .I2(\rgf_c1bus_wb[4]_i_53 ),
        .I3(\rgf_c1bus_wb[4]_i_53_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [5]),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_112 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_115 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [7]),
        .I2(\rgf_c1bus_wb[4]_i_57 ),
        .I3(\rgf_c1bus_wb[4]_i_57_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [7]),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_120 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_123 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [9]),
        .I2(\rgf_c1bus_wb[4]_i_61 ),
        .I3(\rgf_c1bus_wb[4]_i_61_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [8]),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_128 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_131 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [11]),
        .I2(\rgf_c1bus_wb[4]_i_65 ),
        .I3(\rgf_c1bus_wb[4]_i_65_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [10]),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_133 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_134 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [2]),
        .I2(\rgf_c1bus_wb[4]_i_67 ),
        .I3(\rgf_c1bus_wb[4]_i_67_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [2]),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_69 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_72 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [3]),
        .I2(\rgf_c1bus_wb[4]_i_33 ),
        .I3(\rgf_c1bus_wb[4]_i_33_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [3]),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_77 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_80 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [1]),
        .I2(\rgf_c1bus_wb[4]_i_37 ),
        .I3(\rgf_c1bus_wb[4]_i_37_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [1]),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_85 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_88 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [14]),
        .I2(\rgf_c1bus_wb[4]_i_41 ),
        .I3(\rgf_c1bus_wb[4]_i_41_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [13]),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_93 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c1bus_wb[4]_i_95 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_96 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [15]),
        .I2(\rgf_c1bus_wb[4]_i_47_1 ),
        .I3(\rgf_c1bus_wb[4]_i_47_2 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [14]),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/sr[4]_i_246 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/sr[4]_i_247 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [12]),
        .I2(\sr[4]_i_235 ),
        .I3(\sr[4]_i_235_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [11]),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/sr[4]_i_248 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/sr[4]_i_249 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [10]),
        .I2(\sr[4]_i_237 ),
        .I3(\sr[4]_i_237_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [9]),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/sr[4]_i_250 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/sr[4]_i_252 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [0]),
        .I2(\sr[4]_i_240 ),
        .I3(\sr[4]_i_240_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [0]),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/sr[4]_i_253 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/sr[4]_i_254 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/sr[4]_i_255 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [4]),
        .I2(\sr[4]_i_243 ),
        .I3(\sr[4]_i_243_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [4]),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/sr[4]_i_256 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_39 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_1 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/sr[4]_i_257 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_39 [6]),
        .I2(\sr[4]_i_245 ),
        .I3(\sr[4]_i_245_0 ),
        .I4(\sr_reg[0] ),
        .I5(\rgf_c1bus_wb[4]_i_47_3 [6]),
        .O(\grn_reg[6]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_32
   (p_1_in3_in,
    \grn_reg[4] ,
    out,
    \bdatw[15]_INST_0_i_1 ,
    \i_/bdatw[15]_INST_0_i_9_0 ,
    \bbus_o[4]_INST_0_i_1 ,
    \bbus_o[3]_INST_0_i_1 ,
    \bbus_o[2]_INST_0_i_1 ,
    \bbus_o[1]_INST_0_i_1 ,
    \bbus_o[0]_INST_0_i_1 ,
    bank_sel,
    \i_/bdatw[15]_INST_0_i_9_1 ,
    \i_/bdatw[15]_INST_0_i_9_2 ,
    \i_/bdatw[15]_INST_0_i_9_3 ,
    \i_/bdatw[15]_INST_0_i_9_4 ,
    ctl_selb0_0,
    \i_/bdatw[15]_INST_0_i_9_5 ,
    \i_/bdatw[15]_INST_0_i_9_6 ,
    \i_/bdatw[15]_INST_0_i_24_0 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_9_7 ,
    \i_/bdatw[15]_INST_0_i_27_0 ,
    \i_/bdatw[15]_INST_0_i_27_1 ,
    \i_/bdatw[15]_INST_0_i_77_0 ,
    \i_/bdatw[15]_INST_0_i_27_2 ,
    b0bus_sel_0,
    \i_/bdatw[15]_INST_0_i_9_8 ,
    \i_/bdatw[15]_INST_0_i_24_1 );
  output [10:0]p_1_in3_in;
  output [4:0]\grn_reg[4] ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_9_0 ;
  input \bbus_o[4]_INST_0_i_1 ;
  input \bbus_o[3]_INST_0_i_1 ;
  input \bbus_o[2]_INST_0_i_1 ;
  input \bbus_o[1]_INST_0_i_1 ;
  input \bbus_o[0]_INST_0_i_1 ;
  input [0:0]bank_sel;
  input \i_/bdatw[15]_INST_0_i_9_1 ;
  input \i_/bdatw[15]_INST_0_i_9_2 ;
  input \i_/bdatw[15]_INST_0_i_9_3 ;
  input \i_/bdatw[15]_INST_0_i_9_4 ;
  input [0:0]ctl_selb0_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_9_5 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_9_6 ;
  input \i_/bdatw[15]_INST_0_i_24_0 ;
  input [1:0]ctl_selb0_rn;
  input [10:0]\i_/bdatw[15]_INST_0_i_9_7 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_1 ;
  input \i_/bdatw[15]_INST_0_i_77_0 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_27_2 ;
  input [1:0]b0bus_sel_0;
  input \i_/bdatw[15]_INST_0_i_9_8 ;
  input \i_/bdatw[15]_INST_0_i_24_1 ;

  wire [1:0]b0bus_sel_0;
  wire [0:0]bank_sel;
  wire \bbus_o[0]_INST_0_i_1 ;
  wire \bbus_o[1]_INST_0_i_1 ;
  wire \bbus_o[2]_INST_0_i_1 ;
  wire \bbus_o[3]_INST_0_i_1 ;
  wire \bbus_o[4]_INST_0_i_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_1 ;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [4:0]\grn_reg[4] ;
  wire \i_/bbus_o[0]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[0]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[0]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_11_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_8_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_13_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_19_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_19_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_9_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_10_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_19_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_9_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_24_0 ;
  wire \i_/bdatw[15]_INST_0_i_24_1 ;
  wire \i_/bdatw[15]_INST_0_i_24_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_1 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_27_2 ;
  wire \i_/bdatw[15]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_77_0 ;
  wire \i_/bdatw[15]_INST_0_i_77_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_9_0 ;
  wire \i_/bdatw[15]_INST_0_i_9_1 ;
  wire \i_/bdatw[15]_INST_0_i_9_2 ;
  wire \i_/bdatw[15]_INST_0_i_9_3 ;
  wire \i_/bdatw[15]_INST_0_i_9_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_9_5 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_9_6 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_9_7 ;
  wire \i_/bdatw[15]_INST_0_i_9_8 ;
  wire \i_/bdatw[8]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_18_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_19_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_45_n_0 ;
  wire [15:0]out;
  wire [10:0]p_1_in3_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_10 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [0]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[0]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_12 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [0]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [0]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[0]_INST_0_i_5 
       (.I0(\i_/bbus_o[0]_INST_0_i_9_n_0 ),
        .I1(\i_/bbus_o[0]_INST_0_i_10_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_0 [0]),
        .I3(gr2_bus1),
        .I4(\bbus_o[0]_INST_0_i_1 ),
        .I5(\i_/bbus_o[0]_INST_0_i_12_n_0 ),
        .O(\grn_reg[4] [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [0]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[0]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [1]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [1]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[1]_INST_0_i_5 
       (.I0(\i_/bbus_o[1]_INST_0_i_8_n_0 ),
        .I1(\i_/bbus_o[1]_INST_0_i_9_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_0 [1]),
        .I3(gr2_bus1),
        .I4(\bbus_o[1]_INST_0_i_1 ),
        .I5(\i_/bbus_o[1]_INST_0_i_11_n_0 ),
        .O(\grn_reg[4] [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_8 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [1]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[1]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_9 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [1]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[1]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_10 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [2]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[2]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_12 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [2]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [2]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[2]_INST_0_i_5 
       (.I0(\i_/bbus_o[2]_INST_0_i_9_n_0 ),
        .I1(\i_/bbus_o[2]_INST_0_i_10_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_0 [2]),
        .I3(gr2_bus1),
        .I4(\bbus_o[2]_INST_0_i_1 ),
        .I5(\i_/bbus_o[2]_INST_0_i_12_n_0 ),
        .O(\grn_reg[4] [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [2]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[2]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_10 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [3]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[3]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_12 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [3]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [3]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[3]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[3]_INST_0_i_5 
       (.I0(\i_/bbus_o[3]_INST_0_i_9_n_0 ),
        .I1(\i_/bbus_o[3]_INST_0_i_10_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_0 [3]),
        .I3(gr2_bus1),
        .I4(\bbus_o[3]_INST_0_i_1 ),
        .I5(\i_/bbus_o[3]_INST_0_i_12_n_0 ),
        .O(\grn_reg[4] [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [3]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[3]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_10 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [4]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[4]_INST_0_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bbus_o[4]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_27_2 [0]),
        .I2(b0bus_sel_0[1]),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_13 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [4]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [4]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[4]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_27 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_77_0 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I4(\i_/bdatw[15]_INST_0_i_9_4 ),
        .I5(ctl_selb0_0),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_28 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_9_8 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 ),
        .I3(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I4(\i_/bdatw[15]_INST_0_i_9_4 ),
        .I5(ctl_selb0_0),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[4]_INST_0_i_5 
       (.I0(\i_/bbus_o[4]_INST_0_i_9_n_0 ),
        .I1(\i_/bbus_o[4]_INST_0_i_10_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_0 [4]),
        .I3(gr2_bus1),
        .I4(\bbus_o[4]_INST_0_i_1 ),
        .I5(\i_/bbus_o[4]_INST_0_i_13_n_0 ),
        .O(\grn_reg[4] [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [4]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[4]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bbus_o[5]_INST_0_i_10 
       (.I0(\i_/bbus_o[5]_INST_0_i_19_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [0]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [5]),
        .O(\i_/bbus_o[5]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [5]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [5]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[5]_INST_0_i_5 
       (.I0(\i_/bbus_o[5]_INST_0_i_9_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[5]_INST_0_i_10_n_0 ),
        .O(p_1_in3_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [5]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bbus_o[6]_INST_0_i_10 
       (.I0(\i_/bbus_o[6]_INST_0_i_19_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [1]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [6]),
        .O(\i_/bbus_o[6]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [6]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [6]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[6]_INST_0_i_5 
       (.I0(\i_/bbus_o[6]_INST_0_i_9_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[6]_INST_0_i_10_n_0 ),
        .O(p_1_in3_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [6]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bbus_o[7]_INST_0_i_10 
       (.I0(\i_/bbus_o[7]_INST_0_i_19_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [2]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [7]),
        .O(\i_/bbus_o[7]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [7]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [7]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[7]_INST_0_i_5 
       (.I0(\i_/bbus_o[7]_INST_0_i_9_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[7]_INST_0_i_10_n_0 ),
        .O(p_1_in3_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [7]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_20 
       (.I0(\i_/bdatw[10]_INST_0_i_46_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [5]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [10]),
        .O(\i_/bdatw[10]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [10]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [10]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[10]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_7 
       (.I0(\i_/bdatw[10]_INST_0_i_19_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_20_n_0 ),
        .O(p_1_in3_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_19 
       (.I0(\i_/bdatw[11]_INST_0_i_46_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [6]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [11]),
        .O(\i_/bdatw[11]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [11]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [11]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[11]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_7 
       (.I0(\i_/bdatw[11]_INST_0_i_18_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_19_n_0 ),
        .O(p_1_in3_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_19 
       (.I0(\i_/bdatw[12]_INST_0_i_44_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [7]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [12]),
        .O(\i_/bdatw[12]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [12]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [12]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[12]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_7 
       (.I0(\i_/bdatw[12]_INST_0_i_18_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_19_n_0 ),
        .O(p_1_in3_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_19 
       (.I0(\i_/bdatw[13]_INST_0_i_46_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [8]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [13]),
        .O(\i_/bdatw[13]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [13]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [13]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[13]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_7 
       (.I0(\i_/bdatw[13]_INST_0_i_18_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_19_n_0 ),
        .O(p_1_in3_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_20 
       (.I0(\i_/bdatw[14]_INST_0_i_51_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [9]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [14]),
        .O(\i_/bdatw[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [14]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [14]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[14]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_7 
       (.I0(\i_/bdatw[14]_INST_0_i_19_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_20_n_0 ),
        .O(p_1_in3_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_25 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_9_1 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_2 ),
        .I3(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I4(\i_/bdatw[15]_INST_0_i_9_4 ),
        .I5(ctl_selb0_0),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/bdatw[15]_INST_0_i_26 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_9_8 ),
        .I2(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_9_4 ),
        .I4(ctl_selb0_0),
        .I5(\i_/bdatw[15]_INST_0_i_9_2 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_77_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [10]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [15]),
        .O(\i_/bdatw[15]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_72 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I4(\i_/bdatw[15]_INST_0_i_9_4 ),
        .I5(ctl_selb0_0),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_73 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_24_1 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_9_3 ),
        .I4(\i_/bdatw[15]_INST_0_i_9_4 ),
        .I5(ctl_selb0_0),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_77 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [15]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [15]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[15]_INST_0_i_77_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \i_/bdatw[15]_INST_0_i_78 
       (.I0(\i_/bdatw[15]_INST_0_i_27_2 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_27_2 [0]),
        .I2(b0bus_sel_0[0]),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_9 
       (.I0(\i_/bdatw[15]_INST_0_i_24_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_27_n_0 ),
        .O(p_1_in3_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_19 
       (.I0(\i_/bdatw[8]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [3]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [8]),
        .O(\i_/bdatw[8]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [8]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [8]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_7 
       (.I0(\i_/bdatw[8]_INST_0_i_18_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_19_n_0 ),
        .O(p_1_in3_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_9_5 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_6 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_19 
       (.I0(\i_/bdatw[9]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_9_7 [4]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_9_0 [9]),
        .O(\i_/bdatw[9]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 [9]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 [9]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[9]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_7 
       (.I0(\i_/bdatw[9]_INST_0_i_18_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_19_n_0 ),
        .O(p_1_in3_in[4]));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_33
   (p_0_in2_in,
    \grn_reg[4] ,
    out,
    \bdatw[15]_INST_0_i_1 ,
    \i_/bdatw[15]_INST_0_i_10_0 ,
    \i_/bdatw[15]_INST_0_i_10_1 ,
    \i_/bdatw[15]_INST_0_i_31_0 ,
    \i_/bdatw[15]_INST_0_i_31_1 ,
    \bbus_o[4]_INST_0_i_1 ,
    \bbus_o[3]_INST_0_i_1 ,
    \bbus_o[2]_INST_0_i_1 ,
    \bbus_o[1]_INST_0_i_1 ,
    \bbus_o[0]_INST_0_i_1 ,
    \i_/bdatw[15]_INST_0_i_82_0 ,
    \i_/bdatw[15]_INST_0_i_10_2 ,
    \i_/bdatw[15]_INST_0_i_10_3 ,
    \i_/bdatw[15]_INST_0_i_28_0 ,
    \i_/bdatw[15]_INST_0_i_28_1 ,
    ctl_selb0_0,
    \i_/bdatw[15]_INST_0_i_10_4 ,
    \i_/bdatw[15]_INST_0_i_10_5 ,
    \i_/bdatw[15]_INST_0_i_28_2 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_10_6 ,
    \i_/bdatw[15]_INST_0_i_31_2 ,
    b0bus_sel_0,
    \i_/bdatw[15]_INST_0_i_82_1 ,
    \i_/bdatw[15]_INST_0_i_28_3 );
  output [10:0]p_0_in2_in;
  output [4:0]\grn_reg[4] ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_1 ;
  input [10:0]\i_/bdatw[15]_INST_0_i_10_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_10_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_31_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_31_1 ;
  input \bbus_o[4]_INST_0_i_1 ;
  input \bbus_o[3]_INST_0_i_1 ;
  input \bbus_o[2]_INST_0_i_1 ;
  input \bbus_o[1]_INST_0_i_1 ;
  input \bbus_o[0]_INST_0_i_1 ;
  input \i_/bdatw[15]_INST_0_i_82_0 ;
  input \i_/bdatw[15]_INST_0_i_10_2 ;
  input \i_/bdatw[15]_INST_0_i_10_3 ;
  input \i_/bdatw[15]_INST_0_i_28_0 ;
  input \i_/bdatw[15]_INST_0_i_28_1 ;
  input [0:0]ctl_selb0_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_10_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_10_5 ;
  input \i_/bdatw[15]_INST_0_i_28_2 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_10_6 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_31_2 ;
  input [1:0]b0bus_sel_0;
  input \i_/bdatw[15]_INST_0_i_82_1 ;
  input \i_/bdatw[15]_INST_0_i_28_3 ;

  wire [1:0]b0bus_sel_0;
  wire \bbus_o[0]_INST_0_i_1 ;
  wire \bbus_o[1]_INST_0_i_1 ;
  wire \bbus_o[2]_INST_0_i_1 ;
  wire \bbus_o[3]_INST_0_i_1 ;
  wire \bbus_o[4]_INST_0_i_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_1 ;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire [4:0]\grn_reg[4] ;
  wire \i_/bbus_o[0]_INST_0_i_13_n_0 ;
  wire \i_/bbus_o[0]_INST_0_i_14_n_0 ;
  wire \i_/bbus_o[0]_INST_0_i_16_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_13_n_0 ;
  wire \i_/bbus_o[1]_INST_0_i_15_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_13_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_14_n_0 ;
  wire \i_/bbus_o[2]_INST_0_i_16_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_13_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_14_n_0 ;
  wire \i_/bbus_o[3]_INST_0_i_16_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_14_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_15_n_0 ;
  wire \i_/bbus_o[4]_INST_0_i_18_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_11_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_20_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_11_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_20_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_11_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_12_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_52_n_0 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_10_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_10_1 ;
  wire \i_/bdatw[15]_INST_0_i_10_2 ;
  wire \i_/bdatw[15]_INST_0_i_10_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_10_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_10_5 ;
  wire \i_/bdatw[15]_INST_0_i_10_6 ;
  wire \i_/bdatw[15]_INST_0_i_28_0 ;
  wire \i_/bdatw[15]_INST_0_i_28_1 ;
  wire \i_/bdatw[15]_INST_0_i_28_2 ;
  wire \i_/bdatw[15]_INST_0_i_28_3 ;
  wire \i_/bdatw[15]_INST_0_i_28_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_31_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_31_1 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_31_2 ;
  wire \i_/bdatw[15]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_82_0 ;
  wire \i_/bdatw[15]_INST_0_i_82_1 ;
  wire \i_/bdatw[15]_INST_0_i_82_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_46_n_0 ;
  wire [15:0]out;
  wire [10:0]p_0_in2_in;

  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_13 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [0]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[0]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_14 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [0]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[0]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[0]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [0]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [0]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[0]_INST_0_i_6 
       (.I0(\i_/bbus_o[0]_INST_0_i_13_n_0 ),
        .I1(\i_/bbus_o[0]_INST_0_i_14_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_10_1 [0]),
        .I3(gr2_bus1),
        .I4(\bbus_o[0]_INST_0_i_1 ),
        .I5(\i_/bbus_o[0]_INST_0_i_16_n_0 ),
        .O(\grn_reg[4] [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_12 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [1]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[1]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_13 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [1]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[1]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[1]_INST_0_i_15 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [1]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [1]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[1]_INST_0_i_6 
       (.I0(\i_/bbus_o[1]_INST_0_i_12_n_0 ),
        .I1(\i_/bbus_o[1]_INST_0_i_13_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_10_1 [1]),
        .I3(gr2_bus1),
        .I4(\bbus_o[1]_INST_0_i_1 ),
        .I5(\i_/bbus_o[1]_INST_0_i_15_n_0 ),
        .O(\grn_reg[4] [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_13 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [2]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[2]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_14 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [2]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[2]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[2]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [2]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [2]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[2]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[2]_INST_0_i_6 
       (.I0(\i_/bbus_o[2]_INST_0_i_13_n_0 ),
        .I1(\i_/bbus_o[2]_INST_0_i_14_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_10_1 [2]),
        .I3(gr2_bus1),
        .I4(\bbus_o[2]_INST_0_i_1 ),
        .I5(\i_/bbus_o[2]_INST_0_i_16_n_0 ),
        .O(\grn_reg[4] [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_13 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [3]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[3]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_14 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [3]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[3]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[3]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [3]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [3]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[3]_INST_0_i_6 
       (.I0(\i_/bbus_o[3]_INST_0_i_13_n_0 ),
        .I1(\i_/bbus_o[3]_INST_0_i_14_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_10_1 [3]),
        .I3(gr2_bus1),
        .I4(\bbus_o[3]_INST_0_i_1 ),
        .I5(\i_/bbus_o[3]_INST_0_i_16_n_0 ),
        .O(\grn_reg[4] [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_14 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [4]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[4]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_15 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_1 [4]),
        .I3(gr7_bus1),
        .O(\i_/bbus_o[4]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bbus_o[4]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_31_2 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_31_2 [1]),
        .I2(b0bus_sel_0[1]),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[4]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [4]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [4]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[4]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_82_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_82_1 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_28_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_28_1 ),
        .I5(ctl_selb0_0),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_82_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_10_2 ),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_28_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_28_1 ),
        .I5(ctl_selb0_0),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \i_/bbus_o[4]_INST_0_i_6 
       (.I0(\i_/bbus_o[4]_INST_0_i_14_n_0 ),
        .I1(\i_/bbus_o[4]_INST_0_i_15_n_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_10_1 [4]),
        .I3(gr2_bus1),
        .I4(\bbus_o[4]_INST_0_i_1 ),
        .I5(\i_/bbus_o[4]_INST_0_i_18_n_0 ),
        .O(\grn_reg[4] [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [5]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bbus_o[5]_INST_0_i_12 
       (.I0(\i_/bbus_o[5]_INST_0_i_20_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [0]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [5]),
        .O(\i_/bbus_o[5]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [5]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [5]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[5]_INST_0_i_6 
       (.I0(\i_/bbus_o[5]_INST_0_i_11_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[5]_INST_0_i_12_n_0 ),
        .O(p_0_in2_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [6]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bbus_o[6]_INST_0_i_12 
       (.I0(\i_/bbus_o[6]_INST_0_i_20_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [1]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [6]),
        .O(\i_/bbus_o[6]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [6]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [6]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[6]_INST_0_i_6 
       (.I0(\i_/bbus_o[6]_INST_0_i_11_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[6]_INST_0_i_12_n_0 ),
        .O(p_0_in2_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_11 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [7]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bbus_o[7]_INST_0_i_12 
       (.I0(\i_/bbus_o[7]_INST_0_i_20_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [2]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [7]),
        .O(\i_/bbus_o[7]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [7]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [7]),
        .I3(gr3_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bbus_o[7]_INST_0_i_6 
       (.I0(\i_/bbus_o[7]_INST_0_i_11_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bbus_o[7]_INST_0_i_12_n_0 ),
        .O(p_0_in2_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_22 
       (.I0(\i_/bdatw[10]_INST_0_i_47_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [5]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [10]),
        .O(\i_/bdatw[10]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [10]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [10]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[10]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_8 
       (.I0(\i_/bdatw[10]_INST_0_i_21_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_22_n_0 ),
        .O(p_0_in2_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_21 
       (.I0(\i_/bdatw[11]_INST_0_i_47_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [6]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [11]),
        .O(\i_/bdatw[11]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [11]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [11]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[11]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_8 
       (.I0(\i_/bdatw[11]_INST_0_i_20_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_21_n_0 ),
        .O(p_0_in2_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_21 
       (.I0(\i_/bdatw[12]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [7]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [12]),
        .O(\i_/bdatw[12]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [12]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [12]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_8 
       (.I0(\i_/bdatw[12]_INST_0_i_20_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_21_n_0 ),
        .O(p_0_in2_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_21 
       (.I0(\i_/bdatw[13]_INST_0_i_47_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [8]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [13]),
        .O(\i_/bdatw[13]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [13]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [13]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[13]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_8 
       (.I0(\i_/bdatw[13]_INST_0_i_20_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_21_n_0 ),
        .O(p_0_in2_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_22 
       (.I0(\i_/bdatw[14]_INST_0_i_52_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [9]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [14]),
        .O(\i_/bdatw[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [14]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [14]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[14]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_8 
       (.I0(\i_/bdatw[14]_INST_0_i_21_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_22_n_0 ),
        .O(p_0_in2_in[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_10 
       (.I0(\i_/bdatw[15]_INST_0_i_28_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_31_n_0 ),
        .O(p_0_in2_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_82_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_10_6 ),
        .I2(\i_/bdatw[15]_INST_0_i_10_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_28_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_28_1 ),
        .I5(ctl_selb0_0),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/bdatw[15]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_82_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_10_2 ),
        .I2(\i_/bdatw[15]_INST_0_i_28_0 ),
        .I3(\i_/bdatw[15]_INST_0_i_28_1 ),
        .I4(ctl_selb0_0),
        .I5(\i_/bdatw[15]_INST_0_i_10_3 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_82_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [10]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [15]),
        .O(\i_/bdatw[15]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_79 
       (.I0(\i_/bdatw[15]_INST_0_i_82_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_28_3 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_28_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_28_1 ),
        .I5(ctl_selb0_0),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_80 
       (.I0(\i_/bdatw[15]_INST_0_i_82_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_28_2 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_28_0 ),
        .I4(\i_/bdatw[15]_INST_0_i_28_1 ),
        .I5(ctl_selb0_0),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_82 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [15]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [15]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[15]_INST_0_i_82_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/bdatw[15]_INST_0_i_83 
       (.I0(\i_/bdatw[15]_INST_0_i_31_2 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_31_2 [1]),
        .I2(b0bus_sel_0[0]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_21 
       (.I0(\i_/bdatw[8]_INST_0_i_46_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [3]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [8]),
        .O(\i_/bdatw[8]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [8]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [8]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_8 
       (.I0(\i_/bdatw[8]_INST_0_i_20_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_21_n_0 ),
        .O(p_0_in2_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_10_4 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_5 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_21 
       (.I0(\i_/bdatw[9]_INST_0_i_46_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_10_0 [4]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_10_1 [9]),
        .O(\i_/bdatw[9]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_31_0 [9]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_31_1 [9]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[9]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_8 
       (.I0(\i_/bdatw[9]_INST_0_i_20_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_1 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_21_n_0 ),
        .O(p_0_in2_in[4]));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_34
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_14 ,
    \i_/bdatw[15]_INST_0_i_44_0 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_113_0 ,
    \i_/bdatw[15]_INST_0_i_44_1 ,
    \i_/bdatw[15]_INST_0_i_44_2 ,
    \i_/bdatw[15]_INST_0_i_44_3 ,
    \i_/bdatw[15]_INST_0_i_44_4 ,
    \i_/bdatw[15]_INST_0_i_44_5 ,
    \i_/bdatw[15]_INST_0_i_113_1 ,
    \i_/bdatw[15]_INST_0_i_113_2 ,
    bank_sel,
    \i_/bdatw[15]_INST_0_i_112_0 ,
    \i_/bdatw[15]_INST_0_i_112_1 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_112_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_14 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_44_0 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_113_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_44_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_44_2 ;
  input \i_/bdatw[15]_INST_0_i_44_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_44_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_44_5 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_113_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_113_2 ;
  input [0:0]bank_sel;
  input \i_/bdatw[15]_INST_0_i_112_0 ;
  input \i_/bdatw[15]_INST_0_i_112_1 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_112_2 ;

  wire [0:0]bank_sel;
  wire [15:0]\bdatw[15]_INST_0_i_14 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_69_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_59_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_60_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_69_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_78_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_79_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_99_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_112_0 ;
  wire \i_/bdatw[15]_INST_0_i_112_1 ;
  wire \i_/bdatw[15]_INST_0_i_112_2 ;
  wire \i_/bdatw[15]_INST_0_i_112_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_113_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_113_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_113_2 ;
  wire \i_/bdatw[15]_INST_0_i_113_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_130_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_131_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_201_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_216_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_44_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_44_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_44_2 ;
  wire \i_/bdatw[15]_INST_0_i_44_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_44_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_44_5 ;
  wire \i_/bdatw[8]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_70_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_70_n_0 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_13 
       (.I0(\i_/bdatw[10]_INST_0_i_30_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_31_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_52_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_58 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [2]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [2]),
        .I4(\i_/bdatw[10]_INST_0_i_71_n_0 ),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_59 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[10]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_113_2 [2]),
        .I2(bank_sel),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(\i_/bdatw[10]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_13 
       (.I0(\i_/bdatw[11]_INST_0_i_30_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_31_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_52_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_59 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [3]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [3]),
        .I4(\i_/bdatw[11]_INST_0_i_71_n_0 ),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_60 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[11]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_113_2 [3]),
        .I2(bank_sel),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(\i_/bdatw[11]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_13 
       (.I0(\i_/bdatw[12]_INST_0_i_28_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_29_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_50_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_57 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [4]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [4]),
        .I4(\i_/bdatw[12]_INST_0_i_69_n_0 ),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_58 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[12]_INST_0_i_69 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_113_2 [4]),
        .I2(bank_sel),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(\i_/bdatw[12]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_13 
       (.I0(\i_/bdatw[13]_INST_0_i_30_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_31_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_52_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_43 
       (.I0(\i_/bdatw[13]_INST_0_i_59_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_60_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_59_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_60 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_69_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_69 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_13 
       (.I0(\i_/bdatw[14]_INST_0_i_31_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_34_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \i_/bdatw[14]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \i_/bdatw[14]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_44_3 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_34 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_63_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_48 
       (.I0(\i_/bdatw[14]_INST_0_i_78_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_79_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \i_/bdatw[14]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I2(ctl_selb1_rn[2]),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_44_3 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[14]_INST_0_i_58 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_112_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_112_1 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_112_2 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'h00001000)) 
    \i_/bdatw[14]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \i_/bdatw[14]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_44_3 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_78 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_78_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_79 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_99_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_79_n_0 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[14]_INST_0_i_91 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I2(ctl_selb1_rn[0]),
        .I3(ctl_selb1_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000100)) 
    \i_/bdatw[14]_INST_0_i_92 
       (.I0(\i_/bdatw[15]_INST_0_i_44_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_44_0 [0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_99 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_99_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_112 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_112_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_113 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_201_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_113_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_130 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_130_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_131 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_216_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_131_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_201 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_201_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_216 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_216_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_112_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_113_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_130_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_131_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_13 
       (.I0(\i_/bdatw[8]_INST_0_i_29_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_30_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_51_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_58 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [0]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [0]),
        .I4(\i_/bdatw[8]_INST_0_i_70_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_59 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[8]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_113_2 [0]),
        .I2(bank_sel),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(\i_/bdatw[8]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_13 
       (.I0(\i_/bdatw[9]_INST_0_i_29_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_30_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_51_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_113_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_57 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_44_4 [1]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_44_5 [1]),
        .I4(\i_/bdatw[9]_INST_0_i_70_n_0 ),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_58 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_44_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_44_2 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[9]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_113_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_113_2 [1]),
        .I2(bank_sel),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_113_0 ),
        .O(\i_/bdatw[9]_INST_0_i_70_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_35
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_14 ,
    \i_/bdatw[15]_INST_0_i_43_0 ,
    \i_/bdatw[15]_INST_0_i_43_1 ,
    \i_/bdatw[15]_INST_0_i_200_0 ,
    ctl_selb1_rn,
    \i_/bdatw[15]_INST_0_i_200_1 ,
    \i_/bdatw[15]_INST_0_i_111_0 ,
    \i_/bdatw[15]_INST_0_i_43_2 ,
    \i_/bdatw[15]_INST_0_i_43_3 ,
    \i_/bdatw[15]_INST_0_i_110_0 ,
    \i_/bdatw[15]_INST_0_i_110_1 ,
    \i_/bdatw[15]_INST_0_i_110_2 ,
    ctl_selb1_0,
    \i_/bdatw[15]_INST_0_i_110_3 ,
    \i_/bdatw[15]_INST_0_i_111_1 ,
    \i_/bdatw[15]_INST_0_i_111_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_14 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_43_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_43_1 ;
  input [1:0]\i_/bdatw[15]_INST_0_i_200_0 ;
  input [2:0]ctl_selb1_rn;
  input \i_/bdatw[15]_INST_0_i_200_1 ;
  input \i_/bdatw[15]_INST_0_i_111_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_43_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_43_3 ;
  input \i_/bdatw[15]_INST_0_i_110_0 ;
  input \i_/bdatw[15]_INST_0_i_110_1 ;
  input \i_/bdatw[15]_INST_0_i_110_2 ;
  input [0:0]ctl_selb1_0;
  input \i_/bdatw[15]_INST_0_i_110_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_111_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_111_2 ;

  wire [15:0]\bdatw[15]_INST_0_i_14 ;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_72_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_72_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_70_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_61_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_62_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_70_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_100_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_68_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_80_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_81_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_110_0 ;
  wire \i_/bdatw[15]_INST_0_i_110_1 ;
  wire \i_/bdatw[15]_INST_0_i_110_2 ;
  wire \i_/bdatw[15]_INST_0_i_110_3 ;
  wire \i_/bdatw[15]_INST_0_i_110_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_111_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_111_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_111_2 ;
  wire \i_/bdatw[15]_INST_0_i_111_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_132_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_133_n_0 ;
  wire [1:0]\i_/bdatw[15]_INST_0_i_200_0 ;
  wire \i_/bdatw[15]_INST_0_i_200_1 ;
  wire \i_/bdatw[15]_INST_0_i_200_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_217_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_43_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_43_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_43_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_43_3 ;
  wire \i_/bdatw[8]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_71_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_71_n_0 ;
  wire [15:0]out;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_14 
       (.I0(\i_/bdatw[10]_INST_0_i_32_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_33_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [10]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_53_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_61 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [2]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [2]),
        .I4(\i_/bdatw[10]_INST_0_i_72_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_62 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [2]),
        .I3(gr5_bus1),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[10]_INST_0_i_72 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_111_2 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_110_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(\i_/bdatw[10]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_14 
       (.I0(\i_/bdatw[11]_INST_0_i_32_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_33_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [11]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_53_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_62 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [3]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [3]),
        .I4(\i_/bdatw[11]_INST_0_i_72_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_63 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [3]),
        .I3(gr5_bus1),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[11]_INST_0_i_72 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [3]),
        .I1(\i_/bdatw[15]_INST_0_i_111_2 [3]),
        .I2(\i_/bdatw[15]_INST_0_i_110_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(\i_/bdatw[11]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_14 
       (.I0(\i_/bdatw[12]_INST_0_i_30_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_31_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_31 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [12]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_51_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_60 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [4]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [4]),
        .I4(\i_/bdatw[12]_INST_0_i_70_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_61 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [4]),
        .I3(gr5_bus1),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[12]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [4]),
        .I1(\i_/bdatw[15]_INST_0_i_111_2 [4]),
        .I2(\i_/bdatw[15]_INST_0_i_110_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(\i_/bdatw[12]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_14 
       (.I0(\i_/bdatw[13]_INST_0_i_32_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_33_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [13]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_53_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_44 
       (.I0(\i_/bdatw[13]_INST_0_i_61_n_0 ),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [5]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_62_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_61_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_62 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [5]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_70_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_70 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [5]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [5]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_70_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_100 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_14 
       (.I0(\i_/bdatw[14]_INST_0_i_35_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_38_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \i_/bdatw[14]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_200_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_200_0 [1]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \i_/bdatw[14]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_200_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_200_0 [1]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_111_0 ),
        .I5(ctl_selb1_rn[2]),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_38 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [14]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_68_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_49 
       (.I0(\i_/bdatw[14]_INST_0_i_80_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_81_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \i_/bdatw[14]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_200_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_200_0 [1]),
        .I2(ctl_selb1_rn[2]),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_111_0 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \i_/bdatw[14]_INST_0_i_65 
       (.I0(\i_/bdatw[15]_INST_0_i_110_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_110_1 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_110_2 ),
        .I4(ctl_selb1_0),
        .I5(\i_/bdatw[15]_INST_0_i_110_3 ),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'h00004000)) 
    \i_/bdatw[14]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_200_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_200_0 [1]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \i_/bdatw[14]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_200_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_200_0 [1]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_111_0 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_68 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_68_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_80 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_80_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_81 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [6]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_100_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_81_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[14]_INST_0_i_93 
       (.I0(\i_/bdatw[15]_INST_0_i_200_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_200_0 [1]),
        .I2(ctl_selb1_rn[0]),
        .I3(ctl_selb1_rn[1]),
        .I4(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(gr2_bus1));
  LUT5 #(
    .INIT(32'h00000400)) 
    \i_/bdatw[14]_INST_0_i_94 
       (.I0(\i_/bdatw[15]_INST_0_i_200_0 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_200_0 [1]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_110 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_110_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_111 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [15]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_200_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_111_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_132 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_132_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_133 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [7]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_217_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_133_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_200 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_200_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_217 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_217_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_110_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_111_n_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_132_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_133_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_14 
       (.I0(\i_/bdatw[8]_INST_0_i_31_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_32_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [8]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_52_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_61 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [0]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [0]),
        .I4(\i_/bdatw[8]_INST_0_i_71_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_62 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [0]),
        .I3(gr5_bus1),
        .O(\grn_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[8]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [0]),
        .I1(\i_/bdatw[15]_INST_0_i_111_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_110_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(\i_/bdatw[8]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_14 
       (.I0(\i_/bdatw[9]_INST_0_i_31_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_14 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_32_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [9]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_52_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_111_2 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_60 
       (.I0(gr3_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_43_0 [1]),
        .I2(gr4_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_43_1 [1]),
        .I4(\i_/bdatw[9]_INST_0_i_71_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_61 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_14 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_43_2 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_43_3 [1]),
        .I3(gr5_bus1),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/bdatw[9]_INST_0_i_71 
       (.I0(\i_/bdatw[15]_INST_0_i_111_1 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_111_2 [1]),
        .I2(\i_/bdatw[15]_INST_0_i_110_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(\i_/bdatw[15]_INST_0_i_200_1 ),
        .O(\i_/bdatw[9]_INST_0_i_71_n_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_6
   (p_0_in,
    \grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \i_/rgf_c0bus_wb[4]_i_108_0 ,
    \i_/badr[15]_INST_0_i_52_0 ,
    \i_/badr[15]_INST_0_i_52_1 ,
    ctl_sela0_rn,
    ctl_sela0,
    \i_/badr[15]_INST_0_i_52_2 ,
    \i_/rgf_c0bus_wb[4]_i_108_1 ,
    \i_/rgf_c0bus_wb[4]_i_108_2 ,
    \i_/rgf_c0bus_wb[4]_i_108_3 ,
    \i_/rgf_c0bus_wb[4]_i_108_4 ,
    \i_/rgf_c0bus_wb[4]_i_108_5 ,
    \i_/rgf_c0bus_wb[4]_i_108_6 );
  output [15:0]p_0_in;
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\i_/rgf_c0bus_wb[4]_i_108_0 ;
  input \i_/badr[15]_INST_0_i_52_0 ;
  input \i_/badr[15]_INST_0_i_52_1 ;
  input [1:0]ctl_sela0_rn;
  input [0:0]ctl_sela0;
  input \i_/badr[15]_INST_0_i_52_2 ;
  input [15:0]\i_/rgf_c0bus_wb[4]_i_108_1 ;
  input [15:0]\i_/rgf_c0bus_wb[4]_i_108_2 ;
  input [15:0]\i_/rgf_c0bus_wb[4]_i_108_3 ;
  input [15:0]\i_/rgf_c0bus_wb[4]_i_108_4 ;
  input [15:0]\i_/rgf_c0bus_wb[4]_i_108_5 ;
  input [15:0]\i_/rgf_c0bus_wb[4]_i_108_6 ;

  wire [0:0]ctl_sela0;
  wire [1:0]ctl_sela0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_40_n_0 ;
  wire \i_/badr[0]_INST_0_i_41_n_0 ;
  wire \i_/badr[10]_INST_0_i_38_n_0 ;
  wire \i_/badr[10]_INST_0_i_39_n_0 ;
  wire \i_/badr[11]_INST_0_i_43_n_0 ;
  wire \i_/badr[11]_INST_0_i_44_n_0 ;
  wire \i_/badr[12]_INST_0_i_38_n_0 ;
  wire \i_/badr[12]_INST_0_i_39_n_0 ;
  wire \i_/badr[13]_INST_0_i_38_n_0 ;
  wire \i_/badr[13]_INST_0_i_39_n_0 ;
  wire \i_/badr[14]_INST_0_i_38_n_0 ;
  wire \i_/badr[14]_INST_0_i_39_n_0 ;
  wire \i_/badr[15]_INST_0_i_129_n_0 ;
  wire \i_/badr[15]_INST_0_i_132_n_0 ;
  wire \i_/badr[15]_INST_0_i_52_0 ;
  wire \i_/badr[15]_INST_0_i_52_1 ;
  wire \i_/badr[15]_INST_0_i_52_2 ;
  wire \i_/badr[1]_INST_0_i_38_n_0 ;
  wire \i_/badr[1]_INST_0_i_39_n_0 ;
  wire \i_/badr[2]_INST_0_i_38_n_0 ;
  wire \i_/badr[2]_INST_0_i_39_n_0 ;
  wire \i_/badr[3]_INST_0_i_42_n_0 ;
  wire \i_/badr[3]_INST_0_i_43_n_0 ;
  wire \i_/badr[4]_INST_0_i_38_n_0 ;
  wire \i_/badr[4]_INST_0_i_39_n_0 ;
  wire \i_/badr[5]_INST_0_i_38_n_0 ;
  wire \i_/badr[5]_INST_0_i_39_n_0 ;
  wire \i_/badr[6]_INST_0_i_38_n_0 ;
  wire \i_/badr[6]_INST_0_i_39_n_0 ;
  wire \i_/badr[7]_INST_0_i_43_n_0 ;
  wire \i_/badr[7]_INST_0_i_44_n_0 ;
  wire \i_/badr[8]_INST_0_i_38_n_0 ;
  wire \i_/badr[8]_INST_0_i_39_n_0 ;
  wire \i_/badr[9]_INST_0_i_38_n_0 ;
  wire \i_/badr[9]_INST_0_i_39_n_0 ;
  wire \i_/rgf_c0bus_wb[13]_i_38_n_0 ;
  wire \i_/rgf_c0bus_wb[13]_i_39_n_0 ;
  wire \i_/rgf_c0bus_wb[13]_i_40_n_0 ;
  wire \i_/rgf_c0bus_wb[13]_i_41_n_0 ;
  wire \i_/rgf_c0bus_wb[15]_i_33_n_0 ;
  wire \i_/rgf_c0bus_wb[15]_i_34_n_0 ;
  wire [15:0]\i_/rgf_c0bus_wb[4]_i_108_0 ;
  wire [15:0]\i_/rgf_c0bus_wb[4]_i_108_1 ;
  wire [15:0]\i_/rgf_c0bus_wb[4]_i_108_2 ;
  wire [15:0]\i_/rgf_c0bus_wb[4]_i_108_3 ;
  wire [15:0]\i_/rgf_c0bus_wb[4]_i_108_4 ;
  wire [15:0]\i_/rgf_c0bus_wb[4]_i_108_5 ;
  wire [15:0]\i_/rgf_c0bus_wb[4]_i_108_6 ;
  wire \i_/rgf_c0bus_wb[4]_i_109_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_110_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_111_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_112_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_113_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_114_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_115_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_116_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_117_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_118_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_119_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_120_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_121_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_122_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_123_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_124_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_125_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_126_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_127_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_128_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_129_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_130_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_131_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_132_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_133_n_0 ;
  wire \i_/rgf_c0bus_wb[4]_i_134_n_0 ;
  wire [15:0]out;
  wire [15:0]p_0_in;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [0]),
        .I4(\i_/badr[0]_INST_0_i_40_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [0]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [0]),
        .I4(\i_/badr[0]_INST_0_i_41_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_40 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/badr[0]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_41 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [0]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [0]),
        .I3(gr1_bus1),
        .O(\i_/badr[0]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [10]),
        .I4(\i_/badr[10]_INST_0_i_38_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [10]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [10]),
        .I4(\i_/badr[10]_INST_0_i_39_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/badr[10]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [10]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [10]),
        .I3(gr1_bus1),
        .O(\i_/badr[10]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [11]),
        .I4(\i_/badr[11]_INST_0_i_43_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [11]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [11]),
        .I4(\i_/badr[11]_INST_0_i_44_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_43 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/badr[11]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_44 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [11]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [11]),
        .I3(gr1_bus1),
        .O(\i_/badr[11]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [12]),
        .I4(\i_/badr[12]_INST_0_i_38_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [12]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [12]),
        .I4(\i_/badr[12]_INST_0_i_39_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/badr[12]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [12]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [12]),
        .I3(gr1_bus1),
        .O(\i_/badr[12]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [13]),
        .I4(\i_/badr[13]_INST_0_i_38_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [13]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [13]),
        .I4(\i_/badr[13]_INST_0_i_39_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/badr[13]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [13]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [13]),
        .I3(gr1_bus1),
        .O(\i_/badr[13]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [14]),
        .I4(\i_/badr[14]_INST_0_i_38_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [14]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [14]),
        .I4(\i_/badr[14]_INST_0_i_39_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/badr[14]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [14]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [14]),
        .I3(gr1_bus1),
        .O(\i_/badr[14]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \i_/badr[15]_INST_0_i_127 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(\i_/badr[15]_INST_0_i_52_1 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0),
        .I4(\i_/badr[15]_INST_0_i_52_2 ),
        .I5(ctl_sela0_rn[1]),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \i_/badr[15]_INST_0_i_128 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(\i_/badr[15]_INST_0_i_52_1 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_52_2 ),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_129 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/badr[15]_INST_0_i_129_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_130 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(\i_/badr[15]_INST_0_i_52_1 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_52_2 ),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_131 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(\i_/badr[15]_INST_0_i_52_1 ),
        .I2(ctl_sela0_rn[1]),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_52_2 ),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_132 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [15]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [15]),
        .I3(gr1_bus1),
        .O(\i_/badr[15]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_216 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(\i_/badr[15]_INST_0_i_52_1 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_52_2 ),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \i_/badr[15]_INST_0_i_217 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(ctl_sela0_rn[1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\i_/badr[15]_INST_0_i_52_1 ),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_52_2 ),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_218 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\i_/badr[15]_INST_0_i_52_1 ),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_52_2 ),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/badr[15]_INST_0_i_219 
       (.I0(\i_/badr[15]_INST_0_i_52_0 ),
        .I1(\i_/badr[15]_INST_0_i_52_1 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[1]),
        .I4(ctl_sela0),
        .I5(\i_/badr[15]_INST_0_i_52_2 ),
        .O(gr1_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_52 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [15]),
        .I4(\i_/badr[15]_INST_0_i_129_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_53 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [15]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [15]),
        .I4(\i_/badr[15]_INST_0_i_132_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [1]),
        .I4(\i_/badr[1]_INST_0_i_38_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [1]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [1]),
        .I4(\i_/badr[1]_INST_0_i_39_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/badr[1]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [1]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [1]),
        .I3(gr1_bus1),
        .O(\i_/badr[1]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [2]),
        .I4(\i_/badr[2]_INST_0_i_38_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [2]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [2]),
        .I4(\i_/badr[2]_INST_0_i_39_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/badr[2]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [2]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [2]),
        .I3(gr1_bus1),
        .O(\i_/badr[2]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [3]),
        .I4(\i_/badr[3]_INST_0_i_42_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [3]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [3]),
        .I4(\i_/badr[3]_INST_0_i_43_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_42 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/badr[3]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_43 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [3]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [3]),
        .I3(gr1_bus1),
        .O(\i_/badr[3]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [4]),
        .I4(\i_/badr[4]_INST_0_i_38_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [4]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [4]),
        .I4(\i_/badr[4]_INST_0_i_39_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/badr[4]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [4]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [4]),
        .I3(gr1_bus1),
        .O(\i_/badr[4]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [5]),
        .I4(\i_/badr[5]_INST_0_i_38_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [5]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [5]),
        .I4(\i_/badr[5]_INST_0_i_39_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/badr[5]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [5]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [5]),
        .I3(gr1_bus1),
        .O(\i_/badr[5]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [6]),
        .I4(\i_/badr[6]_INST_0_i_38_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [6]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [6]),
        .I4(\i_/badr[6]_INST_0_i_39_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/badr[6]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [6]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [6]),
        .I3(gr1_bus1),
        .O(\i_/badr[6]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_29 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [7]),
        .I4(\i_/badr[7]_INST_0_i_43_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_30 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [7]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [7]),
        .I4(\i_/badr[7]_INST_0_i_44_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_43 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/badr[7]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_44 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [7]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [7]),
        .I3(gr1_bus1),
        .O(\i_/badr[7]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [8]),
        .I4(\i_/badr[8]_INST_0_i_38_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [8]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [8]),
        .I4(\i_/badr[8]_INST_0_i_39_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/badr[8]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [8]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [8]),
        .I3(gr1_bus1),
        .O(\i_/badr[8]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_0 [9]),
        .I4(\i_/badr[9]_INST_0_i_38_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(\i_/rgf_c0bus_wb[4]_i_108_3 [9]),
        .I2(gr4_bus1),
        .I3(\i_/rgf_c0bus_wb[4]_i_108_4 [9]),
        .I4(\i_/badr[9]_INST_0_i_39_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/badr[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_5 [9]),
        .I1(gr2_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_6 [9]),
        .I3(gr1_bus1),
        .O(\i_/badr[9]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[13]_i_36 
       (.I0(\i_/badr[4]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[13]_i_38_n_0 ),
        .I2(\i_/badr[4]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[13]_i_39_n_0 ),
        .O(p_0_in[4]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[13]_i_37 
       (.I0(\i_/badr[0]_INST_0_i_40_n_0 ),
        .I1(\i_/rgf_c0bus_wb[13]_i_40_n_0 ),
        .I2(\i_/badr[0]_INST_0_i_41_n_0 ),
        .I3(\i_/rgf_c0bus_wb[13]_i_41_n_0 ),
        .O(p_0_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[13]_i_38 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [4]),
        .I1(gr0_bus1),
        .I2(out[4]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[13]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[13]_i_39 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [4]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [4]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[13]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[13]_i_40 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [0]),
        .I1(gr0_bus1),
        .I2(out[0]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[13]_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[13]_i_41 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [0]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [0]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[13]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[15]_i_32 
       (.I0(\i_/badr[13]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[15]_i_33_n_0 ),
        .I2(\i_/badr[13]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(p_0_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[15]_i_33 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [13]),
        .I1(gr0_bus1),
        .I2(out[13]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[15]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[15]_i_34 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [13]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [13]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[15]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_101 
       (.I0(\i_/badr[2]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_123_n_0 ),
        .I2(\i_/badr[2]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_124_n_0 ),
        .O(p_0_in[2]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_102 
       (.I0(\i_/badr[7]_INST_0_i_43_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_125_n_0 ),
        .I2(\i_/badr[7]_INST_0_i_44_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_126_n_0 ),
        .O(p_0_in[7]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_103 
       (.I0(\i_/badr[5]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_127_n_0 ),
        .I2(\i_/badr[5]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_128_n_0 ),
        .O(p_0_in[5]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_106 
       (.I0(\i_/badr[11]_INST_0_i_43_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_129_n_0 ),
        .I2(\i_/badr[11]_INST_0_i_44_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_130_n_0 ),
        .O(p_0_in[11]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_107 
       (.I0(\i_/badr[9]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_131_n_0 ),
        .I2(\i_/badr[9]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_132_n_0 ),
        .O(p_0_in[9]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_108 
       (.I0(\i_/badr[15]_INST_0_i_129_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_133_n_0 ),
        .I2(\i_/badr[15]_INST_0_i_132_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_134_n_0 ),
        .O(p_0_in[15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_109 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [1]),
        .I1(gr0_bus1),
        .I2(out[1]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_109_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_110 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [1]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [1]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_110_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_111 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [3]),
        .I1(gr0_bus1),
        .I2(out[3]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_111_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_112 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [3]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [3]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_112_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_113 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [14]),
        .I1(gr0_bus1),
        .I2(out[14]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_113_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_114 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [14]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [14]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_114_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_115 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [10]),
        .I1(gr0_bus1),
        .I2(out[10]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_115_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_116 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [10]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [10]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_116_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_117 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [12]),
        .I1(gr0_bus1),
        .I2(out[12]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_117_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_118 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [12]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [12]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_118_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_119 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [6]),
        .I1(gr0_bus1),
        .I2(out[6]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_119_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_120 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [6]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [6]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_120_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_121 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [8]),
        .I1(gr0_bus1),
        .I2(out[8]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_121_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_122 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [8]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [8]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_122_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_123 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [2]),
        .I1(gr0_bus1),
        .I2(out[2]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_123_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_124 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [2]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [2]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_124_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_125 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [7]),
        .I1(gr0_bus1),
        .I2(out[7]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_125_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_126 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [7]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [7]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_126_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_127 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [5]),
        .I1(gr0_bus1),
        .I2(out[5]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_127_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_128 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [5]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [5]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_128_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_129 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [11]),
        .I1(gr0_bus1),
        .I2(out[11]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_129_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_130 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [11]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [11]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_130_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_131 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [9]),
        .I1(gr0_bus1),
        .I2(out[9]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_131_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_132 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [9]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [9]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_132_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_133 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_0 [15]),
        .I1(gr0_bus1),
        .I2(out[15]),
        .I3(gr7_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_133_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/rgf_c0bus_wb[4]_i_134 
       (.I0(\i_/rgf_c0bus_wb[4]_i_108_4 [15]),
        .I1(gr4_bus1),
        .I2(\i_/rgf_c0bus_wb[4]_i_108_3 [15]),
        .I3(gr3_bus1),
        .O(\i_/rgf_c0bus_wb[4]_i_134_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_66 
       (.I0(\i_/badr[1]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_109_n_0 ),
        .I2(\i_/badr[1]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_110_n_0 ),
        .O(p_0_in[1]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_71 
       (.I0(\i_/badr[3]_INST_0_i_42_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_111_n_0 ),
        .I2(\i_/badr[3]_INST_0_i_43_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_112_n_0 ),
        .O(p_0_in[3]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_78 
       (.I0(\i_/badr[14]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_113_n_0 ),
        .I2(\i_/badr[14]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_114_n_0 ),
        .O(p_0_in[14]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_83 
       (.I0(\i_/badr[10]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_115_n_0 ),
        .I2(\i_/badr[10]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_116_n_0 ),
        .O(p_0_in[10]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_88 
       (.I0(\i_/badr[12]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_117_n_0 ),
        .I2(\i_/badr[12]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_118_n_0 ),
        .O(p_0_in[12]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_93 
       (.I0(\i_/badr[6]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_119_n_0 ),
        .I2(\i_/badr[6]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_120_n_0 ),
        .O(p_0_in[6]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \i_/rgf_c0bus_wb[4]_i_98 
       (.I0(\i_/badr[8]_INST_0_i_38_n_0 ),
        .I1(\i_/rgf_c0bus_wb[4]_i_121_n_0 ),
        .I2(\i_/badr[8]_INST_0_i_39_n_0 ),
        .I3(\i_/rgf_c0bus_wb[4]_i_122_n_0 ),
        .O(p_0_in[8]));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_7
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \sr_reg[1] ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_0 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_0 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_0 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_0 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_0 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_0 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_0 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_0 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_0 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_0 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_0 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_0 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_0 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_0 ,
    \grn_reg[0]_1 ,
    out,
    \rgf_c1bus_wb[4]_i_45 ,
    \badr[15]_INST_0_i_31 ,
    \i_/badr[0]_INST_0_i_18_0 ,
    \i_/badr[0]_INST_0_i_18_1 ,
    \i_/badr[0]_INST_0_i_18_2 ,
    \rgf_c1bus_wb[4]_i_45_0 ,
    \rgf_c1bus_wb[4]_i_40 ,
    \rgf_c1bus_wb[4]_i_40_0 ,
    \rgf_c1bus_wb[4]_i_40_1 ,
    \rgf_c1bus_wb[4]_i_45_1 ,
    \rgf_c1bus_wb[4]_i_42 ,
    \rgf_c1bus_wb[4]_i_42_0 ,
    \rgf_c1bus_wb[4]_i_50 ,
    \rgf_c1bus_wb[4]_i_50_0 ,
    \rgf_c1bus_wb[4]_i_48 ,
    \rgf_c1bus_wb[4]_i_48_0 ,
    \rgf_c1bus_wb[4]_i_64 ,
    \rgf_c1bus_wb[4]_i_64_0 ,
    \rgf_c1bus_wb[4]_i_62 ,
    \rgf_c1bus_wb[4]_i_62_0 ,
    \rgf_c1bus_wb[4]_i_60 ,
    \rgf_c1bus_wb[4]_i_60_0 ,
    \rgf_c1bus_wb[4]_i_58 ,
    \rgf_c1bus_wb[4]_i_58_0 ,
    \rgf_c1bus_wb[4]_i_56 ,
    \rgf_c1bus_wb[4]_i_56_0 ,
    \rgf_c1bus_wb[4]_i_54 ,
    \rgf_c1bus_wb[4]_i_54_0 ,
    \rgf_c1bus_wb[4]_i_52 ,
    \rgf_c1bus_wb[4]_i_52_0 ,
    \rgf_c1bus_wb[4]_i_32 ,
    \rgf_c1bus_wb[4]_i_32_0 ,
    \rgf_c1bus_wb[4]_i_34 ,
    \rgf_c1bus_wb[4]_i_34_0 ,
    \rgf_c1bus_wb[4]_i_36 ,
    \rgf_c1bus_wb[4]_i_36_0 ,
    \rgf_c1bus_wb[4]_i_38 ,
    \rgf_c1bus_wb[4]_i_38_0 ,
    \sr[4]_i_239 ,
    \sr[4]_i_239_0 ,
    a1bus_sel_0,
    \i_/badr[15]_INST_0_i_29_0 ,
    \i_/badr[15]_INST_0_i_29_1 ,
    \i_/badr[0]_INST_0_i_18_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \sr_reg[1] ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\rgf_c1bus_wb[4]_i_45 ;
  input [1:0]\badr[15]_INST_0_i_31 ;
  input \i_/badr[0]_INST_0_i_18_0 ;
  input \i_/badr[0]_INST_0_i_18_1 ;
  input \i_/badr[0]_INST_0_i_18_2 ;
  input [15:0]\rgf_c1bus_wb[4]_i_45_0 ;
  input \rgf_c1bus_wb[4]_i_40 ;
  input \rgf_c1bus_wb[4]_i_40_0 ;
  input [15:0]\rgf_c1bus_wb[4]_i_40_1 ;
  input [15:0]\rgf_c1bus_wb[4]_i_45_1 ;
  input \rgf_c1bus_wb[4]_i_42 ;
  input \rgf_c1bus_wb[4]_i_42_0 ;
  input \rgf_c1bus_wb[4]_i_50 ;
  input \rgf_c1bus_wb[4]_i_50_0 ;
  input \rgf_c1bus_wb[4]_i_48 ;
  input \rgf_c1bus_wb[4]_i_48_0 ;
  input \rgf_c1bus_wb[4]_i_64 ;
  input \rgf_c1bus_wb[4]_i_64_0 ;
  input \rgf_c1bus_wb[4]_i_62 ;
  input \rgf_c1bus_wb[4]_i_62_0 ;
  input \rgf_c1bus_wb[4]_i_60 ;
  input \rgf_c1bus_wb[4]_i_60_0 ;
  input \rgf_c1bus_wb[4]_i_58 ;
  input \rgf_c1bus_wb[4]_i_58_0 ;
  input \rgf_c1bus_wb[4]_i_56 ;
  input \rgf_c1bus_wb[4]_i_56_0 ;
  input \rgf_c1bus_wb[4]_i_54 ;
  input \rgf_c1bus_wb[4]_i_54_0 ;
  input \rgf_c1bus_wb[4]_i_52 ;
  input \rgf_c1bus_wb[4]_i_52_0 ;
  input \rgf_c1bus_wb[4]_i_32 ;
  input \rgf_c1bus_wb[4]_i_32_0 ;
  input \rgf_c1bus_wb[4]_i_34 ;
  input \rgf_c1bus_wb[4]_i_34_0 ;
  input \rgf_c1bus_wb[4]_i_36 ;
  input \rgf_c1bus_wb[4]_i_36_0 ;
  input \rgf_c1bus_wb[4]_i_38 ;
  input \rgf_c1bus_wb[4]_i_38_0 ;
  input \sr[4]_i_239 ;
  input \sr[4]_i_239_0 ;
  input [2:0]a1bus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_29_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_29_1 ;
  input \i_/badr[0]_INST_0_i_18_3 ;

  wire [2:0]a1bus_sel_0;
  wire [1:0]\badr[15]_INST_0_i_31 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \i_/badr[0]_INST_0_i_18_0 ;
  wire \i_/badr[0]_INST_0_i_18_1 ;
  wire \i_/badr[0]_INST_0_i_18_2 ;
  wire \i_/badr[0]_INST_0_i_18_3 ;
  wire \i_/badr[0]_INST_0_i_35_n_0 ;
  wire \i_/badr[10]_INST_0_i_34_n_0 ;
  wire \i_/badr[11]_INST_0_i_35_n_0 ;
  wire \i_/badr[12]_INST_0_i_34_n_0 ;
  wire \i_/badr[13]_INST_0_i_34_n_0 ;
  wire \i_/badr[14]_INST_0_i_34_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_29_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_29_1 ;
  wire \i_/badr[15]_INST_0_i_93_n_0 ;
  wire \i_/badr[1]_INST_0_i_34_n_0 ;
  wire \i_/badr[2]_INST_0_i_34_n_0 ;
  wire \i_/badr[3]_INST_0_i_35_n_0 ;
  wire \i_/badr[4]_INST_0_i_34_n_0 ;
  wire \i_/badr[5]_INST_0_i_34_n_0 ;
  wire \i_/badr[6]_INST_0_i_34_n_0 ;
  wire \i_/badr[7]_INST_0_i_35_n_0 ;
  wire \i_/badr[8]_INST_0_i_34_n_0 ;
  wire \i_/badr[9]_INST_0_i_34_n_0 ;
  wire [15:0]out;
  wire \rgf_c1bus_wb[4]_i_32 ;
  wire \rgf_c1bus_wb[4]_i_32_0 ;
  wire \rgf_c1bus_wb[4]_i_34 ;
  wire \rgf_c1bus_wb[4]_i_34_0 ;
  wire \rgf_c1bus_wb[4]_i_36 ;
  wire \rgf_c1bus_wb[4]_i_36_0 ;
  wire \rgf_c1bus_wb[4]_i_38 ;
  wire \rgf_c1bus_wb[4]_i_38_0 ;
  wire \rgf_c1bus_wb[4]_i_40 ;
  wire \rgf_c1bus_wb[4]_i_40_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_40_1 ;
  wire \rgf_c1bus_wb[4]_i_42 ;
  wire \rgf_c1bus_wb[4]_i_42_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45_1 ;
  wire \rgf_c1bus_wb[4]_i_48 ;
  wire \rgf_c1bus_wb[4]_i_48_0 ;
  wire \rgf_c1bus_wb[4]_i_50 ;
  wire \rgf_c1bus_wb[4]_i_50_0 ;
  wire \rgf_c1bus_wb[4]_i_52 ;
  wire \rgf_c1bus_wb[4]_i_52_0 ;
  wire \rgf_c1bus_wb[4]_i_54 ;
  wire \rgf_c1bus_wb[4]_i_54_0 ;
  wire \rgf_c1bus_wb[4]_i_56 ;
  wire \rgf_c1bus_wb[4]_i_56_0 ;
  wire \rgf_c1bus_wb[4]_i_58 ;
  wire \rgf_c1bus_wb[4]_i_58_0 ;
  wire \rgf_c1bus_wb[4]_i_60 ;
  wire \rgf_c1bus_wb[4]_i_60_0 ;
  wire \rgf_c1bus_wb[4]_i_62 ;
  wire \rgf_c1bus_wb[4]_i_62_0 ;
  wire \rgf_c1bus_wb[4]_i_64 ;
  wire \rgf_c1bus_wb[4]_i_64_0 ;
  wire \sr[4]_i_239 ;
  wire \sr[4]_i_239_0 ;
  wire \sr_reg[1] ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [0]),
        .I4(\i_/badr[0]_INST_0_i_35_n_0 ),
        .O(\grn_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [0]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [0]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [0]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[0]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [10]),
        .I4(\i_/badr[10]_INST_0_i_34_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [10]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [10]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [10]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[10]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [11]),
        .I4(\i_/badr[11]_INST_0_i_35_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [11]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [11]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [11]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[11]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [12]),
        .I4(\i_/badr[12]_INST_0_i_34_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [12]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [12]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [12]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[12]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [13]),
        .I4(\i_/badr[13]_INST_0_i_34_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [13]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [13]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [13]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[13]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [14]),
        .I4(\i_/badr[14]_INST_0_i_34_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [14]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [14]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [14]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[14]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_29 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [15]),
        .I4(\i_/badr[15]_INST_0_i_93_n_0 ),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_30 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [15]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_1 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \i_/badr[15]_INST_0_i_91 
       (.I0(\badr[15]_INST_0_i_31 [1]),
        .I1(\badr[15]_INST_0_i_31 [0]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 ),
        .I4(\i_/badr[0]_INST_0_i_18_2 ),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_92 
       (.I0(\badr[15]_INST_0_i_31 [1]),
        .I1(\badr[15]_INST_0_i_31 [0]),
        .I2(a1bus_sel_0[0]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_93 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [15]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [15]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[15]_INST_0_i_93_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \i_/badr[15]_INST_0_i_94 
       (.I0(\badr[15]_INST_0_i_31 [1]),
        .I1(\badr[15]_INST_0_i_31 [0]),
        .I2(\i_/badr[0]_INST_0_i_18_0 ),
        .I3(\i_/badr[0]_INST_0_i_18_1 ),
        .I4(\i_/badr[0]_INST_0_i_18_2 ),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_95 
       (.I0(\badr[15]_INST_0_i_31 [1]),
        .I1(\badr[15]_INST_0_i_31 [0]),
        .I2(a1bus_sel_0[2]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[15]_INST_0_i_96 
       (.I0(\badr[15]_INST_0_i_31 [1]),
        .I1(\badr[15]_INST_0_i_31 [0]),
        .I2(a1bus_sel_0[1]),
        .O(\sr_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [1]),
        .I4(\i_/badr[1]_INST_0_i_34_n_0 ),
        .O(\grn_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [1]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [1]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[1]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [2]),
        .I4(\i_/badr[2]_INST_0_i_34_n_0 ),
        .O(\grn_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [2]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [2]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[2]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [3]),
        .I4(\i_/badr[3]_INST_0_i_35_n_0 ),
        .O(\grn_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [3]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [3]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [3]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[3]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [4]),
        .I4(\i_/badr[4]_INST_0_i_34_n_0 ),
        .O(\grn_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [4]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [4]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [4]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[4]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [5]),
        .I4(\i_/badr[5]_INST_0_i_34_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [5]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [5]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [5]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[5]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [6]),
        .I4(\i_/badr[6]_INST_0_i_34_n_0 ),
        .O(\grn_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [6]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [6]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [6]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[6]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [7]),
        .I4(\i_/badr[7]_INST_0_i_35_n_0 ),
        .O(\grn_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [7]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [7]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [7]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[7]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [8]),
        .I4(\i_/badr[8]_INST_0_i_34_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [8]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [8]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [8]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[8]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45 [9]),
        .I4(\i_/badr[9]_INST_0_i_34_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_45_1 [9]),
        .I1(gr0_bus1),
        .I2(\rgf_c1bus_wb[4]_i_45_0 [9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_29_0 [9]),
        .I1(\i_/badr[15]_INST_0_i_29_1 [9]),
        .I2(\i_/badr[0]_INST_0_i_18_3 ),
        .I3(\i_/badr[0]_INST_0_i_18_0 ),
        .I4(\i_/badr[0]_INST_0_i_18_1 ),
        .I5(\i_/badr[0]_INST_0_i_18_2 ),
        .O(\i_/badr[9]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_101 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [13]),
        .I2(\rgf_c1bus_wb[4]_i_50 ),
        .I3(\rgf_c1bus_wb[4]_i_50_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [13]),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_105 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [5]),
        .I2(\rgf_c1bus_wb[4]_i_52 ),
        .I3(\rgf_c1bus_wb[4]_i_52_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [5]),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_109 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [6]),
        .I2(\rgf_c1bus_wb[4]_i_54 ),
        .I3(\rgf_c1bus_wb[4]_i_54_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [6]),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_113 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [7]),
        .I2(\rgf_c1bus_wb[4]_i_56 ),
        .I3(\rgf_c1bus_wb[4]_i_56_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [7]),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_117 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [8]),
        .I2(\rgf_c1bus_wb[4]_i_58 ),
        .I3(\rgf_c1bus_wb[4]_i_58_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [8]),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_121 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [9]),
        .I2(\rgf_c1bus_wb[4]_i_60 ),
        .I3(\rgf_c1bus_wb[4]_i_60_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [9]),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_125 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [10]),
        .I2(\rgf_c1bus_wb[4]_i_62 ),
        .I3(\rgf_c1bus_wb[4]_i_62_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [10]),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_129 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [11]),
        .I2(\rgf_c1bus_wb[4]_i_64 ),
        .I3(\rgf_c1bus_wb[4]_i_64_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [11]),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_70 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [4]),
        .I2(\rgf_c1bus_wb[4]_i_32 ),
        .I3(\rgf_c1bus_wb[4]_i_32_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_74 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [3]),
        .I2(\rgf_c1bus_wb[4]_i_34 ),
        .I3(\rgf_c1bus_wb[4]_i_34_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_78 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [2]),
        .I2(\rgf_c1bus_wb[4]_i_36 ),
        .I3(\rgf_c1bus_wb[4]_i_36_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_82 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [1]),
        .I2(\rgf_c1bus_wb[4]_i_38 ),
        .I3(\rgf_c1bus_wb[4]_i_38_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_86 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [15]),
        .I2(\rgf_c1bus_wb[4]_i_40 ),
        .I3(\rgf_c1bus_wb[4]_i_40_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [15]),
        .O(\grn_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_90 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [14]),
        .I2(\rgf_c1bus_wb[4]_i_42 ),
        .I3(\rgf_c1bus_wb[4]_i_42_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [14]),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_97 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [12]),
        .I2(\rgf_c1bus_wb[4]_i_48 ),
        .I3(\rgf_c1bus_wb[4]_i_48_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [12]),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/sr[4]_i_251 
       (.I0(gr7_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_0 [0]),
        .I2(\sr[4]_i_239 ),
        .I3(\sr[4]_i_239_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_40_1 [0]),
        .O(\grn_reg[0]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_8
   (\grn_reg[15] ,
    \sr_reg[1] ,
    \grn_reg[15]_0 ,
    \grn_reg[14] ,
    \grn_reg[14]_0 ,
    \grn_reg[13] ,
    \grn_reg[13]_0 ,
    \grn_reg[12] ,
    \grn_reg[12]_0 ,
    \grn_reg[11] ,
    \grn_reg[11]_0 ,
    \grn_reg[10] ,
    \grn_reg[10]_0 ,
    \grn_reg[9] ,
    \grn_reg[9]_0 ,
    \grn_reg[8] ,
    \grn_reg[8]_0 ,
    \grn_reg[7] ,
    \grn_reg[7]_0 ,
    \grn_reg[6] ,
    \grn_reg[6]_0 ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \grn_reg[4] ,
    \grn_reg[4]_0 ,
    \grn_reg[3] ,
    \grn_reg[3]_0 ,
    \grn_reg[2] ,
    \grn_reg[2]_0 ,
    \grn_reg[1] ,
    \grn_reg[1]_0 ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    out,
    \rgf_c1bus_wb[4]_i_45 ,
    \rgf_c1bus_wb[4]_i_45_0 ,
    \rgf_c1bus_wb[4]_i_45_1 ,
    \badr[15]_INST_0_i_7 ,
    \rgf_c1bus_wb[4]_i_42 ,
    \rgf_c1bus_wb[4]_i_42_0 ,
    \rgf_c1bus_wb[4]_i_50 ,
    \rgf_c1bus_wb[4]_i_50_0 ,
    \rgf_c1bus_wb[4]_i_48 ,
    \rgf_c1bus_wb[4]_i_48_0 ,
    \rgf_c1bus_wb[4]_i_64 ,
    \rgf_c1bus_wb[4]_i_64_0 ,
    \rgf_c1bus_wb[4]_i_62 ,
    \rgf_c1bus_wb[4]_i_62_0 ,
    \rgf_c1bus_wb[4]_i_60 ,
    \rgf_c1bus_wb[4]_i_60_0 ,
    \rgf_c1bus_wb[4]_i_58 ,
    \rgf_c1bus_wb[4]_i_58_0 ,
    \rgf_c1bus_wb[4]_i_56 ,
    \rgf_c1bus_wb[4]_i_56_0 ,
    \rgf_c1bus_wb[4]_i_54 ,
    \rgf_c1bus_wb[4]_i_54_0 ,
    \rgf_c1bus_wb[4]_i_52 ,
    \rgf_c1bus_wb[4]_i_52_0 ,
    \rgf_c1bus_wb[4]_i_32 ,
    \rgf_c1bus_wb[4]_i_32_0 ,
    \rgf_c1bus_wb[4]_i_34 ,
    \rgf_c1bus_wb[4]_i_34_0 ,
    \rgf_c1bus_wb[4]_i_36 ,
    \rgf_c1bus_wb[4]_i_36_0 ,
    \rgf_c1bus_wb[4]_i_38 ,
    \rgf_c1bus_wb[4]_i_38_0 ,
    \rgf_c1bus_wb[4]_i_44 ,
    \rgf_c1bus_wb[4]_i_44_0 ,
    \i_/rgf_c1bus_wb[4]_i_87_0 ,
    \i_/badr[15]_INST_0_i_32_0 ,
    \i_/badr[15]_INST_0_i_32_1 ,
    \i_/badr[15]_INST_0_i_32_2 ,
    a1bus_sel_0,
    \rgf_c1bus_wb[4]_i_45_2 ,
    \rgf_c1bus_wb[4]_i_45_3 ,
    \i_/badr[15]_INST_0_i_32_3 ,
    \i_/badr[15]_INST_0_i_32_4 ,
    \i_/badr[0]_INST_0_i_21_0 );
  output \grn_reg[15] ;
  output \sr_reg[1] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14] ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13] ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12] ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11] ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10] ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9] ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8] ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7] ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6] ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4] ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3] ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2] ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1] ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_1 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input \rgf_c1bus_wb[4]_i_45 ;
  input \rgf_c1bus_wb[4]_i_45_0 ;
  input [15:0]\rgf_c1bus_wb[4]_i_45_1 ;
  input [15:0]\badr[15]_INST_0_i_7 ;
  input \rgf_c1bus_wb[4]_i_42 ;
  input \rgf_c1bus_wb[4]_i_42_0 ;
  input \rgf_c1bus_wb[4]_i_50 ;
  input \rgf_c1bus_wb[4]_i_50_0 ;
  input \rgf_c1bus_wb[4]_i_48 ;
  input \rgf_c1bus_wb[4]_i_48_0 ;
  input \rgf_c1bus_wb[4]_i_64 ;
  input \rgf_c1bus_wb[4]_i_64_0 ;
  input \rgf_c1bus_wb[4]_i_62 ;
  input \rgf_c1bus_wb[4]_i_62_0 ;
  input \rgf_c1bus_wb[4]_i_60 ;
  input \rgf_c1bus_wb[4]_i_60_0 ;
  input \rgf_c1bus_wb[4]_i_58 ;
  input \rgf_c1bus_wb[4]_i_58_0 ;
  input \rgf_c1bus_wb[4]_i_56 ;
  input \rgf_c1bus_wb[4]_i_56_0 ;
  input \rgf_c1bus_wb[4]_i_54 ;
  input \rgf_c1bus_wb[4]_i_54_0 ;
  input \rgf_c1bus_wb[4]_i_52 ;
  input \rgf_c1bus_wb[4]_i_52_0 ;
  input \rgf_c1bus_wb[4]_i_32 ;
  input \rgf_c1bus_wb[4]_i_32_0 ;
  input \rgf_c1bus_wb[4]_i_34 ;
  input \rgf_c1bus_wb[4]_i_34_0 ;
  input \rgf_c1bus_wb[4]_i_36 ;
  input \rgf_c1bus_wb[4]_i_36_0 ;
  input \rgf_c1bus_wb[4]_i_38 ;
  input \rgf_c1bus_wb[4]_i_38_0 ;
  input \rgf_c1bus_wb[4]_i_44 ;
  input \rgf_c1bus_wb[4]_i_44_0 ;
  input [1:0]\i_/rgf_c1bus_wb[4]_i_87_0 ;
  input \i_/badr[15]_INST_0_i_32_0 ;
  input \i_/badr[15]_INST_0_i_32_1 ;
  input \i_/badr[15]_INST_0_i_32_2 ;
  input [2:0]a1bus_sel_0;
  input [15:0]\rgf_c1bus_wb[4]_i_45_2 ;
  input [15:0]\rgf_c1bus_wb[4]_i_45_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_32_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_32_4 ;
  input \i_/badr[0]_INST_0_i_21_0 ;

  wire [2:0]a1bus_sel_0;
  wire [15:0]\badr[15]_INST_0_i_7 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[15]_1 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \i_/badr[0]_INST_0_i_21_0 ;
  wire \i_/badr[0]_INST_0_i_36_n_0 ;
  wire \i_/badr[10]_INST_0_i_35_n_0 ;
  wire \i_/badr[11]_INST_0_i_36_n_0 ;
  wire \i_/badr[12]_INST_0_i_35_n_0 ;
  wire \i_/badr[13]_INST_0_i_35_n_0 ;
  wire \i_/badr[14]_INST_0_i_35_n_0 ;
  wire \i_/badr[15]_INST_0_i_32_0 ;
  wire \i_/badr[15]_INST_0_i_32_1 ;
  wire \i_/badr[15]_INST_0_i_32_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_32_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_32_4 ;
  wire \i_/badr[15]_INST_0_i_99_n_0 ;
  wire \i_/badr[1]_INST_0_i_35_n_0 ;
  wire \i_/badr[2]_INST_0_i_35_n_0 ;
  wire \i_/badr[3]_INST_0_i_36_n_0 ;
  wire \i_/badr[4]_INST_0_i_35_n_0 ;
  wire \i_/badr[5]_INST_0_i_35_n_0 ;
  wire \i_/badr[6]_INST_0_i_35_n_0 ;
  wire \i_/badr[7]_INST_0_i_36_n_0 ;
  wire \i_/badr[8]_INST_0_i_35_n_0 ;
  wire \i_/badr[9]_INST_0_i_35_n_0 ;
  wire [1:0]\i_/rgf_c1bus_wb[4]_i_87_0 ;
  wire [15:0]out;
  wire \rgf_c1bus_wb[4]_i_32 ;
  wire \rgf_c1bus_wb[4]_i_32_0 ;
  wire \rgf_c1bus_wb[4]_i_34 ;
  wire \rgf_c1bus_wb[4]_i_34_0 ;
  wire \rgf_c1bus_wb[4]_i_36 ;
  wire \rgf_c1bus_wb[4]_i_36_0 ;
  wire \rgf_c1bus_wb[4]_i_38 ;
  wire \rgf_c1bus_wb[4]_i_38_0 ;
  wire \rgf_c1bus_wb[4]_i_42 ;
  wire \rgf_c1bus_wb[4]_i_42_0 ;
  wire \rgf_c1bus_wb[4]_i_44 ;
  wire \rgf_c1bus_wb[4]_i_44_0 ;
  wire \rgf_c1bus_wb[4]_i_45 ;
  wire \rgf_c1bus_wb[4]_i_45_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45_1 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45_2 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45_3 ;
  wire \rgf_c1bus_wb[4]_i_48 ;
  wire \rgf_c1bus_wb[4]_i_48_0 ;
  wire \rgf_c1bus_wb[4]_i_50 ;
  wire \rgf_c1bus_wb[4]_i_50_0 ;
  wire \rgf_c1bus_wb[4]_i_52 ;
  wire \rgf_c1bus_wb[4]_i_52_0 ;
  wire \rgf_c1bus_wb[4]_i_54 ;
  wire \rgf_c1bus_wb[4]_i_54_0 ;
  wire \rgf_c1bus_wb[4]_i_56 ;
  wire \rgf_c1bus_wb[4]_i_56_0 ;
  wire \rgf_c1bus_wb[4]_i_58 ;
  wire \rgf_c1bus_wb[4]_i_58_0 ;
  wire \rgf_c1bus_wb[4]_i_60 ;
  wire \rgf_c1bus_wb[4]_i_60_0 ;
  wire \rgf_c1bus_wb[4]_i_62 ;
  wire \rgf_c1bus_wb[4]_i_62_0 ;
  wire \rgf_c1bus_wb[4]_i_64 ;
  wire \rgf_c1bus_wb[4]_i_64_0 ;
  wire \sr_reg[1] ;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [0]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [0]),
        .I4(\i_/badr[0]_INST_0_i_36_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [0]),
        .I1(gr0_bus1),
        .I2(out[0]),
        .I3(gr7_bus1),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[0]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [0]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [0]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[0]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [10]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [10]),
        .I4(\i_/badr[10]_INST_0_i_35_n_0 ),
        .O(\grn_reg[10]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [10]),
        .I1(gr0_bus1),
        .I2(out[10]),
        .I3(gr7_bus1),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[10]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [10]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [10]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[10]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [11]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [11]),
        .I4(\i_/badr[11]_INST_0_i_36_n_0 ),
        .O(\grn_reg[11]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [11]),
        .I1(gr0_bus1),
        .I2(out[11]),
        .I3(gr7_bus1),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[11]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [11]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [11]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[11]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [12]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [12]),
        .I4(\i_/badr[12]_INST_0_i_35_n_0 ),
        .O(\grn_reg[12]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [12]),
        .I1(gr0_bus1),
        .I2(out[12]),
        .I3(gr7_bus1),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[12]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [12]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [12]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[12]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [13]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [13]),
        .I4(\i_/badr[13]_INST_0_i_35_n_0 ),
        .O(\grn_reg[13]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [13]),
        .I1(gr0_bus1),
        .I2(out[13]),
        .I3(gr7_bus1),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[13]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [13]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [13]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[13]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [14]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [14]),
        .I4(\i_/badr[14]_INST_0_i_35_n_0 ),
        .O(\grn_reg[14]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [14]),
        .I1(gr0_bus1),
        .I2(out[14]),
        .I3(gr7_bus1),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[14]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [14]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [14]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[14]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \i_/badr[15]_INST_0_i_100 
       (.I0(\i_/rgf_c1bus_wb[4]_i_87_0 [1]),
        .I1(\i_/rgf_c1bus_wb[4]_i_87_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_32_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_1 ),
        .I4(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[15]_INST_0_i_101 
       (.I0(\i_/rgf_c1bus_wb[4]_i_87_0 [1]),
        .I1(\i_/rgf_c1bus_wb[4]_i_87_0 [0]),
        .I2(a1bus_sel_0[2]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[15]_INST_0_i_102 
       (.I0(\i_/rgf_c1bus_wb[4]_i_87_0 [1]),
        .I1(\i_/rgf_c1bus_wb[4]_i_87_0 [0]),
        .I2(a1bus_sel_0[1]),
        .O(\sr_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_32 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [15]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [15]),
        .I4(\i_/badr[15]_INST_0_i_99_n_0 ),
        .O(\grn_reg[15]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_33 
       (.I0(\badr[15]_INST_0_i_7 [15]),
        .I1(gr0_bus1),
        .I2(out[15]),
        .I3(gr7_bus1),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \i_/badr[15]_INST_0_i_97 
       (.I0(\i_/rgf_c1bus_wb[4]_i_87_0 [1]),
        .I1(\i_/rgf_c1bus_wb[4]_i_87_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_32_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_1 ),
        .I4(\i_/badr[15]_INST_0_i_32_2 ),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[15]_INST_0_i_98 
       (.I0(\i_/rgf_c1bus_wb[4]_i_87_0 [1]),
        .I1(\i_/rgf_c1bus_wb[4]_i_87_0 [0]),
        .I2(a1bus_sel_0[0]),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[15]_INST_0_i_99 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [15]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [15]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[15]_INST_0_i_99_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [1]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [1]),
        .I4(\i_/badr[1]_INST_0_i_35_n_0 ),
        .O(\grn_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [1]),
        .I1(gr0_bus1),
        .I2(out[1]),
        .I3(gr7_bus1),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[1]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [1]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [1]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[1]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [2]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [2]),
        .I4(\i_/badr[2]_INST_0_i_35_n_0 ),
        .O(\grn_reg[2]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [2]),
        .I1(gr0_bus1),
        .I2(out[2]),
        .I3(gr7_bus1),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[2]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [2]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [2]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[2]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [3]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [3]),
        .I4(\i_/badr[3]_INST_0_i_36_n_0 ),
        .O(\grn_reg[3]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [3]),
        .I1(gr0_bus1),
        .I2(out[3]),
        .I3(gr7_bus1),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[3]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [3]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [3]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[3]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [4]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [4]),
        .I4(\i_/badr[4]_INST_0_i_35_n_0 ),
        .O(\grn_reg[4]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [4]),
        .I1(gr0_bus1),
        .I2(out[4]),
        .I3(gr7_bus1),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[4]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [4]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [4]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[4]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [5]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [5]),
        .I4(\i_/badr[5]_INST_0_i_35_n_0 ),
        .O(\grn_reg[5]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [5]),
        .I1(gr0_bus1),
        .I2(out[5]),
        .I3(gr7_bus1),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[5]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [5]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [5]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[5]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [6]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [6]),
        .I4(\i_/badr[6]_INST_0_i_35_n_0 ),
        .O(\grn_reg[6]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [6]),
        .I1(gr0_bus1),
        .I2(out[6]),
        .I3(gr7_bus1),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[6]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [6]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [6]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[6]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [7]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [7]),
        .I4(\i_/badr[7]_INST_0_i_36_n_0 ),
        .O(\grn_reg[7]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [7]),
        .I1(gr0_bus1),
        .I2(out[7]),
        .I3(gr7_bus1),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[7]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [7]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [7]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[7]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [8]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [8]),
        .I4(\i_/badr[8]_INST_0_i_35_n_0 ),
        .O(\grn_reg[8]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [8]),
        .I1(gr0_bus1),
        .I2(out[8]),
        .I3(gr7_bus1),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[8]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [8]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [8]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[8]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_21 
       (.I0(gr3_bus1),
        .I1(\rgf_c1bus_wb[4]_i_45_2 [9]),
        .I2(gr4_bus1),
        .I3(\rgf_c1bus_wb[4]_i_45_3 [9]),
        .I4(\i_/badr[9]_INST_0_i_35_n_0 ),
        .O(\grn_reg[9]_1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_22 
       (.I0(\badr[15]_INST_0_i_7 [9]),
        .I1(gr0_bus1),
        .I2(out[9]),
        .I3(gr7_bus1),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \i_/badr[9]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_32_3 [9]),
        .I1(\i_/badr[15]_INST_0_i_32_4 [9]),
        .I2(\i_/badr[0]_INST_0_i_21_0 ),
        .I3(\i_/badr[15]_INST_0_i_32_0 ),
        .I4(\i_/badr[15]_INST_0_i_32_1 ),
        .I5(\i_/badr[15]_INST_0_i_32_2 ),
        .O(\i_/badr[9]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_102 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(\rgf_c1bus_wb[4]_i_50 ),
        .I3(\rgf_c1bus_wb[4]_i_50_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [13]),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_106 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(\rgf_c1bus_wb[4]_i_52 ),
        .I3(\rgf_c1bus_wb[4]_i_52_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [5]),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_110 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(\rgf_c1bus_wb[4]_i_54 ),
        .I3(\rgf_c1bus_wb[4]_i_54_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [6]),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_114 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(\rgf_c1bus_wb[4]_i_56 ),
        .I3(\rgf_c1bus_wb[4]_i_56_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [7]),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_118 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(\rgf_c1bus_wb[4]_i_58 ),
        .I3(\rgf_c1bus_wb[4]_i_58_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [8]),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_122 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(\rgf_c1bus_wb[4]_i_60 ),
        .I3(\rgf_c1bus_wb[4]_i_60_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [9]),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_126 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(\rgf_c1bus_wb[4]_i_62 ),
        .I3(\rgf_c1bus_wb[4]_i_62_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [10]),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_130 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(\rgf_c1bus_wb[4]_i_64 ),
        .I3(\rgf_c1bus_wb[4]_i_64_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [11]),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_71 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(\rgf_c1bus_wb[4]_i_32 ),
        .I3(\rgf_c1bus_wb[4]_i_32_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_75 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(\rgf_c1bus_wb[4]_i_34 ),
        .I3(\rgf_c1bus_wb[4]_i_34_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_79 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(\rgf_c1bus_wb[4]_i_36 ),
        .I3(\rgf_c1bus_wb[4]_i_36_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_83 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(\rgf_c1bus_wb[4]_i_38 ),
        .I3(\rgf_c1bus_wb[4]_i_38_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_87 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(\rgf_c1bus_wb[4]_i_45 ),
        .I3(\rgf_c1bus_wb[4]_i_45_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [15]),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_91 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(\rgf_c1bus_wb[4]_i_42 ),
        .I3(\rgf_c1bus_wb[4]_i_42_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [14]),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_94 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(\rgf_c1bus_wb[4]_i_44 ),
        .I3(\rgf_c1bus_wb[4]_i_44_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFF8FFF8)) 
    \i_/rgf_c1bus_wb[4]_i_98 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(\rgf_c1bus_wb[4]_i_48 ),
        .I3(\rgf_c1bus_wb[4]_i_48_0 ),
        .I4(\sr_reg[1] ),
        .I5(\rgf_c1bus_wb[4]_i_45_1 [12]),
        .O(\grn_reg[12] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bank_bus" *) 
module mcss_rgf_bank_bus_9
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_11 ,
    \bbus_o[4]_INST_0_i_7 ,
    \bbus_o[4]_INST_0_i_7_0 ,
    \i_/bdatw[15]_INST_0_i_33_0 ,
    \i_/bdatw[15]_INST_0_i_33_1 ,
    \bbus_o[3]_INST_0_i_7 ,
    \bbus_o[3]_INST_0_i_7_0 ,
    \bbus_o[2]_INST_0_i_7 ,
    \bbus_o[2]_INST_0_i_7_0 ,
    \bbus_o[1]_INST_0_i_7 ,
    \bbus_o[1]_INST_0_i_7_0 ,
    \bbus_o[0]_INST_0_i_7 ,
    \bbus_o[0]_INST_0_i_7_0 ,
    \i_/bbus_o[4]_INST_0_i_21_0 ,
    \i_/bdatw[15]_INST_0_i_34_0 ,
    \i_/bbus_o[4]_INST_0_i_20_0 ,
    \i_/bbus_o[4]_INST_0_i_21_1 ,
    \i_/bbus_o[4]_INST_0_i_21_2 ,
    ctl_selb0_0,
    \bdatw[15]_INST_0_i_11_0 ,
    \bdatw[15]_INST_0_i_11_1 ,
    \bbus_o[4]_INST_0_i_7_1 ,
    \bbus_o[4]_INST_0_i_7_2 ,
    \i_/bdatw[15]_INST_0_i_34_1 ,
    \bbus_o[3]_INST_0_i_7_1 ,
    \bbus_o[3]_INST_0_i_7_2 ,
    \bbus_o[2]_INST_0_i_7_1 ,
    \bbus_o[2]_INST_0_i_7_2 ,
    \bbus_o[1]_INST_0_i_7_1 ,
    \bbus_o[1]_INST_0_i_7_2 ,
    \bbus_o[0]_INST_0_i_7_1 ,
    \bbus_o[0]_INST_0_i_7_2 ,
    \i_/bdatw[15]_INST_0_i_34_2 ,
    \i_/bdatw[15]_INST_0_i_92_0 ,
    ctl_selb0_rn,
    \i_/bdatw[15]_INST_0_i_34_3 ,
    b0bus_sel_0,
    \i_/bbus_o[5]_INST_0_i_14_0 ,
    \i_/bbus_o[4]_INST_0_i_20_1 ,
    \i_/bbus_o[4]_INST_0_i_20_2 ,
    \i_/bdatw[15]_INST_0_i_33_2 ,
    \i_/bbus_o[4]_INST_0_i_21_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [10:0]out;
  input [10:0]\bdatw[15]_INST_0_i_11 ;
  input \bbus_o[4]_INST_0_i_7 ;
  input \bbus_o[4]_INST_0_i_7_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_33_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_33_1 ;
  input \bbus_o[3]_INST_0_i_7 ;
  input \bbus_o[3]_INST_0_i_7_0 ;
  input \bbus_o[2]_INST_0_i_7 ;
  input \bbus_o[2]_INST_0_i_7_0 ;
  input \bbus_o[1]_INST_0_i_7 ;
  input \bbus_o[1]_INST_0_i_7_0 ;
  input \bbus_o[0]_INST_0_i_7 ;
  input \bbus_o[0]_INST_0_i_7_0 ;
  input \i_/bbus_o[4]_INST_0_i_21_0 ;
  input \i_/bdatw[15]_INST_0_i_34_0 ;
  input \i_/bbus_o[4]_INST_0_i_20_0 ;
  input \i_/bbus_o[4]_INST_0_i_21_1 ;
  input \i_/bbus_o[4]_INST_0_i_21_2 ;
  input [0:0]ctl_selb0_0;
  input [10:0]\bdatw[15]_INST_0_i_11_0 ;
  input [15:0]\bdatw[15]_INST_0_i_11_1 ;
  input \bbus_o[4]_INST_0_i_7_1 ;
  input \bbus_o[4]_INST_0_i_7_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_34_1 ;
  input \bbus_o[3]_INST_0_i_7_1 ;
  input \bbus_o[3]_INST_0_i_7_2 ;
  input \bbus_o[2]_INST_0_i_7_1 ;
  input \bbus_o[2]_INST_0_i_7_2 ;
  input \bbus_o[1]_INST_0_i_7_1 ;
  input \bbus_o[1]_INST_0_i_7_2 ;
  input \bbus_o[0]_INST_0_i_7_1 ;
  input \bbus_o[0]_INST_0_i_7_2 ;
  input [10:0]\i_/bdatw[15]_INST_0_i_34_2 ;
  input \i_/bdatw[15]_INST_0_i_92_0 ;
  input [1:0]ctl_selb0_rn;
  input \i_/bdatw[15]_INST_0_i_34_3 ;
  input [1:0]b0bus_sel_0;
  input [1:0]\i_/bbus_o[5]_INST_0_i_14_0 ;
  input \i_/bbus_o[4]_INST_0_i_20_1 ;
  input \i_/bbus_o[4]_INST_0_i_20_2 ;
  input \i_/bdatw[15]_INST_0_i_33_2 ;
  input \i_/bbus_o[4]_INST_0_i_21_3 ;

  wire [1:0]b0bus_sel_0;
  wire \bbus_o[0]_INST_0_i_7 ;
  wire \bbus_o[0]_INST_0_i_7_0 ;
  wire \bbus_o[0]_INST_0_i_7_1 ;
  wire \bbus_o[0]_INST_0_i_7_2 ;
  wire \bbus_o[1]_INST_0_i_7 ;
  wire \bbus_o[1]_INST_0_i_7_0 ;
  wire \bbus_o[1]_INST_0_i_7_1 ;
  wire \bbus_o[1]_INST_0_i_7_2 ;
  wire \bbus_o[2]_INST_0_i_7 ;
  wire \bbus_o[2]_INST_0_i_7_0 ;
  wire \bbus_o[2]_INST_0_i_7_1 ;
  wire \bbus_o[2]_INST_0_i_7_2 ;
  wire \bbus_o[3]_INST_0_i_7 ;
  wire \bbus_o[3]_INST_0_i_7_0 ;
  wire \bbus_o[3]_INST_0_i_7_1 ;
  wire \bbus_o[3]_INST_0_i_7_2 ;
  wire \bbus_o[4]_INST_0_i_7 ;
  wire \bbus_o[4]_INST_0_i_7_0 ;
  wire \bbus_o[4]_INST_0_i_7_1 ;
  wire \bbus_o[4]_INST_0_i_7_2 ;
  wire [10:0]\bdatw[15]_INST_0_i_11 ;
  wire [10:0]\bdatw[15]_INST_0_i_11_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_1 ;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/bbus_o[4]_INST_0_i_20_0 ;
  wire \i_/bbus_o[4]_INST_0_i_20_1 ;
  wire \i_/bbus_o[4]_INST_0_i_20_2 ;
  wire \i_/bbus_o[4]_INST_0_i_21_0 ;
  wire \i_/bbus_o[4]_INST_0_i_21_1 ;
  wire \i_/bbus_o[4]_INST_0_i_21_2 ;
  wire \i_/bbus_o[4]_INST_0_i_21_3 ;
  wire [1:0]\i_/bbus_o[5]_INST_0_i_14_0 ;
  wire \i_/bbus_o[5]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[5]_INST_0_i_22_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[6]_INST_0_i_22_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_21_n_0 ;
  wire \i_/bbus_o[7]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_54_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_33_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_33_1 ;
  wire \i_/bdatw[15]_INST_0_i_33_2 ;
  wire \i_/bdatw[15]_INST_0_i_34_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_34_1 ;
  wire [10:0]\i_/bdatw[15]_INST_0_i_34_2 ;
  wire \i_/bdatw[15]_INST_0_i_34_3 ;
  wire \i_/bdatw[15]_INST_0_i_89_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_92_0 ;
  wire \i_/bdatw[15]_INST_0_i_92_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_48_n_0 ;
  wire [10:0]out;

  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[0]_INST_0_i_18 
       (.I0(\bbus_o[0]_INST_0_i_7 ),
        .I1(\bbus_o[0]_INST_0_i_7_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_33_0 [0]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_33_1 [0]),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[0]_INST_0_i_19 
       (.I0(\bbus_o[0]_INST_0_i_7_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [0]),
        .I3(\bbus_o[0]_INST_0_i_7_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_1 [0]),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[1]_INST_0_i_17 
       (.I0(\bbus_o[1]_INST_0_i_7 ),
        .I1(\bbus_o[1]_INST_0_i_7_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_33_0 [1]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_33_1 [1]),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[1]_INST_0_i_18 
       (.I0(\bbus_o[1]_INST_0_i_7_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [1]),
        .I3(\bbus_o[1]_INST_0_i_7_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_1 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[2]_INST_0_i_18 
       (.I0(\bbus_o[2]_INST_0_i_7 ),
        .I1(\bbus_o[2]_INST_0_i_7_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_33_0 [2]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_33_1 [2]),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[2]_INST_0_i_19 
       (.I0(\bbus_o[2]_INST_0_i_7_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [2]),
        .I3(\bbus_o[2]_INST_0_i_7_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_1 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[3]_INST_0_i_18 
       (.I0(\bbus_o[3]_INST_0_i_7 ),
        .I1(\bbus_o[3]_INST_0_i_7_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_33_0 [3]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_33_1 [3]),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[3]_INST_0_i_19 
       (.I0(\bbus_o[3]_INST_0_i_7_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [3]),
        .I3(\bbus_o[3]_INST_0_i_7_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_1 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bbus_o[4]_INST_0_i_20 
       (.I0(\bbus_o[4]_INST_0_i_7 ),
        .I1(\bbus_o[4]_INST_0_i_7_0 ),
        .I2(gr1_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_33_0 [4]),
        .I4(gr2_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_33_1 [4]),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \i_/bbus_o[4]_INST_0_i_21 
       (.I0(\bbus_o[4]_INST_0_i_7_1 ),
        .I1(gr0_bus1),
        .I2(\bdatw[15]_INST_0_i_11_1 [4]),
        .I3(\bbus_o[4]_INST_0_i_7_2 ),
        .I4(gr6_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_34_1 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_33 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bbus_o[4]_INST_0_i_20_1 ),
        .I2(\i_/bbus_o[4]_INST_0_i_20_0 ),
        .I3(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I4(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I5(ctl_selb0_0),
        .O(gr1_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_34 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bbus_o[4]_INST_0_i_20_2 ),
        .I2(\i_/bbus_o[4]_INST_0_i_20_0 ),
        .I3(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I4(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I5(ctl_selb0_0),
        .O(gr2_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bbus_o[4]_INST_0_i_37 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bbus_o[4]_INST_0_i_21_3 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I4(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I5(ctl_selb0_0),
        .O(gr6_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [0]),
        .I4(\i_/bbus_o[5]_INST_0_i_21_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[5]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [0]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [5]),
        .I4(\i_/bbus_o[5]_INST_0_i_22_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bbus_o[5]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [5]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [5]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bbus_o[5]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[5]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[5]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [1]),
        .I4(\i_/bbus_o[6]_INST_0_i_21_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[6]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [1]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [6]),
        .I4(\i_/bbus_o[6]_INST_0_i_22_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bbus_o[6]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [6]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [6]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bbus_o[6]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[6]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[6]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [2]),
        .I4(\i_/bbus_o[7]_INST_0_i_21_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bbus_o[7]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [2]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [7]),
        .I4(\i_/bbus_o[7]_INST_0_i_22_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bbus_o[7]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [7]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [7]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bbus_o[7]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bbus_o[7]_INST_0_i_22 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/bbus_o[7]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [5]),
        .I4(\i_/bdatw[10]_INST_0_i_48_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [5]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_49_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[10]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [10]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [10]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[10]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [6]),
        .I4(\i_/bdatw[11]_INST_0_i_48_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_49_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[11]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [11]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [11]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[11]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [7]),
        .I4(\i_/bdatw[12]_INST_0_i_46_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_47_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[12]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [12]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [12]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[12]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [8]),
        .I4(\i_/bdatw[13]_INST_0_i_48_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_49_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[13]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [13]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [13]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[13]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_24 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [9]),
        .I4(\i_/bdatw[14]_INST_0_i_53_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_54_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[14]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [14]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [14]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[14]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_175 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_92_0 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I4(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I5(ctl_selb0_0),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_33 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [10]),
        .I4(\i_/bdatw[15]_INST_0_i_89_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_92_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_87 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_34_0 ),
        .I2(\i_/bbus_o[4]_INST_0_i_20_0 ),
        .I3(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I4(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I5(ctl_selb0_0),
        .O(gr3_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_88 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_33_2 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I4(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I5(ctl_selb0_0),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[15]_INST_0_i_89 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [15]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [15]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/bdatw[15]_INST_0_i_90 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_34_0 ),
        .I2(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I3(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I4(ctl_selb0_0),
        .I5(\i_/bbus_o[4]_INST_0_i_20_0 ),
        .O(gr7_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_91 
       (.I0(\i_/bbus_o[4]_INST_0_i_21_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_34_3 ),
        .I2(\i_/bbus_o[4]_INST_0_i_20_0 ),
        .I3(\i_/bbus_o[4]_INST_0_i_21_1 ),
        .I4(\i_/bbus_o[4]_INST_0_i_21_2 ),
        .I5(ctl_selb0_0),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_92 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_92_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [3]),
        .I4(\i_/bdatw[8]_INST_0_i_47_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [3]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_48_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[8]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [8]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [8]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[8]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_23 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\bdatw[15]_INST_0_i_11 [4]),
        .I4(\i_/bdatw[9]_INST_0_i_47_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_11_0 [4]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_11_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_48_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT6 #(
    .INIT(64'h00F8000000880000)) 
    \i_/bdatw[9]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_33_1 [9]),
        .I1(b0bus_sel_0[1]),
        .I2(\i_/bdatw[15]_INST_0_i_33_0 [9]),
        .I3(\i_/bbus_o[5]_INST_0_i_14_0 [1]),
        .I4(\i_/bbus_o[5]_INST_0_i_14_0 [0]),
        .I5(b0bus_sel_0[0]),
        .O(\i_/bdatw[9]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_34_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_34_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_48_n_0 ));
endmodule

module mcss_rgf_bus
   (\tr_reg[15] ,
    \sr_reg[15] ,
    \sp_reg[15] ,
    \grn_reg[15] ,
    \tr_reg[14] ,
    \sr_reg[14] ,
    \sp_reg[14] ,
    \grn_reg[14] ,
    \tr_reg[13] ,
    \sr_reg[13] ,
    \sp_reg[13] ,
    \grn_reg[13] ,
    \tr_reg[12] ,
    \sr_reg[12] ,
    \sp_reg[12] ,
    \grn_reg[12] ,
    \tr_reg[11] ,
    \sr_reg[11] ,
    \sp_reg[11] ,
    \grn_reg[11] ,
    \tr_reg[10] ,
    \sr_reg[10] ,
    \sp_reg[10] ,
    \grn_reg[10] ,
    \tr_reg[9] ,
    \sr_reg[9] ,
    \sp_reg[9] ,
    \grn_reg[9] ,
    \tr_reg[8] ,
    \sr_reg[8] ,
    \sp_reg[8] ,
    \grn_reg[8] ,
    \tr_reg[7] ,
    \sr_reg[7] ,
    \sp_reg[7] ,
    \grn_reg[7] ,
    \tr_reg[6] ,
    \sr_reg[6] ,
    \sp_reg[6] ,
    \grn_reg[6] ,
    \tr_reg[5] ,
    \sr_reg[5] ,
    \sp_reg[5] ,
    \grn_reg[5] ,
    \tr_reg[4] ,
    \sr_reg[4] ,
    \sp_reg[4] ,
    \grn_reg[4] ,
    \tr_reg[3] ,
    \sr_reg[3] ,
    \sp_reg[3] ,
    \grn_reg[3] ,
    \tr_reg[2] ,
    \sr_reg[2] ,
    \sp_reg[2] ,
    \grn_reg[2] ,
    \tr_reg[1] ,
    \sr_reg[1] ,
    \sp_reg[1] ,
    \grn_reg[1] ,
    \tr_reg[0] ,
    \sr_reg[0] ,
    \sp_reg[0] ,
    \grn_reg[0] ,
    \sr_reg[15]_0 ,
    \sr_reg[14]_0 ,
    \sr_reg[13]_0 ,
    \sr_reg[12]_0 ,
    \sr_reg[11]_0 ,
    \sr_reg[10]_0 ,
    \sr_reg[9]_0 ,
    \sr_reg[8]_0 ,
    \sr_reg[7]_0 ,
    \sr_reg[6]_0 ,
    \sr_reg[5]_0 ,
    \sr_reg[4]_0 ,
    \sr_reg[3]_0 ,
    \sr_reg[2]_0 ,
    \sr_reg[1]_0 ,
    \sr_reg[0]_0 ,
    \abus_o[15] ,
    p_1_in,
    p_0_in,
    \rgf_c0bus_wb[4]_i_21 ,
    \rgf_c0bus_wb[4]_i_21_0 ,
    \rgf_c0bus_wb[4]_i_21_1 ,
    \rgf_c0bus_wb[4]_i_21_2 ,
    \abus_o[14] ,
    \rgf_c0bus_wb[4]_i_21_3 ,
    \rgf_c0bus_wb[4]_i_21_4 ,
    \rgf_c0bus_wb[4]_i_21_5 ,
    \rgf_c0bus_wb[4]_i_21_6 ,
    \abus_o[13] ,
    \sr[4]_i_226 ,
    \sr[4]_i_226_0 ,
    \sr[4]_i_226_1 ,
    \sr[4]_i_226_2 ,
    \abus_o[12] ,
    \rgf_c0bus_wb[12]_i_23 ,
    \rgf_c0bus_wb[12]_i_23_0 ,
    \rgf_c0bus_wb[12]_i_23_1 ,
    \rgf_c0bus_wb[12]_i_23_2 ,
    \abus_o[11] ,
    \rgf_c0bus_wb[12]_i_23_3 ,
    \rgf_c0bus_wb[12]_i_23_4 ,
    \rgf_c0bus_wb[12]_i_23_5 ,
    \rgf_c0bus_wb[12]_i_23_6 ,
    \abus_o[10] ,
    \rgf_c0bus_wb[12]_i_22 ,
    \rgf_c0bus_wb[12]_i_22_0 ,
    \rgf_c0bus_wb[12]_i_22_1 ,
    \rgf_c0bus_wb[12]_i_22_2 ,
    \abus_o[9] ,
    \rgf_c0bus_wb[12]_i_22_3 ,
    \rgf_c0bus_wb[12]_i_22_4 ,
    \rgf_c0bus_wb[12]_i_22_5 ,
    \rgf_c0bus_wb[12]_i_22_6 ,
    \abus_o[8] ,
    \rgf_c0bus_wb[12]_i_25 ,
    \rgf_c0bus_wb[12]_i_25_0 ,
    \rgf_c0bus_wb[12]_i_25_1 ,
    \rgf_c0bus_wb[12]_i_25_2 ,
    \abus_o[7] ,
    \rgf_c0bus_wb[12]_i_25_3 ,
    \rgf_c0bus_wb[12]_i_25_4 ,
    \rgf_c0bus_wb[12]_i_25_5 ,
    \rgf_c0bus_wb[12]_i_25_6 ,
    \abus_o[6] ,
    \rgf_c0bus_wb[4]_i_25 ,
    \rgf_c0bus_wb[4]_i_25_0 ,
    \rgf_c0bus_wb[4]_i_25_1 ,
    \rgf_c0bus_wb[4]_i_25_2 ,
    \abus_o[5] ,
    \rgf_c0bus_wb[13]_i_31 ,
    \rgf_c0bus_wb[13]_i_31_0 ,
    \rgf_c0bus_wb[13]_i_31_1 ,
    \rgf_c0bus_wb[13]_i_31_2 ,
    \abus_o[4] ,
    \rgf_c0bus_wb[13]_i_31_3 ,
    \rgf_c0bus_wb[13]_i_31_4 ,
    \rgf_c0bus_wb[13]_i_31_5 ,
    \rgf_c0bus_wb[13]_i_31_6 ,
    \abus_o[3] ,
    \rgf_c0bus_wb[13]_i_30 ,
    \rgf_c0bus_wb[13]_i_30_0 ,
    \rgf_c0bus_wb[13]_i_30_1 ,
    \rgf_c0bus_wb[13]_i_30_2 ,
    \abus_o[2] ,
    \rgf_c0bus_wb[13]_i_30_3 ,
    \rgf_c0bus_wb[13]_i_30_4 ,
    \rgf_c0bus_wb[13]_i_30_5 ,
    \rgf_c0bus_wb[13]_i_30_6 ,
    \abus_o[1] ,
    \rgf_c0bus_wb[13]_i_32 ,
    \rgf_c0bus_wb[13]_i_32_0 ,
    \rgf_c0bus_wb[13]_i_32_1 ,
    \rgf_c0bus_wb[13]_i_32_2 ,
    \abus_o[0] ,
    \abus_o[0]_0 ,
    \abus_o[0]_1 ,
    \rgf_c0bus_wb[13]_i_32_3 ,
    \rgf_c0bus_wb[13]_i_32_4 ,
    \rgf_c0bus_wb[13]_i_32_5 ,
    \rgf_c0bus_wb[13]_i_32_6 ,
    \rgf_c0bus_wb[4]_i_21_7 ,
    \rgf_c0bus_wb[4]_i_21_8 ,
    p_0_in_0,
    a0bus_sel_cr,
    out,
    \rgf_c0bus_wb[4]_i_21_9 ,
    \rgf_c0bus_wb[4]_i_21_10 ,
    \sr[4]_i_226_3 ,
    \sr[4]_i_226_4 ,
    \sr[4]_i_226_5 ,
    \sr[4]_i_226_6 ,
    \rgf_c0bus_wb[4]_i_24 ,
    \rgf_c0bus_wb[4]_i_24_0 ,
    \rgf_c0bus_wb[4]_i_24_1 ,
    \rgf_c0bus_wb[4]_i_24_2 ,
    \rgf_c0bus_wb[12]_i_23_7 ,
    \rgf_c0bus_wb[12]_i_23_8 ,
    \rgf_c0bus_wb[12]_i_23_9 ,
    \rgf_c0bus_wb[12]_i_23_10 ,
    \rgf_c0bus_wb[4]_i_23 ,
    \rgf_c0bus_wb[4]_i_23_0 ,
    \rgf_c0bus_wb[4]_i_23_1 ,
    \rgf_c0bus_wb[4]_i_23_2 ,
    \rgf_c0bus_wb[12]_i_22_7 ,
    \rgf_c0bus_wb[12]_i_22_8 ,
    \rgf_c0bus_wb[12]_i_22_9 ,
    \rgf_c0bus_wb[12]_i_22_10 ,
    \rgf_c0bus_wb[4]_i_26 ,
    \rgf_c0bus_wb[4]_i_26_0 ,
    \rgf_c0bus_wb[4]_i_26_1 ,
    \rgf_c0bus_wb[4]_i_26_2 ,
    \rgf_c0bus_wb[12]_i_25_7 ,
    \rgf_c0bus_wb[12]_i_25_8 ,
    \rgf_c0bus_wb[12]_i_25_9 ,
    \rgf_c0bus_wb[12]_i_25_10 ,
    \rgf_c0bus_wb[4]_i_25_3 ,
    \rgf_c0bus_wb[4]_i_25_4 ,
    \rgf_c0bus_wb[4]_i_25_5 ,
    \rgf_c0bus_wb[4]_i_25_6 ,
    \rgf_c0bus_wb[4]_i_29 ,
    \rgf_c0bus_wb[4]_i_29_0 ,
    \rgf_c0bus_wb[4]_i_29_1 ,
    \rgf_c0bus_wb[4]_i_29_2 ,
    \rgf_c0bus_wb[13]_i_31_7 ,
    \rgf_c0bus_wb[13]_i_31_8 ,
    \rgf_c0bus_wb[13]_i_31_9 ,
    \rgf_c0bus_wb[13]_i_31_10 ,
    \rgf_c0bus_wb[4]_i_30 ,
    \rgf_c0bus_wb[4]_i_30_0 ,
    \rgf_c0bus_wb[4]_i_30_1 ,
    \rgf_c0bus_wb[4]_i_30_2 ,
    \rgf_c0bus_wb[13]_i_30_7 ,
    \rgf_c0bus_wb[13]_i_30_8 ,
    \rgf_c0bus_wb[13]_i_30_9 ,
    \rgf_c0bus_wb[13]_i_30_10 ,
    \rgf_c0bus_wb[15]_i_30 ,
    \rgf_c0bus_wb[15]_i_30_0 ,
    \rgf_c0bus_wb[15]_i_30_1 ,
    \rgf_c0bus_wb[15]_i_30_2 ,
    \rgf_c0bus_wb[13]_i_32_7 ,
    \rgf_c0bus_wb[13]_i_32_8 ,
    \rgf_c0bus_wb[13]_i_32_9 ,
    \rgf_c0bus_wb[13]_i_32_10 ,
    \rgf_c0bus_wb[4]_i_20 ,
    \rgf_c0bus_wb[4]_i_20_0 ,
    \rgf_c0bus_wb[4]_i_20_1 ,
    \rgf_c0bus_wb[4]_i_20_2 ,
    O,
    \rgf_c0bus_wb[4]_i_21_11 ,
    \rgf_c0bus_wb[4]_i_21_12 ,
    data3);
  output \tr_reg[15] ;
  output \sr_reg[15] ;
  output \sp_reg[15] ;
  output \grn_reg[15] ;
  output \tr_reg[14] ;
  output \sr_reg[14] ;
  output \sp_reg[14] ;
  output \grn_reg[14] ;
  output \tr_reg[13] ;
  output \sr_reg[13] ;
  output \sp_reg[13] ;
  output \grn_reg[13] ;
  output \tr_reg[12] ;
  output \sr_reg[12] ;
  output \sp_reg[12] ;
  output \grn_reg[12] ;
  output \tr_reg[11] ;
  output \sr_reg[11] ;
  output \sp_reg[11] ;
  output \grn_reg[11] ;
  output \tr_reg[10] ;
  output \sr_reg[10] ;
  output \sp_reg[10] ;
  output \grn_reg[10] ;
  output \tr_reg[9] ;
  output \sr_reg[9] ;
  output \sp_reg[9] ;
  output \grn_reg[9] ;
  output \tr_reg[8] ;
  output \sr_reg[8] ;
  output \sp_reg[8] ;
  output \grn_reg[8] ;
  output \tr_reg[7] ;
  output \sr_reg[7] ;
  output \sp_reg[7] ;
  output \grn_reg[7] ;
  output \tr_reg[6] ;
  output \sr_reg[6] ;
  output \sp_reg[6] ;
  output \grn_reg[6] ;
  output \tr_reg[5] ;
  output \sr_reg[5] ;
  output \sp_reg[5] ;
  output \grn_reg[5] ;
  output \tr_reg[4] ;
  output \sr_reg[4] ;
  output \sp_reg[4] ;
  output \grn_reg[4] ;
  output \tr_reg[3] ;
  output \sr_reg[3] ;
  output \sp_reg[3] ;
  output \grn_reg[3] ;
  output \tr_reg[2] ;
  output \sr_reg[2] ;
  output \sp_reg[2] ;
  output \grn_reg[2] ;
  output \tr_reg[1] ;
  output \sr_reg[1] ;
  output \sp_reg[1] ;
  output \grn_reg[1] ;
  output \tr_reg[0] ;
  output \sr_reg[0] ;
  output \sp_reg[0] ;
  output \grn_reg[0] ;
  output \sr_reg[15]_0 ;
  output \sr_reg[14]_0 ;
  output \sr_reg[13]_0 ;
  output \sr_reg[12]_0 ;
  output \sr_reg[11]_0 ;
  output \sr_reg[10]_0 ;
  output \sr_reg[9]_0 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[4]_0 ;
  output \sr_reg[3]_0 ;
  output \sr_reg[2]_0 ;
  output \sr_reg[1]_0 ;
  output \sr_reg[0]_0 ;
  input \abus_o[15] ;
  input [14:0]p_1_in;
  input [14:0]p_0_in;
  input \rgf_c0bus_wb[4]_i_21 ;
  input \rgf_c0bus_wb[4]_i_21_0 ;
  input \rgf_c0bus_wb[4]_i_21_1 ;
  input \rgf_c0bus_wb[4]_i_21_2 ;
  input \abus_o[14] ;
  input \rgf_c0bus_wb[4]_i_21_3 ;
  input \rgf_c0bus_wb[4]_i_21_4 ;
  input \rgf_c0bus_wb[4]_i_21_5 ;
  input \rgf_c0bus_wb[4]_i_21_6 ;
  input \abus_o[13] ;
  input \sr[4]_i_226 ;
  input \sr[4]_i_226_0 ;
  input \sr[4]_i_226_1 ;
  input \sr[4]_i_226_2 ;
  input \abus_o[12] ;
  input \rgf_c0bus_wb[12]_i_23 ;
  input \rgf_c0bus_wb[12]_i_23_0 ;
  input \rgf_c0bus_wb[12]_i_23_1 ;
  input \rgf_c0bus_wb[12]_i_23_2 ;
  input \abus_o[11] ;
  input \rgf_c0bus_wb[12]_i_23_3 ;
  input \rgf_c0bus_wb[12]_i_23_4 ;
  input \rgf_c0bus_wb[12]_i_23_5 ;
  input \rgf_c0bus_wb[12]_i_23_6 ;
  input \abus_o[10] ;
  input \rgf_c0bus_wb[12]_i_22 ;
  input \rgf_c0bus_wb[12]_i_22_0 ;
  input \rgf_c0bus_wb[12]_i_22_1 ;
  input \rgf_c0bus_wb[12]_i_22_2 ;
  input \abus_o[9] ;
  input \rgf_c0bus_wb[12]_i_22_3 ;
  input \rgf_c0bus_wb[12]_i_22_4 ;
  input \rgf_c0bus_wb[12]_i_22_5 ;
  input \rgf_c0bus_wb[12]_i_22_6 ;
  input \abus_o[8] ;
  input \rgf_c0bus_wb[12]_i_25 ;
  input \rgf_c0bus_wb[12]_i_25_0 ;
  input \rgf_c0bus_wb[12]_i_25_1 ;
  input \rgf_c0bus_wb[12]_i_25_2 ;
  input \abus_o[7] ;
  input \rgf_c0bus_wb[12]_i_25_3 ;
  input \rgf_c0bus_wb[12]_i_25_4 ;
  input \rgf_c0bus_wb[12]_i_25_5 ;
  input \rgf_c0bus_wb[12]_i_25_6 ;
  input \abus_o[6] ;
  input \rgf_c0bus_wb[4]_i_25 ;
  input \rgf_c0bus_wb[4]_i_25_0 ;
  input \rgf_c0bus_wb[4]_i_25_1 ;
  input \rgf_c0bus_wb[4]_i_25_2 ;
  input \abus_o[5] ;
  input \rgf_c0bus_wb[13]_i_31 ;
  input \rgf_c0bus_wb[13]_i_31_0 ;
  input \rgf_c0bus_wb[13]_i_31_1 ;
  input \rgf_c0bus_wb[13]_i_31_2 ;
  input \abus_o[4] ;
  input \rgf_c0bus_wb[13]_i_31_3 ;
  input \rgf_c0bus_wb[13]_i_31_4 ;
  input \rgf_c0bus_wb[13]_i_31_5 ;
  input \rgf_c0bus_wb[13]_i_31_6 ;
  input \abus_o[3] ;
  input \rgf_c0bus_wb[13]_i_30 ;
  input \rgf_c0bus_wb[13]_i_30_0 ;
  input \rgf_c0bus_wb[13]_i_30_1 ;
  input \rgf_c0bus_wb[13]_i_30_2 ;
  input \abus_o[2] ;
  input \rgf_c0bus_wb[13]_i_30_3 ;
  input \rgf_c0bus_wb[13]_i_30_4 ;
  input \rgf_c0bus_wb[13]_i_30_5 ;
  input \rgf_c0bus_wb[13]_i_30_6 ;
  input \abus_o[1] ;
  input \rgf_c0bus_wb[13]_i_32 ;
  input \rgf_c0bus_wb[13]_i_32_0 ;
  input \rgf_c0bus_wb[13]_i_32_1 ;
  input \rgf_c0bus_wb[13]_i_32_2 ;
  input \abus_o[0] ;
  input [0:0]\abus_o[0]_0 ;
  input [0:0]\abus_o[0]_1 ;
  input \rgf_c0bus_wb[13]_i_32_3 ;
  input \rgf_c0bus_wb[13]_i_32_4 ;
  input \rgf_c0bus_wb[13]_i_32_5 ;
  input \rgf_c0bus_wb[13]_i_32_6 ;
  input \rgf_c0bus_wb[4]_i_21_7 ;
  input \rgf_c0bus_wb[4]_i_21_8 ;
  input [15:0]p_0_in_0;
  input [3:0]a0bus_sel_cr;
  input [15:0]out;
  input \rgf_c0bus_wb[4]_i_21_9 ;
  input \rgf_c0bus_wb[4]_i_21_10 ;
  input \sr[4]_i_226_3 ;
  input \sr[4]_i_226_4 ;
  input \sr[4]_i_226_5 ;
  input \sr[4]_i_226_6 ;
  input \rgf_c0bus_wb[4]_i_24 ;
  input \rgf_c0bus_wb[4]_i_24_0 ;
  input \rgf_c0bus_wb[4]_i_24_1 ;
  input \rgf_c0bus_wb[4]_i_24_2 ;
  input \rgf_c0bus_wb[12]_i_23_7 ;
  input \rgf_c0bus_wb[12]_i_23_8 ;
  input \rgf_c0bus_wb[12]_i_23_9 ;
  input \rgf_c0bus_wb[12]_i_23_10 ;
  input \rgf_c0bus_wb[4]_i_23 ;
  input \rgf_c0bus_wb[4]_i_23_0 ;
  input \rgf_c0bus_wb[4]_i_23_1 ;
  input \rgf_c0bus_wb[4]_i_23_2 ;
  input \rgf_c0bus_wb[12]_i_22_7 ;
  input \rgf_c0bus_wb[12]_i_22_8 ;
  input \rgf_c0bus_wb[12]_i_22_9 ;
  input \rgf_c0bus_wb[12]_i_22_10 ;
  input \rgf_c0bus_wb[4]_i_26 ;
  input \rgf_c0bus_wb[4]_i_26_0 ;
  input \rgf_c0bus_wb[4]_i_26_1 ;
  input \rgf_c0bus_wb[4]_i_26_2 ;
  input \rgf_c0bus_wb[12]_i_25_7 ;
  input \rgf_c0bus_wb[12]_i_25_8 ;
  input \rgf_c0bus_wb[12]_i_25_9 ;
  input \rgf_c0bus_wb[12]_i_25_10 ;
  input \rgf_c0bus_wb[4]_i_25_3 ;
  input \rgf_c0bus_wb[4]_i_25_4 ;
  input \rgf_c0bus_wb[4]_i_25_5 ;
  input \rgf_c0bus_wb[4]_i_25_6 ;
  input \rgf_c0bus_wb[4]_i_29 ;
  input \rgf_c0bus_wb[4]_i_29_0 ;
  input \rgf_c0bus_wb[4]_i_29_1 ;
  input \rgf_c0bus_wb[4]_i_29_2 ;
  input \rgf_c0bus_wb[13]_i_31_7 ;
  input \rgf_c0bus_wb[13]_i_31_8 ;
  input \rgf_c0bus_wb[13]_i_31_9 ;
  input \rgf_c0bus_wb[13]_i_31_10 ;
  input \rgf_c0bus_wb[4]_i_30 ;
  input \rgf_c0bus_wb[4]_i_30_0 ;
  input \rgf_c0bus_wb[4]_i_30_1 ;
  input \rgf_c0bus_wb[4]_i_30_2 ;
  input \rgf_c0bus_wb[13]_i_30_7 ;
  input \rgf_c0bus_wb[13]_i_30_8 ;
  input \rgf_c0bus_wb[13]_i_30_9 ;
  input \rgf_c0bus_wb[13]_i_30_10 ;
  input \rgf_c0bus_wb[15]_i_30 ;
  input \rgf_c0bus_wb[15]_i_30_0 ;
  input \rgf_c0bus_wb[15]_i_30_1 ;
  input \rgf_c0bus_wb[15]_i_30_2 ;
  input \rgf_c0bus_wb[13]_i_32_7 ;
  input \rgf_c0bus_wb[13]_i_32_8 ;
  input \rgf_c0bus_wb[13]_i_32_9 ;
  input \rgf_c0bus_wb[13]_i_32_10 ;
  input \rgf_c0bus_wb[4]_i_20 ;
  input \rgf_c0bus_wb[4]_i_20_0 ;
  input \rgf_c0bus_wb[4]_i_20_1 ;
  input \rgf_c0bus_wb[4]_i_20_2 ;
  input [0:0]O;
  input [15:0]\rgf_c0bus_wb[4]_i_21_11 ;
  input [15:0]\rgf_c0bus_wb[4]_i_21_12 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [3:0]a0bus_sel_cr;
  wire \abus_o[0] ;
  wire [0:0]\abus_o[0]_0 ;
  wire [0:0]\abus_o[0]_1 ;
  wire \abus_o[10] ;
  wire \abus_o[11] ;
  wire \abus_o[12] ;
  wire \abus_o[13] ;
  wire \abus_o[14] ;
  wire \abus_o[15] ;
  wire \abus_o[1] ;
  wire \abus_o[2] ;
  wire \abus_o[3] ;
  wire \abus_o[4] ;
  wire \abus_o[5] ;
  wire \abus_o[6] ;
  wire \abus_o[7] ;
  wire \abus_o[8] ;
  wire \abus_o[9] ;
  wire [14:0]data3;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire [15:0]out;
  wire [14:0]p_0_in;
  wire [15:0]p_0_in_0;
  wire [14:0]p_1_in;
  wire \rgf_c0bus_wb[12]_i_22 ;
  wire \rgf_c0bus_wb[12]_i_22_0 ;
  wire \rgf_c0bus_wb[12]_i_22_1 ;
  wire \rgf_c0bus_wb[12]_i_22_10 ;
  wire \rgf_c0bus_wb[12]_i_22_2 ;
  wire \rgf_c0bus_wb[12]_i_22_3 ;
  wire \rgf_c0bus_wb[12]_i_22_4 ;
  wire \rgf_c0bus_wb[12]_i_22_5 ;
  wire \rgf_c0bus_wb[12]_i_22_6 ;
  wire \rgf_c0bus_wb[12]_i_22_7 ;
  wire \rgf_c0bus_wb[12]_i_22_8 ;
  wire \rgf_c0bus_wb[12]_i_22_9 ;
  wire \rgf_c0bus_wb[12]_i_23 ;
  wire \rgf_c0bus_wb[12]_i_23_0 ;
  wire \rgf_c0bus_wb[12]_i_23_1 ;
  wire \rgf_c0bus_wb[12]_i_23_10 ;
  wire \rgf_c0bus_wb[12]_i_23_2 ;
  wire \rgf_c0bus_wb[12]_i_23_3 ;
  wire \rgf_c0bus_wb[12]_i_23_4 ;
  wire \rgf_c0bus_wb[12]_i_23_5 ;
  wire \rgf_c0bus_wb[12]_i_23_6 ;
  wire \rgf_c0bus_wb[12]_i_23_7 ;
  wire \rgf_c0bus_wb[12]_i_23_8 ;
  wire \rgf_c0bus_wb[12]_i_23_9 ;
  wire \rgf_c0bus_wb[12]_i_25 ;
  wire \rgf_c0bus_wb[12]_i_25_0 ;
  wire \rgf_c0bus_wb[12]_i_25_1 ;
  wire \rgf_c0bus_wb[12]_i_25_10 ;
  wire \rgf_c0bus_wb[12]_i_25_2 ;
  wire \rgf_c0bus_wb[12]_i_25_3 ;
  wire \rgf_c0bus_wb[12]_i_25_4 ;
  wire \rgf_c0bus_wb[12]_i_25_5 ;
  wire \rgf_c0bus_wb[12]_i_25_6 ;
  wire \rgf_c0bus_wb[12]_i_25_7 ;
  wire \rgf_c0bus_wb[12]_i_25_8 ;
  wire \rgf_c0bus_wb[12]_i_25_9 ;
  wire \rgf_c0bus_wb[13]_i_30 ;
  wire \rgf_c0bus_wb[13]_i_30_0 ;
  wire \rgf_c0bus_wb[13]_i_30_1 ;
  wire \rgf_c0bus_wb[13]_i_30_10 ;
  wire \rgf_c0bus_wb[13]_i_30_2 ;
  wire \rgf_c0bus_wb[13]_i_30_3 ;
  wire \rgf_c0bus_wb[13]_i_30_4 ;
  wire \rgf_c0bus_wb[13]_i_30_5 ;
  wire \rgf_c0bus_wb[13]_i_30_6 ;
  wire \rgf_c0bus_wb[13]_i_30_7 ;
  wire \rgf_c0bus_wb[13]_i_30_8 ;
  wire \rgf_c0bus_wb[13]_i_30_9 ;
  wire \rgf_c0bus_wb[13]_i_31 ;
  wire \rgf_c0bus_wb[13]_i_31_0 ;
  wire \rgf_c0bus_wb[13]_i_31_1 ;
  wire \rgf_c0bus_wb[13]_i_31_10 ;
  wire \rgf_c0bus_wb[13]_i_31_2 ;
  wire \rgf_c0bus_wb[13]_i_31_3 ;
  wire \rgf_c0bus_wb[13]_i_31_4 ;
  wire \rgf_c0bus_wb[13]_i_31_5 ;
  wire \rgf_c0bus_wb[13]_i_31_6 ;
  wire \rgf_c0bus_wb[13]_i_31_7 ;
  wire \rgf_c0bus_wb[13]_i_31_8 ;
  wire \rgf_c0bus_wb[13]_i_31_9 ;
  wire \rgf_c0bus_wb[13]_i_32 ;
  wire \rgf_c0bus_wb[13]_i_32_0 ;
  wire \rgf_c0bus_wb[13]_i_32_1 ;
  wire \rgf_c0bus_wb[13]_i_32_10 ;
  wire \rgf_c0bus_wb[13]_i_32_2 ;
  wire \rgf_c0bus_wb[13]_i_32_3 ;
  wire \rgf_c0bus_wb[13]_i_32_4 ;
  wire \rgf_c0bus_wb[13]_i_32_5 ;
  wire \rgf_c0bus_wb[13]_i_32_6 ;
  wire \rgf_c0bus_wb[13]_i_32_7 ;
  wire \rgf_c0bus_wb[13]_i_32_8 ;
  wire \rgf_c0bus_wb[13]_i_32_9 ;
  wire \rgf_c0bus_wb[15]_i_30 ;
  wire \rgf_c0bus_wb[15]_i_30_0 ;
  wire \rgf_c0bus_wb[15]_i_30_1 ;
  wire \rgf_c0bus_wb[15]_i_30_2 ;
  wire \rgf_c0bus_wb[4]_i_20 ;
  wire \rgf_c0bus_wb[4]_i_20_0 ;
  wire \rgf_c0bus_wb[4]_i_20_1 ;
  wire \rgf_c0bus_wb[4]_i_20_2 ;
  wire \rgf_c0bus_wb[4]_i_21 ;
  wire \rgf_c0bus_wb[4]_i_21_0 ;
  wire \rgf_c0bus_wb[4]_i_21_1 ;
  wire \rgf_c0bus_wb[4]_i_21_10 ;
  wire [15:0]\rgf_c0bus_wb[4]_i_21_11 ;
  wire [15:0]\rgf_c0bus_wb[4]_i_21_12 ;
  wire \rgf_c0bus_wb[4]_i_21_2 ;
  wire \rgf_c0bus_wb[4]_i_21_3 ;
  wire \rgf_c0bus_wb[4]_i_21_4 ;
  wire \rgf_c0bus_wb[4]_i_21_5 ;
  wire \rgf_c0bus_wb[4]_i_21_6 ;
  wire \rgf_c0bus_wb[4]_i_21_7 ;
  wire \rgf_c0bus_wb[4]_i_21_8 ;
  wire \rgf_c0bus_wb[4]_i_21_9 ;
  wire \rgf_c0bus_wb[4]_i_23 ;
  wire \rgf_c0bus_wb[4]_i_23_0 ;
  wire \rgf_c0bus_wb[4]_i_23_1 ;
  wire \rgf_c0bus_wb[4]_i_23_2 ;
  wire \rgf_c0bus_wb[4]_i_24 ;
  wire \rgf_c0bus_wb[4]_i_24_0 ;
  wire \rgf_c0bus_wb[4]_i_24_1 ;
  wire \rgf_c0bus_wb[4]_i_24_2 ;
  wire \rgf_c0bus_wb[4]_i_25 ;
  wire \rgf_c0bus_wb[4]_i_25_0 ;
  wire \rgf_c0bus_wb[4]_i_25_1 ;
  wire \rgf_c0bus_wb[4]_i_25_2 ;
  wire \rgf_c0bus_wb[4]_i_25_3 ;
  wire \rgf_c0bus_wb[4]_i_25_4 ;
  wire \rgf_c0bus_wb[4]_i_25_5 ;
  wire \rgf_c0bus_wb[4]_i_25_6 ;
  wire \rgf_c0bus_wb[4]_i_26 ;
  wire \rgf_c0bus_wb[4]_i_26_0 ;
  wire \rgf_c0bus_wb[4]_i_26_1 ;
  wire \rgf_c0bus_wb[4]_i_26_2 ;
  wire \rgf_c0bus_wb[4]_i_29 ;
  wire \rgf_c0bus_wb[4]_i_29_0 ;
  wire \rgf_c0bus_wb[4]_i_29_1 ;
  wire \rgf_c0bus_wb[4]_i_29_2 ;
  wire \rgf_c0bus_wb[4]_i_30 ;
  wire \rgf_c0bus_wb[4]_i_30_0 ;
  wire \rgf_c0bus_wb[4]_i_30_1 ;
  wire \rgf_c0bus_wb[4]_i_30_2 ;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[4]_i_226 ;
  wire \sr[4]_i_226_0 ;
  wire \sr[4]_i_226_1 ;
  wire \sr[4]_i_226_2 ;
  wire \sr[4]_i_226_3 ;
  wire \sr[4]_i_226_4 ;
  wire \sr[4]_i_226_5 ;
  wire \sr[4]_i_226_6 ;
  wire \sr_reg[0] ;
  wire \sr_reg[0]_0 ;
  wire \sr_reg[10] ;
  wire \sr_reg[10]_0 ;
  wire \sr_reg[11] ;
  wire \sr_reg[11]_0 ;
  wire \sr_reg[12] ;
  wire \sr_reg[12]_0 ;
  wire \sr_reg[13] ;
  wire \sr_reg[13]_0 ;
  wire \sr_reg[14] ;
  wire \sr_reg[14]_0 ;
  wire \sr_reg[15] ;
  wire \sr_reg[15]_0 ;
  wire \sr_reg[1] ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[2] ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[3] ;
  wire \sr_reg[3]_0 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[9] ;
  wire \sr_reg[9]_0 ;
  wire \tr_reg[0] ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[15] ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[0]_INST_0_i_12 
       (.I0(out[0]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_20_1 ),
        .I3(\rgf_c0bus_wb[4]_i_20_2 ),
        .I4(\rgf_c0bus_wb[4]_i_20_0 ),
        .I5(\rgf_c0bus_wb[4]_i_20 ),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[0]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(O),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [0]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [0]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[0]_INST_0_i_2 
       (.I0(\abus_o[0] ),
        .I1(\abus_o[0]_0 ),
        .I2(\abus_o[0]_1 ),
        .I3(\sr_reg[0] ),
        .I4(\sp_reg[0] ),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[10]_INST_0_i_12 
       (.I0(out[10]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[12]_i_22_9 ),
        .I3(\rgf_c0bus_wb[12]_i_22_10 ),
        .I4(\rgf_c0bus_wb[12]_i_22_8 ),
        .I5(\rgf_c0bus_wb[12]_i_22_7 ),
        .O(\sr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[9]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [10]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [10]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[10]_INST_0_i_2 
       (.I0(\abus_o[10] ),
        .I1(p_1_in[9]),
        .I2(p_0_in[9]),
        .I3(\sr_reg[10] ),
        .I4(\sp_reg[10] ),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[11]_INST_0_i_12 
       (.I0(out[11]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_23_1 ),
        .I3(\rgf_c0bus_wb[4]_i_23_2 ),
        .I4(\rgf_c0bus_wb[4]_i_23_0 ),
        .I5(\rgf_c0bus_wb[4]_i_23 ),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[10]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [11]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [11]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[11]_INST_0_i_2 
       (.I0(\abus_o[11] ),
        .I1(p_1_in[10]),
        .I2(p_0_in[10]),
        .I3(\sr_reg[11] ),
        .I4(\sp_reg[11] ),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[12]_INST_0_i_12 
       (.I0(out[12]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[12]_i_23_9 ),
        .I3(\rgf_c0bus_wb[12]_i_23_10 ),
        .I4(\rgf_c0bus_wb[12]_i_23_8 ),
        .I5(\rgf_c0bus_wb[12]_i_23_7 ),
        .O(\sr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[11]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [12]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [12]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[12]_INST_0_i_2 
       (.I0(\abus_o[12] ),
        .I1(p_1_in[11]),
        .I2(p_0_in[11]),
        .I3(\sr_reg[12] ),
        .I4(\sp_reg[12] ),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[13]_INST_0_i_12 
       (.I0(out[13]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_24_1 ),
        .I3(\rgf_c0bus_wb[4]_i_24_2 ),
        .I4(\rgf_c0bus_wb[4]_i_24_0 ),
        .I5(\rgf_c0bus_wb[4]_i_24 ),
        .O(\sr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[12]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [13]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [13]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[13]_INST_0_i_2 
       (.I0(\abus_o[13] ),
        .I1(p_1_in[12]),
        .I2(p_0_in[12]),
        .I3(\sr_reg[13] ),
        .I4(\sp_reg[13] ),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[14]_INST_0_i_12 
       (.I0(out[14]),
        .I1(a0bus_sel_cr[0]),
        .I2(\sr[4]_i_226_5 ),
        .I3(\sr[4]_i_226_6 ),
        .I4(\sr[4]_i_226_4 ),
        .I5(\sr[4]_i_226_3 ),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[13]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [14]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [14]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[14]_INST_0_i_2 
       (.I0(\abus_o[14] ),
        .I1(p_1_in[13]),
        .I2(p_0_in[13]),
        .I3(\sr_reg[14] ),
        .I4(\sp_reg[14] ),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[15]_INST_0_i_12 
       (.I0(out[15]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_21_9 ),
        .I3(\rgf_c0bus_wb[4]_i_21_10 ),
        .I4(\rgf_c0bus_wb[4]_i_21_8 ),
        .I5(\rgf_c0bus_wb[4]_i_21_7 ),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[14]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [15]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [15]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[15]_INST_0_i_2 
       (.I0(\abus_o[15] ),
        .I1(p_1_in[14]),
        .I2(p_0_in[14]),
        .I3(\sr_reg[15] ),
        .I4(\sp_reg[15] ),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[1]_INST_0_i_12 
       (.I0(out[1]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[13]_i_32_9 ),
        .I3(\rgf_c0bus_wb[13]_i_32_10 ),
        .I4(\rgf_c0bus_wb[13]_i_32_8 ),
        .I5(\rgf_c0bus_wb[13]_i_32_7 ),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[0]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [1]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [1]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[1]_INST_0_i_2 
       (.I0(\abus_o[1] ),
        .I1(p_1_in[0]),
        .I2(p_0_in[0]),
        .I3(\sr_reg[1] ),
        .I4(\sp_reg[1] ),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[2]_INST_0_i_12 
       (.I0(out[2]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[15]_i_30_1 ),
        .I3(\rgf_c0bus_wb[15]_i_30_2 ),
        .I4(\rgf_c0bus_wb[15]_i_30_0 ),
        .I5(\rgf_c0bus_wb[15]_i_30 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[1]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [2]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [2]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[2]_INST_0_i_2 
       (.I0(\abus_o[2] ),
        .I1(p_1_in[1]),
        .I2(p_0_in[1]),
        .I3(\sr_reg[2] ),
        .I4(\sp_reg[2] ),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[3]_INST_0_i_12 
       (.I0(out[3]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[13]_i_30_9 ),
        .I3(\rgf_c0bus_wb[13]_i_30_10 ),
        .I4(\rgf_c0bus_wb[13]_i_30_8 ),
        .I5(\rgf_c0bus_wb[13]_i_30_7 ),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[2]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [3]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [3]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[3]_INST_0_i_2 
       (.I0(\abus_o[3] ),
        .I1(p_1_in[2]),
        .I2(p_0_in[2]),
        .I3(\sr_reg[3] ),
        .I4(\sp_reg[3] ),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[4]_INST_0_i_12 
       (.I0(out[4]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_30_1 ),
        .I3(\rgf_c0bus_wb[4]_i_30_2 ),
        .I4(\rgf_c0bus_wb[4]_i_30_0 ),
        .I5(\rgf_c0bus_wb[4]_i_30 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[3]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [4]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [4]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[4]_INST_0_i_2 
       (.I0(\abus_o[4] ),
        .I1(p_1_in[3]),
        .I2(p_0_in[3]),
        .I3(\sr_reg[4] ),
        .I4(\sp_reg[4] ),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[5]_INST_0_i_12 
       (.I0(out[5]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[13]_i_31_9 ),
        .I3(\rgf_c0bus_wb[13]_i_31_10 ),
        .I4(\rgf_c0bus_wb[13]_i_31_8 ),
        .I5(\rgf_c0bus_wb[13]_i_31_7 ),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[4]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [5]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [5]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[5]_INST_0_i_2 
       (.I0(\abus_o[5] ),
        .I1(p_1_in[4]),
        .I2(p_0_in[4]),
        .I3(\sr_reg[5] ),
        .I4(\sp_reg[5] ),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[6]_INST_0_i_12 
       (.I0(out[6]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_29_1 ),
        .I3(\rgf_c0bus_wb[4]_i_29_2 ),
        .I4(\rgf_c0bus_wb[4]_i_29_0 ),
        .I5(\rgf_c0bus_wb[4]_i_29 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[5]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [6]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [6]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[6]_INST_0_i_2 
       (.I0(\abus_o[6] ),
        .I1(p_1_in[5]),
        .I2(p_0_in[5]),
        .I3(\sr_reg[6] ),
        .I4(\sp_reg[6] ),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[7]_INST_0_i_12 
       (.I0(out[7]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_25_5 ),
        .I3(\rgf_c0bus_wb[4]_i_25_6 ),
        .I4(\rgf_c0bus_wb[4]_i_25_4 ),
        .I5(\rgf_c0bus_wb[4]_i_25_3 ),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[6]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [7]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [7]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[7]_INST_0_i_2 
       (.I0(\abus_o[7] ),
        .I1(p_1_in[6]),
        .I2(p_0_in[6]),
        .I3(\sr_reg[7] ),
        .I4(\sp_reg[7] ),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[8]_INST_0_i_12 
       (.I0(out[8]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[12]_i_25_9 ),
        .I3(\rgf_c0bus_wb[12]_i_25_10 ),
        .I4(\rgf_c0bus_wb[12]_i_25_8 ),
        .I5(\rgf_c0bus_wb[12]_i_25_7 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[7]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [8]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [8]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[8]_INST_0_i_2 
       (.I0(\abus_o[8] ),
        .I1(p_1_in[7]),
        .I2(p_0_in[7]),
        .I3(\sr_reg[8] ),
        .I4(\sp_reg[8] ),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[9]_INST_0_i_12 
       (.I0(out[9]),
        .I1(a0bus_sel_cr[0]),
        .I2(\rgf_c0bus_wb[4]_i_26_1 ),
        .I3(\rgf_c0bus_wb[4]_i_26_2 ),
        .I4(\rgf_c0bus_wb[4]_i_26_0 ),
        .I5(\rgf_c0bus_wb[4]_i_26 ),
        .O(\sr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_13 
       (.I0(a0bus_sel_cr[3]),
        .I1(data3[8]),
        .I2(a0bus_sel_cr[2]),
        .I3(\rgf_c0bus_wb[4]_i_21_11 [9]),
        .I4(\rgf_c0bus_wb[4]_i_21_12 [9]),
        .I5(a0bus_sel_cr[1]),
        .O(\sp_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[9]_INST_0_i_2 
       (.I0(\abus_o[9] ),
        .I1(p_1_in[8]),
        .I2(p_0_in[8]),
        .I3(\sr_reg[9] ),
        .I4(\sp_reg[9] ),
        .O(\tr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[13]_i_34 
       (.I0(\sp_reg[4] ),
        .I1(\rgf_c0bus_wb[4]_i_30 ),
        .I2(\rgf_c0bus_wb[4]_i_30_0 ),
        .I3(p_0_in_0[4]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[4]),
        .O(\sr_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[13]_i_35 
       (.I0(\sp_reg[0] ),
        .I1(\rgf_c0bus_wb[4]_i_20 ),
        .I2(\rgf_c0bus_wb[4]_i_20_0 ),
        .I3(p_0_in_0[0]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[0]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[15]_i_31 
       (.I0(\sp_reg[13] ),
        .I1(\rgf_c0bus_wb[4]_i_24 ),
        .I2(\rgf_c0bus_wb[4]_i_24_0 ),
        .I3(p_0_in_0[13]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[13]),
        .O(\sr_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_35 
       (.I0(\rgf_c0bus_wb[13]_i_30_3 ),
        .I1(\rgf_c0bus_wb[13]_i_30_4 ),
        .I2(\rgf_c0bus_wb[13]_i_30_5 ),
        .I3(\rgf_c0bus_wb[13]_i_30_6 ),
        .I4(\abus_o[2] ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_36 
       (.I0(\sp_reg[1] ),
        .I1(\rgf_c0bus_wb[13]_i_32_7 ),
        .I2(\rgf_c0bus_wb[13]_i_32_8 ),
        .I3(p_0_in_0[1]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[1]),
        .O(\sr_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_37 
       (.I0(\rgf_c0bus_wb[13]_i_32 ),
        .I1(\rgf_c0bus_wb[13]_i_32_0 ),
        .I2(\rgf_c0bus_wb[13]_i_32_1 ),
        .I3(\rgf_c0bus_wb[13]_i_32_2 ),
        .I4(\abus_o[1] ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_38 
       (.I0(\rgf_c0bus_wb[13]_i_31_3 ),
        .I1(\rgf_c0bus_wb[13]_i_31_4 ),
        .I2(\rgf_c0bus_wb[13]_i_31_5 ),
        .I3(\rgf_c0bus_wb[13]_i_31_6 ),
        .I4(\abus_o[4] ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_39 
       (.I0(\sp_reg[3] ),
        .I1(\rgf_c0bus_wb[13]_i_30_7 ),
        .I2(\rgf_c0bus_wb[13]_i_30_8 ),
        .I3(p_0_in_0[3]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[3]),
        .O(\sr_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_40 
       (.I0(\rgf_c0bus_wb[13]_i_30 ),
        .I1(\rgf_c0bus_wb[13]_i_30_0 ),
        .I2(\rgf_c0bus_wb[13]_i_30_1 ),
        .I3(\rgf_c0bus_wb[13]_i_30_2 ),
        .I4(\abus_o[3] ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_41 
       (.I0(\rgf_c0bus_wb[4]_i_21 ),
        .I1(\rgf_c0bus_wb[4]_i_21_0 ),
        .I2(\rgf_c0bus_wb[4]_i_21_1 ),
        .I3(\rgf_c0bus_wb[4]_i_21_2 ),
        .I4(\abus_o[15] ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_42 
       (.I0(\rgf_c0bus_wb[4]_i_21_3 ),
        .I1(\rgf_c0bus_wb[4]_i_21_4 ),
        .I2(\rgf_c0bus_wb[4]_i_21_5 ),
        .I3(\rgf_c0bus_wb[4]_i_21_6 ),
        .I4(\abus_o[14] ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_43 
       (.I0(\sp_reg[14] ),
        .I1(\sr[4]_i_226_3 ),
        .I2(\sr[4]_i_226_4 ),
        .I3(p_0_in_0[14]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[14]),
        .O(\sr_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_44 
       (.I0(\rgf_c0bus_wb[13]_i_32_3 ),
        .I1(\rgf_c0bus_wb[13]_i_32_4 ),
        .I2(\rgf_c0bus_wb[13]_i_32_5 ),
        .I3(\rgf_c0bus_wb[13]_i_32_6 ),
        .I4(\abus_o[0] ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_45 
       (.I0(\rgf_c0bus_wb[12]_i_23_3 ),
        .I1(\rgf_c0bus_wb[12]_i_23_4 ),
        .I2(\rgf_c0bus_wb[12]_i_23_5 ),
        .I3(\rgf_c0bus_wb[12]_i_23_6 ),
        .I4(\abus_o[11] ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_46 
       (.I0(\sp_reg[10] ),
        .I1(\rgf_c0bus_wb[12]_i_22_7 ),
        .I2(\rgf_c0bus_wb[12]_i_22_8 ),
        .I3(p_0_in_0[10]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[10]),
        .O(\sr_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_47 
       (.I0(\rgf_c0bus_wb[12]_i_22 ),
        .I1(\rgf_c0bus_wb[12]_i_22_0 ),
        .I2(\rgf_c0bus_wb[12]_i_22_1 ),
        .I3(\rgf_c0bus_wb[12]_i_22_2 ),
        .I4(\abus_o[10] ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_48 
       (.I0(\sr[4]_i_226 ),
        .I1(\sr[4]_i_226_0 ),
        .I2(\sr[4]_i_226_1 ),
        .I3(\sr[4]_i_226_2 ),
        .I4(\abus_o[13] ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_49 
       (.I0(\sp_reg[12] ),
        .I1(\rgf_c0bus_wb[12]_i_23_7 ),
        .I2(\rgf_c0bus_wb[12]_i_23_8 ),
        .I3(p_0_in_0[12]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[12]),
        .O(\sr_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_50 
       (.I0(\rgf_c0bus_wb[12]_i_23 ),
        .I1(\rgf_c0bus_wb[12]_i_23_0 ),
        .I2(\rgf_c0bus_wb[12]_i_23_1 ),
        .I3(\rgf_c0bus_wb[12]_i_23_2 ),
        .I4(\abus_o[12] ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_51 
       (.I0(\rgf_c0bus_wb[12]_i_25_3 ),
        .I1(\rgf_c0bus_wb[12]_i_25_4 ),
        .I2(\rgf_c0bus_wb[12]_i_25_5 ),
        .I3(\rgf_c0bus_wb[12]_i_25_6 ),
        .I4(\abus_o[7] ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_52 
       (.I0(\sp_reg[6] ),
        .I1(\rgf_c0bus_wb[4]_i_29 ),
        .I2(\rgf_c0bus_wb[4]_i_29_0 ),
        .I3(p_0_in_0[6]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[6]),
        .O(\sr_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_53 
       (.I0(\rgf_c0bus_wb[4]_i_25 ),
        .I1(\rgf_c0bus_wb[4]_i_25_0 ),
        .I2(\rgf_c0bus_wb[4]_i_25_1 ),
        .I3(\rgf_c0bus_wb[4]_i_25_2 ),
        .I4(\abus_o[6] ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_54 
       (.I0(\rgf_c0bus_wb[12]_i_22_3 ),
        .I1(\rgf_c0bus_wb[12]_i_22_4 ),
        .I2(\rgf_c0bus_wb[12]_i_22_5 ),
        .I3(\rgf_c0bus_wb[12]_i_22_6 ),
        .I4(\abus_o[9] ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_55 
       (.I0(\sp_reg[8] ),
        .I1(\rgf_c0bus_wb[12]_i_25_7 ),
        .I2(\rgf_c0bus_wb[12]_i_25_8 ),
        .I3(p_0_in_0[8]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[8]),
        .O(\sr_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_56 
       (.I0(\rgf_c0bus_wb[12]_i_25 ),
        .I1(\rgf_c0bus_wb[12]_i_25_0 ),
        .I2(\rgf_c0bus_wb[12]_i_25_1 ),
        .I3(\rgf_c0bus_wb[12]_i_25_2 ),
        .I4(\abus_o[8] ),
        .O(\grn_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_57 
       (.I0(\sp_reg[2] ),
        .I1(\rgf_c0bus_wb[15]_i_30 ),
        .I2(\rgf_c0bus_wb[15]_i_30_0 ),
        .I3(p_0_in_0[2]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[2]),
        .O(\sr_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_58 
       (.I0(\sp_reg[7] ),
        .I1(\rgf_c0bus_wb[4]_i_25_3 ),
        .I2(\rgf_c0bus_wb[4]_i_25_4 ),
        .I3(p_0_in_0[7]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[7]),
        .O(\sr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_59 
       (.I0(\sp_reg[5] ),
        .I1(\rgf_c0bus_wb[13]_i_31_7 ),
        .I2(\rgf_c0bus_wb[13]_i_31_8 ),
        .I3(p_0_in_0[5]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[5]),
        .O(\sr_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_c0bus_wb[4]_i_60 
       (.I0(\rgf_c0bus_wb[13]_i_31 ),
        .I1(\rgf_c0bus_wb[13]_i_31_0 ),
        .I2(\rgf_c0bus_wb[13]_i_31_1 ),
        .I3(\rgf_c0bus_wb[13]_i_31_2 ),
        .I4(\abus_o[5] ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_61 
       (.I0(\sp_reg[11] ),
        .I1(\rgf_c0bus_wb[4]_i_23 ),
        .I2(\rgf_c0bus_wb[4]_i_23_0 ),
        .I3(p_0_in_0[11]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[11]),
        .O(\sr_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_62 
       (.I0(\sp_reg[9] ),
        .I1(\rgf_c0bus_wb[4]_i_26 ),
        .I2(\rgf_c0bus_wb[4]_i_26_0 ),
        .I3(p_0_in_0[9]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[9]),
        .O(\sr_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf_c0bus_wb[4]_i_63 
       (.I0(\sp_reg[15] ),
        .I1(\rgf_c0bus_wb[4]_i_21_7 ),
        .I2(\rgf_c0bus_wb[4]_i_21_8 ),
        .I3(p_0_in_0[15]),
        .I4(a0bus_sel_cr[0]),
        .I5(out[15]),
        .O(\sr_reg[15]_0 ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_2
   (\tr_reg[15] ,
    \tr_reg[15]_0 ,
    \sp_reg[15] ,
    \grn_reg[15] ,
    \tr_reg[14] ,
    \tr_reg[14]_0 ,
    \grn_reg[14] ,
    \tr_reg[13] ,
    \tr_reg[13]_0 ,
    \grn_reg[13] ,
    \tr_reg[12] ,
    \tr_reg[12]_0 ,
    \grn_reg[12] ,
    \tr_reg[11] ,
    \tr_reg[11]_0 ,
    \grn_reg[11] ,
    \tr_reg[10] ,
    \tr_reg[10]_0 ,
    \grn_reg[10] ,
    \tr_reg[9] ,
    \tr_reg[9]_0 ,
    \grn_reg[9] ,
    \tr_reg[8] ,
    \tr_reg[8]_0 ,
    \tr_reg[7] ,
    \tr_reg[7]_0 ,
    \grn_reg[7] ,
    \tr_reg[6] ,
    \tr_reg[6]_0 ,
    \grn_reg[6] ,
    \tr_reg[5] ,
    \tr_reg[5]_0 ,
    \grn_reg[5] ,
    \tr_reg[4] ,
    \tr_reg[4]_0 ,
    \grn_reg[4] ,
    \tr_reg[3] ,
    \tr_reg[3]_0 ,
    \grn_reg[3] ,
    \tr_reg[2] ,
    \tr_reg[2]_0 ,
    \grn_reg[2] ,
    \tr_reg[1] ,
    \tr_reg[1]_0 ,
    \grn_reg[1] ,
    \tr_reg[0] ,
    \tr_reg[0]_0 ,
    \sp_reg[0] ,
    \grn_reg[0] ,
    \sp_reg[15]_0 ,
    \sr_reg[15] ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[4] ,
    \sp_reg[3] ,
    \sp_reg[2] ,
    \sp_reg[1] ,
    \sp_reg[0]_0 ,
    \sr_reg[0] ,
    p_1_in1_in,
    p_0_in0_in,
    a1bus_sr,
    a1bus_b13,
    \rgf_c1bus_wb[4]_i_23 ,
    \rgf_c1bus_wb[4]_i_23_0 ,
    \rgf_c1bus_wb[4]_i_23_1 ,
    \rgf_c1bus_wb[4]_i_23_2 ,
    \rgf_c1bus_wb[4]_i_23_3 ,
    \rgf_c1bus_wb[4]_i_20 ,
    \rgf_c1bus_wb[4]_i_20_0 ,
    \rgf_c1bus_wb[4]_i_20_1 ,
    \rgf_c1bus_wb[4]_i_20_2 ,
    \rgf_c1bus_wb[4]_i_20_3 ,
    \sr[4]_i_216 ,
    \sr[4]_i_216_0 ,
    \sr[4]_i_216_1 ,
    \sr[4]_i_216_2 ,
    \sr[4]_i_216_3 ,
    \sr[4]_i_207 ,
    \sr[4]_i_207_0 ,
    \sr[4]_i_207_1 ,
    \sr[4]_i_207_2 ,
    \sr[4]_i_207_3 ,
    \sr[4]_i_215 ,
    \sr[4]_i_215_0 ,
    \sr[4]_i_215_1 ,
    \sr[4]_i_215_2 ,
    \sr[4]_i_215_3 ,
    \sr[4]_i_208 ,
    \sr[4]_i_208_0 ,
    \sr[4]_i_208_1 ,
    \sr[4]_i_208_2 ,
    \sr[4]_i_208_3 ,
    \sr[4]_i_218 ,
    \sr[4]_i_218_0 ,
    \sr[4]_i_218_1 ,
    \sr[4]_i_218_2 ,
    \sr[4]_i_218_3 ,
    \sr[4]_i_217 ,
    \sr[4]_i_217_0 ,
    \sr[4]_i_217_1 ,
    \sr[4]_i_217_2 ,
    \sr[4]_i_217_3 ,
    \sr[4]_i_225 ,
    \sr[4]_i_225_0 ,
    \sr[4]_i_225_1 ,
    \sr[4]_i_225_2 ,
    \sr[4]_i_225_3 ,
    \sr[4]_i_219 ,
    \sr[4]_i_219_0 ,
    \sr[4]_i_219_1 ,
    \sr[4]_i_219_2 ,
    \sr[4]_i_219_3 ,
    \sr[4]_i_224 ,
    \sr[4]_i_224_0 ,
    \sr[4]_i_224_1 ,
    \sr[4]_i_224_2 ,
    \sr[4]_i_224_3 ,
    \rgf_c1bus_wb[4]_i_18 ,
    \rgf_c1bus_wb[4]_i_18_0 ,
    \rgf_c1bus_wb[4]_i_18_1 ,
    \rgf_c1bus_wb[4]_i_18_2 ,
    \rgf_c1bus_wb[4]_i_18_3 ,
    \sr[4]_i_220 ,
    \sr[4]_i_220_0 ,
    \sr[4]_i_220_1 ,
    \sr[4]_i_220_2 ,
    \sr[4]_i_220_3 ,
    \rgf_c1bus_wb[4]_i_19 ,
    \rgf_c1bus_wb[4]_i_19_0 ,
    \rgf_c1bus_wb[4]_i_19_1 ,
    \rgf_c1bus_wb[4]_i_19_2 ,
    \rgf_c1bus_wb[4]_i_19_3 ,
    \sr[4]_i_213 ,
    \sr[4]_i_213_0 ,
    \sr[4]_i_213_1 ,
    \sr[4]_i_213_2 ,
    \sr[4]_i_213_3 ,
    \rgf_c1bus_wb[4]_i_22 ,
    \rgf_c1bus_wb[4]_i_20_4 ,
    \rgf_c1bus_wb[4]_i_22_0 ,
    \rgf_c1bus_wb[4]_i_22_1 ,
    \rgf_c1bus_wb[4]_i_22_2 ,
    \rgf_c1bus_wb[4]_i_22_3 ,
    \sr[4]_i_216_4 ,
    \sr[4]_i_216_5 ,
    \sr[4]_i_216_6 ,
    \sr[4]_i_216_7 ,
    \sr[4]_i_216_8 ,
    \sr[4]_i_216_9 ,
    \sr[4]_i_216_10 ,
    \sr[4]_i_216_11 ,
    \sr[4]_i_215_4 ,
    \sr[4]_i_215_5 ,
    \sr[4]_i_215_6 ,
    \sr[4]_i_215_7 ,
    \sr[4]_i_215_8 ,
    \sr[4]_i_215_9 ,
    \sr[4]_i_215_10 ,
    \sr[4]_i_215_11 ,
    \sr[4]_i_218_4 ,
    \sr[4]_i_218_5 ,
    \sr[4]_i_218_6 ,
    \sr[4]_i_218_7 ,
    \sr[4]_i_218_8 ,
    \sr[4]_i_218_9 ,
    \sr[4]_i_218_10 ,
    \sr[4]_i_218_11 ,
    \sr[4]_i_217_4 ,
    \sr[4]_i_217_5 ,
    \sr[4]_i_217_6 ,
    \sr[4]_i_217_7 ,
    \sr[4]_i_225_4 ,
    \sr[4]_i_225_5 ,
    \sr[4]_i_225_6 ,
    \sr[4]_i_225_7 ,
    \sr[4]_i_225_8 ,
    \sr[4]_i_225_9 ,
    \sr[4]_i_225_10 ,
    \sr[4]_i_225_11 ,
    \sr[4]_i_224_4 ,
    \sr[4]_i_224_5 ,
    \sr[4]_i_224_6 ,
    \sr[4]_i_224_7 ,
    \sr[4]_i_224_8 ,
    \sr[4]_i_224_9 ,
    \sr[4]_i_224_10 ,
    \sr[4]_i_224_11 ,
    \rgf_c1bus_wb[4]_i_18_4 ,
    \rgf_c1bus_wb[4]_i_18_5 ,
    \rgf_c1bus_wb[4]_i_18_6 ,
    \rgf_c1bus_wb[4]_i_18_7 ,
    \rgf_c1bus_wb[4]_i_19_4 ,
    \rgf_c1bus_wb[4]_i_19_5 ,
    \rgf_c1bus_wb[4]_i_19_6 ,
    \rgf_c1bus_wb[4]_i_19_7 ,
    \rgf_c1bus_wb[4]_i_19_8 ,
    \rgf_c1bus_wb[4]_i_19_9 ,
    \rgf_c1bus_wb[4]_i_19_10 ,
    \rgf_c1bus_wb[4]_i_19_11 ,
    \rgf_c1bus_wb[4]_i_21 ,
    \sr[4]_i_210 ,
    \rgf_c1bus_wb[4]_i_21_0 ,
    \rgf_c1bus_wb[4]_i_21_1 ,
    \rgf_c1bus_wb[4]_i_21_2 ,
    \rgf_c1bus_wb[4]_i_21_3 ,
    out,
    a1bus_sel_cr,
    \rgf_c1bus_wb[4]_i_22_4 ,
    O,
    \rgf_c1bus_wb[4]_i_22_5 ,
    \rgf_c1bus_wb[4]_i_22_6 ,
    data3);
  output \tr_reg[15] ;
  output \tr_reg[15]_0 ;
  output \sp_reg[15] ;
  output \grn_reg[15] ;
  output \tr_reg[14] ;
  output \tr_reg[14]_0 ;
  output \grn_reg[14] ;
  output \tr_reg[13] ;
  output \tr_reg[13]_0 ;
  output \grn_reg[13] ;
  output \tr_reg[12] ;
  output \tr_reg[12]_0 ;
  output \grn_reg[12] ;
  output \tr_reg[11] ;
  output \tr_reg[11]_0 ;
  output \grn_reg[11] ;
  output \tr_reg[10] ;
  output \tr_reg[10]_0 ;
  output \grn_reg[10] ;
  output \tr_reg[9] ;
  output \tr_reg[9]_0 ;
  output \grn_reg[9] ;
  output \tr_reg[8] ;
  output \tr_reg[8]_0 ;
  output \tr_reg[7] ;
  output \tr_reg[7]_0 ;
  output \grn_reg[7] ;
  output \tr_reg[6] ;
  output \tr_reg[6]_0 ;
  output \grn_reg[6] ;
  output \tr_reg[5] ;
  output \tr_reg[5]_0 ;
  output \grn_reg[5] ;
  output \tr_reg[4] ;
  output \tr_reg[4]_0 ;
  output \grn_reg[4] ;
  output \tr_reg[3] ;
  output \tr_reg[3]_0 ;
  output \grn_reg[3] ;
  output \tr_reg[2] ;
  output \tr_reg[2]_0 ;
  output \grn_reg[2] ;
  output \tr_reg[1] ;
  output \tr_reg[1]_0 ;
  output \grn_reg[1] ;
  output \tr_reg[0] ;
  output \tr_reg[0]_0 ;
  output \sp_reg[0] ;
  output \grn_reg[0] ;
  output \sp_reg[15]_0 ;
  output \sr_reg[15] ;
  output \sp_reg[14] ;
  output \sp_reg[13] ;
  output \sp_reg[12] ;
  output \sp_reg[11] ;
  output \sp_reg[10] ;
  output \sp_reg[9] ;
  output \sp_reg[8] ;
  output \sp_reg[7] ;
  output \sp_reg[6] ;
  output \sp_reg[5] ;
  output \sp_reg[4] ;
  output \sp_reg[3] ;
  output \sp_reg[2] ;
  output \sp_reg[1] ;
  output \sp_reg[0]_0 ;
  output \sr_reg[0] ;
  input [15:0]p_1_in1_in;
  input [15:0]p_0_in0_in;
  input [15:0]a1bus_sr;
  input [15:0]a1bus_b13;
  input \rgf_c1bus_wb[4]_i_23 ;
  input \rgf_c1bus_wb[4]_i_23_0 ;
  input \rgf_c1bus_wb[4]_i_23_1 ;
  input \rgf_c1bus_wb[4]_i_23_2 ;
  input \rgf_c1bus_wb[4]_i_23_3 ;
  input \rgf_c1bus_wb[4]_i_20 ;
  input \rgf_c1bus_wb[4]_i_20_0 ;
  input \rgf_c1bus_wb[4]_i_20_1 ;
  input \rgf_c1bus_wb[4]_i_20_2 ;
  input \rgf_c1bus_wb[4]_i_20_3 ;
  input \sr[4]_i_216 ;
  input \sr[4]_i_216_0 ;
  input \sr[4]_i_216_1 ;
  input \sr[4]_i_216_2 ;
  input \sr[4]_i_216_3 ;
  input \sr[4]_i_207 ;
  input \sr[4]_i_207_0 ;
  input \sr[4]_i_207_1 ;
  input \sr[4]_i_207_2 ;
  input \sr[4]_i_207_3 ;
  input \sr[4]_i_215 ;
  input \sr[4]_i_215_0 ;
  input \sr[4]_i_215_1 ;
  input \sr[4]_i_215_2 ;
  input \sr[4]_i_215_3 ;
  input \sr[4]_i_208 ;
  input \sr[4]_i_208_0 ;
  input \sr[4]_i_208_1 ;
  input \sr[4]_i_208_2 ;
  input \sr[4]_i_208_3 ;
  input \sr[4]_i_218 ;
  input \sr[4]_i_218_0 ;
  input \sr[4]_i_218_1 ;
  input \sr[4]_i_218_2 ;
  input \sr[4]_i_218_3 ;
  input \sr[4]_i_217 ;
  input \sr[4]_i_217_0 ;
  input \sr[4]_i_217_1 ;
  input \sr[4]_i_217_2 ;
  input \sr[4]_i_217_3 ;
  input \sr[4]_i_225 ;
  input \sr[4]_i_225_0 ;
  input \sr[4]_i_225_1 ;
  input \sr[4]_i_225_2 ;
  input \sr[4]_i_225_3 ;
  input \sr[4]_i_219 ;
  input \sr[4]_i_219_0 ;
  input \sr[4]_i_219_1 ;
  input \sr[4]_i_219_2 ;
  input \sr[4]_i_219_3 ;
  input \sr[4]_i_224 ;
  input \sr[4]_i_224_0 ;
  input \sr[4]_i_224_1 ;
  input \sr[4]_i_224_2 ;
  input \sr[4]_i_224_3 ;
  input \rgf_c1bus_wb[4]_i_18 ;
  input \rgf_c1bus_wb[4]_i_18_0 ;
  input \rgf_c1bus_wb[4]_i_18_1 ;
  input \rgf_c1bus_wb[4]_i_18_2 ;
  input \rgf_c1bus_wb[4]_i_18_3 ;
  input \sr[4]_i_220 ;
  input \sr[4]_i_220_0 ;
  input \sr[4]_i_220_1 ;
  input \sr[4]_i_220_2 ;
  input \sr[4]_i_220_3 ;
  input \rgf_c1bus_wb[4]_i_19 ;
  input \rgf_c1bus_wb[4]_i_19_0 ;
  input \rgf_c1bus_wb[4]_i_19_1 ;
  input \rgf_c1bus_wb[4]_i_19_2 ;
  input \rgf_c1bus_wb[4]_i_19_3 ;
  input \sr[4]_i_213 ;
  input \sr[4]_i_213_0 ;
  input \sr[4]_i_213_1 ;
  input \sr[4]_i_213_2 ;
  input \sr[4]_i_213_3 ;
  input \rgf_c1bus_wb[4]_i_22 ;
  input \rgf_c1bus_wb[4]_i_20_4 ;
  input \rgf_c1bus_wb[4]_i_22_0 ;
  input \rgf_c1bus_wb[4]_i_22_1 ;
  input \rgf_c1bus_wb[4]_i_22_2 ;
  input \rgf_c1bus_wb[4]_i_22_3 ;
  input \sr[4]_i_216_4 ;
  input \sr[4]_i_216_5 ;
  input \sr[4]_i_216_6 ;
  input \sr[4]_i_216_7 ;
  input \sr[4]_i_216_8 ;
  input \sr[4]_i_216_9 ;
  input \sr[4]_i_216_10 ;
  input \sr[4]_i_216_11 ;
  input \sr[4]_i_215_4 ;
  input \sr[4]_i_215_5 ;
  input \sr[4]_i_215_6 ;
  input \sr[4]_i_215_7 ;
  input \sr[4]_i_215_8 ;
  input \sr[4]_i_215_9 ;
  input \sr[4]_i_215_10 ;
  input \sr[4]_i_215_11 ;
  input \sr[4]_i_218_4 ;
  input \sr[4]_i_218_5 ;
  input \sr[4]_i_218_6 ;
  input \sr[4]_i_218_7 ;
  input \sr[4]_i_218_8 ;
  input \sr[4]_i_218_9 ;
  input \sr[4]_i_218_10 ;
  input \sr[4]_i_218_11 ;
  input \sr[4]_i_217_4 ;
  input \sr[4]_i_217_5 ;
  input \sr[4]_i_217_6 ;
  input \sr[4]_i_217_7 ;
  input \sr[4]_i_225_4 ;
  input \sr[4]_i_225_5 ;
  input \sr[4]_i_225_6 ;
  input \sr[4]_i_225_7 ;
  input \sr[4]_i_225_8 ;
  input \sr[4]_i_225_9 ;
  input \sr[4]_i_225_10 ;
  input \sr[4]_i_225_11 ;
  input \sr[4]_i_224_4 ;
  input \sr[4]_i_224_5 ;
  input \sr[4]_i_224_6 ;
  input \sr[4]_i_224_7 ;
  input \sr[4]_i_224_8 ;
  input \sr[4]_i_224_9 ;
  input \sr[4]_i_224_10 ;
  input \sr[4]_i_224_11 ;
  input \rgf_c1bus_wb[4]_i_18_4 ;
  input \rgf_c1bus_wb[4]_i_18_5 ;
  input \rgf_c1bus_wb[4]_i_18_6 ;
  input \rgf_c1bus_wb[4]_i_18_7 ;
  input \rgf_c1bus_wb[4]_i_19_4 ;
  input \rgf_c1bus_wb[4]_i_19_5 ;
  input \rgf_c1bus_wb[4]_i_19_6 ;
  input \rgf_c1bus_wb[4]_i_19_7 ;
  input \rgf_c1bus_wb[4]_i_19_8 ;
  input \rgf_c1bus_wb[4]_i_19_9 ;
  input \rgf_c1bus_wb[4]_i_19_10 ;
  input \rgf_c1bus_wb[4]_i_19_11 ;
  input \rgf_c1bus_wb[4]_i_21 ;
  input \sr[4]_i_210 ;
  input \rgf_c1bus_wb[4]_i_21_0 ;
  input \rgf_c1bus_wb[4]_i_21_1 ;
  input \rgf_c1bus_wb[4]_i_21_2 ;
  input \rgf_c1bus_wb[4]_i_21_3 ;
  input [15:0]out;
  input [4:0]a1bus_sel_cr;
  input [15:0]\rgf_c1bus_wb[4]_i_22_4 ;
  input [0:0]O;
  input [15:0]\rgf_c1bus_wb[4]_i_22_5 ;
  input [15:0]\rgf_c1bus_wb[4]_i_22_6 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [15:0]a1bus_b13;
  wire [4:0]a1bus_sel_cr;
  wire [15:0]a1bus_sr;
  wire \badr[10]_INST_0_i_8_n_0 ;
  wire \badr[11]_INST_0_i_8_n_0 ;
  wire \badr[12]_INST_0_i_8_n_0 ;
  wire \badr[13]_INST_0_i_8_n_0 ;
  wire \badr[14]_INST_0_i_8_n_0 ;
  wire \badr[1]_INST_0_i_8_n_0 ;
  wire \badr[2]_INST_0_i_8_n_0 ;
  wire \badr[3]_INST_0_i_8_n_0 ;
  wire \badr[4]_INST_0_i_8_n_0 ;
  wire \badr[5]_INST_0_i_8_n_0 ;
  wire \badr[6]_INST_0_i_8_n_0 ;
  wire \badr[7]_INST_0_i_8_n_0 ;
  wire \badr[8]_INST_0_i_8_n_0 ;
  wire \badr[9]_INST_0_i_8_n_0 ;
  wire [14:0]data3;
  wire \grn_reg[0] ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[9] ;
  wire [15:0]out;
  wire [15:0]p_0_in0_in;
  wire [15:0]p_1_in1_in;
  wire \rgf_c1bus_wb[4]_i_18 ;
  wire \rgf_c1bus_wb[4]_i_18_0 ;
  wire \rgf_c1bus_wb[4]_i_18_1 ;
  wire \rgf_c1bus_wb[4]_i_18_2 ;
  wire \rgf_c1bus_wb[4]_i_18_3 ;
  wire \rgf_c1bus_wb[4]_i_18_4 ;
  wire \rgf_c1bus_wb[4]_i_18_5 ;
  wire \rgf_c1bus_wb[4]_i_18_6 ;
  wire \rgf_c1bus_wb[4]_i_18_7 ;
  wire \rgf_c1bus_wb[4]_i_19 ;
  wire \rgf_c1bus_wb[4]_i_19_0 ;
  wire \rgf_c1bus_wb[4]_i_19_1 ;
  wire \rgf_c1bus_wb[4]_i_19_10 ;
  wire \rgf_c1bus_wb[4]_i_19_11 ;
  wire \rgf_c1bus_wb[4]_i_19_2 ;
  wire \rgf_c1bus_wb[4]_i_19_3 ;
  wire \rgf_c1bus_wb[4]_i_19_4 ;
  wire \rgf_c1bus_wb[4]_i_19_5 ;
  wire \rgf_c1bus_wb[4]_i_19_6 ;
  wire \rgf_c1bus_wb[4]_i_19_7 ;
  wire \rgf_c1bus_wb[4]_i_19_8 ;
  wire \rgf_c1bus_wb[4]_i_19_9 ;
  wire \rgf_c1bus_wb[4]_i_20 ;
  wire \rgf_c1bus_wb[4]_i_20_0 ;
  wire \rgf_c1bus_wb[4]_i_20_1 ;
  wire \rgf_c1bus_wb[4]_i_20_2 ;
  wire \rgf_c1bus_wb[4]_i_20_3 ;
  wire \rgf_c1bus_wb[4]_i_20_4 ;
  wire \rgf_c1bus_wb[4]_i_21 ;
  wire \rgf_c1bus_wb[4]_i_21_0 ;
  wire \rgf_c1bus_wb[4]_i_21_1 ;
  wire \rgf_c1bus_wb[4]_i_21_2 ;
  wire \rgf_c1bus_wb[4]_i_21_3 ;
  wire \rgf_c1bus_wb[4]_i_22 ;
  wire \rgf_c1bus_wb[4]_i_22_0 ;
  wire \rgf_c1bus_wb[4]_i_22_1 ;
  wire \rgf_c1bus_wb[4]_i_22_2 ;
  wire \rgf_c1bus_wb[4]_i_22_3 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_22_4 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_22_5 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_22_6 ;
  wire \rgf_c1bus_wb[4]_i_23 ;
  wire \rgf_c1bus_wb[4]_i_23_0 ;
  wire \rgf_c1bus_wb[4]_i_23_1 ;
  wire \rgf_c1bus_wb[4]_i_23_2 ;
  wire \rgf_c1bus_wb[4]_i_23_3 ;
  wire \sp_reg[0] ;
  wire \sp_reg[0]_0 ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[4]_i_207 ;
  wire \sr[4]_i_207_0 ;
  wire \sr[4]_i_207_1 ;
  wire \sr[4]_i_207_2 ;
  wire \sr[4]_i_207_3 ;
  wire \sr[4]_i_208 ;
  wire \sr[4]_i_208_0 ;
  wire \sr[4]_i_208_1 ;
  wire \sr[4]_i_208_2 ;
  wire \sr[4]_i_208_3 ;
  wire \sr[4]_i_210 ;
  wire \sr[4]_i_213 ;
  wire \sr[4]_i_213_0 ;
  wire \sr[4]_i_213_1 ;
  wire \sr[4]_i_213_2 ;
  wire \sr[4]_i_213_3 ;
  wire \sr[4]_i_215 ;
  wire \sr[4]_i_215_0 ;
  wire \sr[4]_i_215_1 ;
  wire \sr[4]_i_215_10 ;
  wire \sr[4]_i_215_11 ;
  wire \sr[4]_i_215_2 ;
  wire \sr[4]_i_215_3 ;
  wire \sr[4]_i_215_4 ;
  wire \sr[4]_i_215_5 ;
  wire \sr[4]_i_215_6 ;
  wire \sr[4]_i_215_7 ;
  wire \sr[4]_i_215_8 ;
  wire \sr[4]_i_215_9 ;
  wire \sr[4]_i_216 ;
  wire \sr[4]_i_216_0 ;
  wire \sr[4]_i_216_1 ;
  wire \sr[4]_i_216_10 ;
  wire \sr[4]_i_216_11 ;
  wire \sr[4]_i_216_2 ;
  wire \sr[4]_i_216_3 ;
  wire \sr[4]_i_216_4 ;
  wire \sr[4]_i_216_5 ;
  wire \sr[4]_i_216_6 ;
  wire \sr[4]_i_216_7 ;
  wire \sr[4]_i_216_8 ;
  wire \sr[4]_i_216_9 ;
  wire \sr[4]_i_217 ;
  wire \sr[4]_i_217_0 ;
  wire \sr[4]_i_217_1 ;
  wire \sr[4]_i_217_2 ;
  wire \sr[4]_i_217_3 ;
  wire \sr[4]_i_217_4 ;
  wire \sr[4]_i_217_5 ;
  wire \sr[4]_i_217_6 ;
  wire \sr[4]_i_217_7 ;
  wire \sr[4]_i_218 ;
  wire \sr[4]_i_218_0 ;
  wire \sr[4]_i_218_1 ;
  wire \sr[4]_i_218_10 ;
  wire \sr[4]_i_218_11 ;
  wire \sr[4]_i_218_2 ;
  wire \sr[4]_i_218_3 ;
  wire \sr[4]_i_218_4 ;
  wire \sr[4]_i_218_5 ;
  wire \sr[4]_i_218_6 ;
  wire \sr[4]_i_218_7 ;
  wire \sr[4]_i_218_8 ;
  wire \sr[4]_i_218_9 ;
  wire \sr[4]_i_219 ;
  wire \sr[4]_i_219_0 ;
  wire \sr[4]_i_219_1 ;
  wire \sr[4]_i_219_2 ;
  wire \sr[4]_i_219_3 ;
  wire \sr[4]_i_220 ;
  wire \sr[4]_i_220_0 ;
  wire \sr[4]_i_220_1 ;
  wire \sr[4]_i_220_2 ;
  wire \sr[4]_i_220_3 ;
  wire \sr[4]_i_224 ;
  wire \sr[4]_i_224_0 ;
  wire \sr[4]_i_224_1 ;
  wire \sr[4]_i_224_10 ;
  wire \sr[4]_i_224_11 ;
  wire \sr[4]_i_224_2 ;
  wire \sr[4]_i_224_3 ;
  wire \sr[4]_i_224_4 ;
  wire \sr[4]_i_224_5 ;
  wire \sr[4]_i_224_6 ;
  wire \sr[4]_i_224_7 ;
  wire \sr[4]_i_224_8 ;
  wire \sr[4]_i_224_9 ;
  wire \sr[4]_i_225 ;
  wire \sr[4]_i_225_0 ;
  wire \sr[4]_i_225_1 ;
  wire \sr[4]_i_225_10 ;
  wire \sr[4]_i_225_11 ;
  wire \sr[4]_i_225_2 ;
  wire \sr[4]_i_225_3 ;
  wire \sr[4]_i_225_4 ;
  wire \sr[4]_i_225_5 ;
  wire \sr[4]_i_225_6 ;
  wire \sr[4]_i_225_7 ;
  wire \sr[4]_i_225_8 ;
  wire \sr[4]_i_225_9 ;
  wire \sr_reg[0] ;
  wire \sr_reg[15] ;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[10] ;
  wire \tr_reg[10]_0 ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire \tr_reg[15] ;
  wire \tr_reg[15]_0 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[2] ;
  wire \tr_reg[2]_0 ;
  wire \tr_reg[3] ;
  wire \tr_reg[3]_0 ;
  wire \tr_reg[4] ;
  wire \tr_reg[4]_0 ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[8] ;
  wire \tr_reg[8]_0 ;
  wire \tr_reg[9] ;
  wire \tr_reg[9]_0 ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[0]_INST_0_i_1 
       (.I0(\tr_reg[0]_0 ),
        .I1(p_1_in1_in[0]),
        .I2(p_0_in0_in[0]),
        .I3(a1bus_sr[0]),
        .I4(a1bus_b13[0]),
        .I5(\sp_reg[0] ),
        .O(\tr_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[0]_INST_0_i_3 
       (.I0(out[0]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [0]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[0]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(O),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [0]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [0]),
        .I5(a1bus_sel_cr[0]),
        .O(\sp_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[10]_INST_0_i_1 
       (.I0(\tr_reg[10]_0 ),
        .I1(p_1_in1_in[10]),
        .I2(p_0_in0_in[10]),
        .I3(a1bus_sr[10]),
        .I4(a1bus_b13[10]),
        .I5(\badr[10]_INST_0_i_8_n_0 ),
        .O(\tr_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[10]_INST_0_i_3 
       (.I0(out[10]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [10]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[10]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[9]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [10]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [10]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[11]_INST_0_i_1 
       (.I0(\tr_reg[11]_0 ),
        .I1(p_1_in1_in[11]),
        .I2(p_0_in0_in[11]),
        .I3(a1bus_sr[11]),
        .I4(a1bus_b13[11]),
        .I5(\badr[11]_INST_0_i_8_n_0 ),
        .O(\tr_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[11]_INST_0_i_3 
       (.I0(out[11]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [11]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[11]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[10]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [11]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [11]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[11]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[12]_INST_0_i_1 
       (.I0(\tr_reg[12]_0 ),
        .I1(p_1_in1_in[12]),
        .I2(p_0_in0_in[12]),
        .I3(a1bus_sr[12]),
        .I4(a1bus_b13[12]),
        .I5(\badr[12]_INST_0_i_8_n_0 ),
        .O(\tr_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[12]_INST_0_i_3 
       (.I0(out[12]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [12]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[12]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[11]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [12]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [12]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[13]_INST_0_i_1 
       (.I0(\tr_reg[13]_0 ),
        .I1(p_1_in1_in[13]),
        .I2(p_0_in0_in[13]),
        .I3(a1bus_sr[13]),
        .I4(a1bus_b13[13]),
        .I5(\badr[13]_INST_0_i_8_n_0 ),
        .O(\tr_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[13]_INST_0_i_3 
       (.I0(out[13]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [13]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[13]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[12]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [13]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [13]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[14]_INST_0_i_1 
       (.I0(\tr_reg[14]_0 ),
        .I1(p_1_in1_in[14]),
        .I2(p_0_in0_in[14]),
        .I3(a1bus_sr[14]),
        .I4(a1bus_b13[14]),
        .I5(\badr[14]_INST_0_i_8_n_0 ),
        .O(\tr_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[14]_INST_0_i_3 
       (.I0(out[14]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [14]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[14]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[13]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [14]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [14]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[14]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_1 
       (.I0(\tr_reg[15]_0 ),
        .I1(p_1_in1_in[15]),
        .I2(p_0_in0_in[15]),
        .I3(a1bus_sr[15]),
        .I4(a1bus_b13[15]),
        .I5(\sp_reg[15] ),
        .O(\tr_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[15]_INST_0_i_3 
       (.I0(out[15]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [15]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[14]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [15]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [15]),
        .I5(a1bus_sel_cr[0]),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[1]_INST_0_i_1 
       (.I0(\tr_reg[1]_0 ),
        .I1(p_1_in1_in[1]),
        .I2(p_0_in0_in[1]),
        .I3(a1bus_sr[1]),
        .I4(a1bus_b13[1]),
        .I5(\badr[1]_INST_0_i_8_n_0 ),
        .O(\tr_reg[1] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[1]_INST_0_i_3 
       (.I0(out[1]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [1]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[0]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [1]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [1]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[2]_INST_0_i_1 
       (.I0(\tr_reg[2]_0 ),
        .I1(p_1_in1_in[2]),
        .I2(p_0_in0_in[2]),
        .I3(a1bus_sr[2]),
        .I4(a1bus_b13[2]),
        .I5(\badr[2]_INST_0_i_8_n_0 ),
        .O(\tr_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[2]_INST_0_i_3 
       (.I0(out[2]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [2]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[1]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [2]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [2]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[3]_INST_0_i_1 
       (.I0(\tr_reg[3]_0 ),
        .I1(p_1_in1_in[3]),
        .I2(p_0_in0_in[3]),
        .I3(a1bus_sr[3]),
        .I4(a1bus_b13[3]),
        .I5(\badr[3]_INST_0_i_8_n_0 ),
        .O(\tr_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[3]_INST_0_i_3 
       (.I0(out[3]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [3]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[2]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [3]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [3]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[4]_INST_0_i_1 
       (.I0(\tr_reg[4]_0 ),
        .I1(p_1_in1_in[4]),
        .I2(p_0_in0_in[4]),
        .I3(a1bus_sr[4]),
        .I4(a1bus_b13[4]),
        .I5(\badr[4]_INST_0_i_8_n_0 ),
        .O(\tr_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[4]_INST_0_i_3 
       (.I0(out[4]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [4]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[3]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [4]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [4]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[5]_INST_0_i_1 
       (.I0(\tr_reg[5]_0 ),
        .I1(p_1_in1_in[5]),
        .I2(p_0_in0_in[5]),
        .I3(a1bus_sr[5]),
        .I4(a1bus_b13[5]),
        .I5(\badr[5]_INST_0_i_8_n_0 ),
        .O(\tr_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[5]_INST_0_i_3 
       (.I0(out[5]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [5]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[4]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [5]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [5]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[5]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[6]_INST_0_i_1 
       (.I0(\tr_reg[6]_0 ),
        .I1(p_1_in1_in[6]),
        .I2(p_0_in0_in[6]),
        .I3(a1bus_sr[6]),
        .I4(a1bus_b13[6]),
        .I5(\badr[6]_INST_0_i_8_n_0 ),
        .O(\tr_reg[6] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[6]_INST_0_i_3 
       (.I0(out[6]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [6]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[5]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [6]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [6]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[7]_INST_0_i_1 
       (.I0(\tr_reg[7]_0 ),
        .I1(p_1_in1_in[7]),
        .I2(p_0_in0_in[7]),
        .I3(a1bus_sr[7]),
        .I4(a1bus_b13[7]),
        .I5(\badr[7]_INST_0_i_8_n_0 ),
        .O(\tr_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[7]_INST_0_i_3 
       (.I0(out[7]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [7]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[6]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [7]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [7]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[8]_INST_0_i_1 
       (.I0(\tr_reg[8]_0 ),
        .I1(p_1_in1_in[8]),
        .I2(p_0_in0_in[8]),
        .I3(a1bus_sr[8]),
        .I4(a1bus_b13[8]),
        .I5(\badr[8]_INST_0_i_8_n_0 ),
        .O(\tr_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[8]_INST_0_i_3 
       (.I0(out[8]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [8]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[7]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [8]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [8]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[9]_INST_0_i_1 
       (.I0(\tr_reg[9]_0 ),
        .I1(p_1_in1_in[9]),
        .I2(p_0_in0_in[9]),
        .I3(a1bus_sr[9]),
        .I4(a1bus_b13[9]),
        .I5(\badr[9]_INST_0_i_8_n_0 ),
        .O(\tr_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[9]_INST_0_i_3 
       (.I0(out[9]),
        .I1(a1bus_sel_cr[3]),
        .I2(\rgf_c1bus_wb[4]_i_22_4 [9]),
        .I3(a1bus_sel_cr[2]),
        .O(\tr_reg[9]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_8 
       (.I0(a1bus_sel_cr[4]),
        .I1(data3[8]),
        .I2(a1bus_sel_cr[1]),
        .I3(\rgf_c1bus_wb[4]_i_22_5 [9]),
        .I4(\rgf_c1bus_wb[4]_i_22_6 [9]),
        .I5(a1bus_sel_cr[0]),
        .O(\badr[9]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_32 
       (.I0(\badr[4]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_224_8 ),
        .I2(\sr[4]_i_224_9 ),
        .I3(\sr[4]_i_224_10 ),
        .I4(\sr[4]_i_224_11 ),
        .I5(a1bus_sr[4]),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_33 
       (.I0(\rgf_c1bus_wb[4]_i_18 ),
        .I1(\rgf_c1bus_wb[4]_i_18_0 ),
        .I2(\rgf_c1bus_wb[4]_i_18_1 ),
        .I3(\rgf_c1bus_wb[4]_i_18_2 ),
        .I4(\rgf_c1bus_wb[4]_i_18_3 ),
        .I5(\tr_reg[3]_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_34 
       (.I0(\badr[3]_INST_0_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_18_4 ),
        .I2(\rgf_c1bus_wb[4]_i_18_5 ),
        .I3(\rgf_c1bus_wb[4]_i_18_6 ),
        .I4(\rgf_c1bus_wb[4]_i_18_7 ),
        .I5(a1bus_sr[3]),
        .O(\sp_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_36 
       (.I0(\badr[2]_INST_0_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_19_4 ),
        .I2(\rgf_c1bus_wb[4]_i_19_5 ),
        .I3(\rgf_c1bus_wb[4]_i_19_6 ),
        .I4(\rgf_c1bus_wb[4]_i_19_7 ),
        .I5(a1bus_sr[2]),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_37 
       (.I0(\rgf_c1bus_wb[4]_i_19 ),
        .I1(\rgf_c1bus_wb[4]_i_19_0 ),
        .I2(\rgf_c1bus_wb[4]_i_19_1 ),
        .I3(\rgf_c1bus_wb[4]_i_19_2 ),
        .I4(\rgf_c1bus_wb[4]_i_19_3 ),
        .I5(\tr_reg[1]_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_38 
       (.I0(\badr[1]_INST_0_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_19_8 ),
        .I2(\rgf_c1bus_wb[4]_i_19_9 ),
        .I3(\rgf_c1bus_wb[4]_i_19_10 ),
        .I4(\rgf_c1bus_wb[4]_i_19_11 ),
        .I5(a1bus_sr[1]),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_40 
       (.I0(\sp_reg[15] ),
        .I1(\rgf_c1bus_wb[4]_i_22 ),
        .I2(\rgf_c1bus_wb[4]_i_20_4 ),
        .I3(\rgf_c1bus_wb[4]_i_22_0 ),
        .I4(\rgf_c1bus_wb[4]_i_22_1 ),
        .I5(a1bus_sr[15]),
        .O(\sp_reg[15]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_41 
       (.I0(\rgf_c1bus_wb[4]_i_20 ),
        .I1(\rgf_c1bus_wb[4]_i_20_0 ),
        .I2(\rgf_c1bus_wb[4]_i_20_1 ),
        .I3(\rgf_c1bus_wb[4]_i_20_2 ),
        .I4(\rgf_c1bus_wb[4]_i_20_3 ),
        .I5(\tr_reg[14]_0 ),
        .O(\grn_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_42 
       (.I0(\badr[14]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_216_4 ),
        .I2(\sr[4]_i_216_5 ),
        .I3(\sr[4]_i_216_6 ),
        .I4(\sr[4]_i_216_7 ),
        .I5(a1bus_sr[14]),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_44 
       (.I0(a1bus_sr[0]),
        .I1(\rgf_c1bus_wb[4]_i_21_1 ),
        .I2(\rgf_c1bus_wb[4]_i_21_0 ),
        .I3(\rgf_c1bus_wb[4]_i_21_2 ),
        .I4(\rgf_c1bus_wb[4]_i_21_3 ),
        .I5(\rgf_c1bus_wb[4]_i_21 ),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_45 
       (.I0(a1bus_sr[15]),
        .I1(\rgf_c1bus_wb[4]_i_22_1 ),
        .I2(\rgf_c1bus_wb[4]_i_22_0 ),
        .I3(\rgf_c1bus_wb[4]_i_22_2 ),
        .I4(\rgf_c1bus_wb[4]_i_22_3 ),
        .I5(\rgf_c1bus_wb[4]_i_22 ),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_47 
       (.I0(\rgf_c1bus_wb[4]_i_23 ),
        .I1(\rgf_c1bus_wb[4]_i_23_0 ),
        .I2(\rgf_c1bus_wb[4]_i_23_1 ),
        .I3(\rgf_c1bus_wb[4]_i_23_2 ),
        .I4(\rgf_c1bus_wb[4]_i_23_3 ),
        .I5(\tr_reg[15]_0 ),
        .O(\grn_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_48 
       (.I0(\badr[12]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_215_4 ),
        .I2(\sr[4]_i_215_5 ),
        .I3(\sr[4]_i_215_6 ),
        .I4(\sr[4]_i_215_7 ),
        .I5(a1bus_sr[12]),
        .O(\sp_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_50 
       (.I0(\badr[13]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_216_8 ),
        .I2(\sr[4]_i_216_9 ),
        .I3(\sr[4]_i_216_10 ),
        .I4(\sr[4]_i_216_11 ),
        .I5(a1bus_sr[13]),
        .O(\sp_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_51 
       (.I0(\sr[4]_i_216 ),
        .I1(\sr[4]_i_216_0 ),
        .I2(\sr[4]_i_216_1 ),
        .I3(\sr[4]_i_216_2 ),
        .I4(\sr[4]_i_216_3 ),
        .I5(\tr_reg[13]_0 ),
        .O(\grn_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_52 
       (.I0(\badr[5]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_224_4 ),
        .I2(\sr[4]_i_224_5 ),
        .I3(\sr[4]_i_224_6 ),
        .I4(\sr[4]_i_224_7 ),
        .I5(a1bus_sr[5]),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_53 
       (.I0(\sr[4]_i_219 ),
        .I1(\sr[4]_i_219_0 ),
        .I2(\sr[4]_i_219_1 ),
        .I3(\sr[4]_i_219_2 ),
        .I4(\sr[4]_i_219_3 ),
        .I5(\tr_reg[5]_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_54 
       (.I0(\badr[6]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_225_8 ),
        .I2(\sr[4]_i_225_9 ),
        .I3(\sr[4]_i_225_10 ),
        .I4(\sr[4]_i_225_11 ),
        .I5(a1bus_sr[6]),
        .O(\sp_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_56 
       (.I0(\badr[7]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_225_4 ),
        .I2(\sr[4]_i_225_5 ),
        .I3(\sr[4]_i_225_6 ),
        .I4(\sr[4]_i_225_7 ),
        .I5(a1bus_sr[7]),
        .O(\sp_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_57 
       (.I0(\sr[4]_i_217 ),
        .I1(\sr[4]_i_217_0 ),
        .I2(\sr[4]_i_217_1 ),
        .I3(\sr[4]_i_217_2 ),
        .I4(\sr[4]_i_217_3 ),
        .I5(\tr_reg[7]_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_58 
       (.I0(\badr[8]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_217_4 ),
        .I2(\sr[4]_i_217_5 ),
        .I3(\sr[4]_i_217_6 ),
        .I4(\sr[4]_i_217_7 ),
        .I5(a1bus_sr[8]),
        .O(\sp_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_60 
       (.I0(\badr[9]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_218_8 ),
        .I2(\sr[4]_i_218_9 ),
        .I3(\sr[4]_i_218_10 ),
        .I4(\sr[4]_i_218_11 ),
        .I5(a1bus_sr[9]),
        .O(\sp_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_61 
       (.I0(\sr[4]_i_218 ),
        .I1(\sr[4]_i_218_0 ),
        .I2(\sr[4]_i_218_1 ),
        .I3(\sr[4]_i_218_2 ),
        .I4(\sr[4]_i_218_3 ),
        .I5(\tr_reg[9]_0 ),
        .O(\grn_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_62 
       (.I0(\badr[10]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_218_4 ),
        .I2(\sr[4]_i_218_5 ),
        .I3(\sr[4]_i_218_6 ),
        .I4(\sr[4]_i_218_7 ),
        .I5(a1bus_sr[10]),
        .O(\sp_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_64 
       (.I0(\badr[11]_INST_0_i_8_n_0 ),
        .I1(\sr[4]_i_215_8 ),
        .I2(\sr[4]_i_215_9 ),
        .I3(\sr[4]_i_215_10 ),
        .I4(\sr[4]_i_215_11 ),
        .I5(a1bus_sr[11]),
        .O(\sp_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_65 
       (.I0(\sr[4]_i_215 ),
        .I1(\sr[4]_i_215_0 ),
        .I2(\sr[4]_i_215_1 ),
        .I3(\sr[4]_i_215_2 ),
        .I4(\sr[4]_i_215_3 ),
        .I5(\tr_reg[11]_0 ),
        .O(\grn_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_c1bus_wb[4]_i_67 
       (.I0(\sr[4]_i_220 ),
        .I1(\sr[4]_i_220_0 ),
        .I2(\sr[4]_i_220_1 ),
        .I3(\sr[4]_i_220_2 ),
        .I4(\sr[4]_i_220_3 ),
        .I5(\tr_reg[2]_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_235 
       (.I0(\sr[4]_i_207 ),
        .I1(\sr[4]_i_207_0 ),
        .I2(\sr[4]_i_207_1 ),
        .I3(\sr[4]_i_207_2 ),
        .I4(\sr[4]_i_207_3 ),
        .I5(\tr_reg[12]_0 ),
        .O(\grn_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_237 
       (.I0(\sr[4]_i_208 ),
        .I1(\sr[4]_i_208_0 ),
        .I2(\sr[4]_i_208_1 ),
        .I3(\sr[4]_i_208_2 ),
        .I4(\sr[4]_i_208_3 ),
        .I5(\tr_reg[10]_0 ),
        .O(\grn_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_239 
       (.I0(\sp_reg[0] ),
        .I1(\rgf_c1bus_wb[4]_i_21 ),
        .I2(\sr[4]_i_210 ),
        .I3(\rgf_c1bus_wb[4]_i_21_0 ),
        .I4(\rgf_c1bus_wb[4]_i_21_1 ),
        .I5(a1bus_sr[0]),
        .O(\sp_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_240 
       (.I0(\sr[4]_i_213 ),
        .I1(\sr[4]_i_213_0 ),
        .I2(\sr[4]_i_213_1 ),
        .I3(\sr[4]_i_213_2 ),
        .I4(\sr[4]_i_213_3 ),
        .I5(\tr_reg[0]_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_243 
       (.I0(\sr[4]_i_224 ),
        .I1(\sr[4]_i_224_0 ),
        .I2(\sr[4]_i_224_1 ),
        .I3(\sr[4]_i_224_2 ),
        .I4(\sr[4]_i_224_3 ),
        .I5(\tr_reg[4]_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_245 
       (.I0(\sr[4]_i_225 ),
        .I1(\sr[4]_i_225_0 ),
        .I2(\sr[4]_i_225_1 ),
        .I3(\sr[4]_i_225_2 ),
        .I4(\sr[4]_i_225_3 ),
        .I5(\tr_reg[6]_0 ),
        .O(\grn_reg[6] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_3
   (\sp_reg[15] ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[4] ,
    \sp_reg[3] ,
    \sp_reg[2] ,
    \sp_reg[1] ,
    \sp_reg[0] ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \tr_reg[15] ,
    \bdatw[15]_INST_0_i_1 ,
    \bdatw[15]_INST_0_i_1_0 ,
    \bdatw[15]_INST_0_i_1_1 ,
    \bdatw[15]_INST_0_i_1_2 ,
    b0bus_sr,
    \bdatw[14]_INST_0_i_1 ,
    \bdatw[14]_INST_0_i_1_0 ,
    \bdatw[14]_INST_0_i_1_1 ,
    \bdatw[14]_INST_0_i_1_2 ,
    \bdatw[13]_INST_0_i_1 ,
    \bdatw[13]_INST_0_i_1_0 ,
    \bdatw[13]_INST_0_i_1_1 ,
    \bdatw[13]_INST_0_i_1_2 ,
    \bdatw[12]_INST_0_i_1 ,
    \bdatw[12]_INST_0_i_1_0 ,
    \bdatw[12]_INST_0_i_1_1 ,
    \bdatw[12]_INST_0_i_1_2 ,
    \bdatw[11]_INST_0_i_1 ,
    \bdatw[11]_INST_0_i_1_0 ,
    \bdatw[11]_INST_0_i_1_1 ,
    \bdatw[11]_INST_0_i_1_2 ,
    \bdatw[10]_INST_0_i_1 ,
    \bdatw[10]_INST_0_i_1_0 ,
    \bdatw[10]_INST_0_i_1_1 ,
    \bdatw[10]_INST_0_i_1_2 ,
    \bdatw[9]_INST_0_i_1 ,
    \bdatw[9]_INST_0_i_1_0 ,
    \bdatw[9]_INST_0_i_1_1 ,
    \bdatw[9]_INST_0_i_1_2 ,
    \bdatw[8]_INST_0_i_1 ,
    \bdatw[8]_INST_0_i_1_0 ,
    \bdatw[8]_INST_0_i_1_1 ,
    \bdatw[8]_INST_0_i_1_2 ,
    \bbus_o[7]_INST_0_i_1 ,
    \bbus_o[7]_INST_0_i_1_0 ,
    \bbus_o[7]_INST_0_i_1_1 ,
    \bbus_o[7]_INST_0_i_1_2 ,
    \bbus_o[6]_INST_0_i_1 ,
    \bbus_o[6]_INST_0_i_1_0 ,
    \bbus_o[6]_INST_0_i_1_1 ,
    \bbus_o[6]_INST_0_i_1_2 ,
    \bbus_o[5]_INST_0_i_1 ,
    \bbus_o[5]_INST_0_i_1_0 ,
    \bbus_o[5]_INST_0_i_1_1 ,
    \bbus_o[5]_INST_0_i_1_2 ,
    \bbus_o[4]_INST_0_i_1 ,
    \bbus_o[4]_INST_0_i_1_0 ,
    \bbus_o[4]_INST_0_i_1_1 ,
    \bbus_o[4]_INST_0_i_1_2 ,
    \bbus_o[3]_INST_0_i_1 ,
    \bbus_o[3]_INST_0_i_1_0 ,
    \bbus_o[3]_INST_0_i_1_1 ,
    \bbus_o[3]_INST_0_i_1_2 ,
    \bbus_o[2]_INST_0_i_1 ,
    \bbus_o[2]_INST_0_i_1_0 ,
    \bbus_o[2]_INST_0_i_1_1 ,
    \bbus_o[2]_INST_0_i_1_2 ,
    \bbus_o[1]_INST_0_i_1 ,
    \bbus_o[1]_INST_0_i_1_0 ,
    \bbus_o[1]_INST_0_i_1_1 ,
    \bbus_o[1]_INST_0_i_1_2 ,
    \bbus_o[0]_INST_0_i_1 ,
    \bbus_o[0]_INST_0_i_1_0 ,
    \bbus_o[0]_INST_0_i_1_1 ,
    \bbus_o[0]_INST_0_i_1_2 ,
    out,
    b0bus_sel_cr,
    \bdatw[15]_INST_0_i_1_3 ,
    O,
    \bdatw[15]_INST_0_i_11_0 ,
    \bdatw[15]_INST_0_i_11_1 ,
    data3);
  output \sp_reg[15] ;
  output \sp_reg[14] ;
  output \sp_reg[13] ;
  output \sp_reg[12] ;
  output \sp_reg[11] ;
  output \sp_reg[10] ;
  output \sp_reg[9] ;
  output \sp_reg[8] ;
  output \sp_reg[7] ;
  output \sp_reg[6] ;
  output \sp_reg[5] ;
  output \sp_reg[4] ;
  output \sp_reg[3] ;
  output \sp_reg[2] ;
  output \sp_reg[1] ;
  output \sp_reg[0] ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \tr_reg[15] ;
  input \bdatw[15]_INST_0_i_1 ;
  input \bdatw[15]_INST_0_i_1_0 ;
  input \bdatw[15]_INST_0_i_1_1 ;
  input \bdatw[15]_INST_0_i_1_2 ;
  input [15:0]b0bus_sr;
  input \bdatw[14]_INST_0_i_1 ;
  input \bdatw[14]_INST_0_i_1_0 ;
  input \bdatw[14]_INST_0_i_1_1 ;
  input \bdatw[14]_INST_0_i_1_2 ;
  input \bdatw[13]_INST_0_i_1 ;
  input \bdatw[13]_INST_0_i_1_0 ;
  input \bdatw[13]_INST_0_i_1_1 ;
  input \bdatw[13]_INST_0_i_1_2 ;
  input \bdatw[12]_INST_0_i_1 ;
  input \bdatw[12]_INST_0_i_1_0 ;
  input \bdatw[12]_INST_0_i_1_1 ;
  input \bdatw[12]_INST_0_i_1_2 ;
  input \bdatw[11]_INST_0_i_1 ;
  input \bdatw[11]_INST_0_i_1_0 ;
  input \bdatw[11]_INST_0_i_1_1 ;
  input \bdatw[11]_INST_0_i_1_2 ;
  input \bdatw[10]_INST_0_i_1 ;
  input \bdatw[10]_INST_0_i_1_0 ;
  input \bdatw[10]_INST_0_i_1_1 ;
  input \bdatw[10]_INST_0_i_1_2 ;
  input \bdatw[9]_INST_0_i_1 ;
  input \bdatw[9]_INST_0_i_1_0 ;
  input \bdatw[9]_INST_0_i_1_1 ;
  input \bdatw[9]_INST_0_i_1_2 ;
  input \bdatw[8]_INST_0_i_1 ;
  input \bdatw[8]_INST_0_i_1_0 ;
  input \bdatw[8]_INST_0_i_1_1 ;
  input \bdatw[8]_INST_0_i_1_2 ;
  input \bbus_o[7]_INST_0_i_1 ;
  input \bbus_o[7]_INST_0_i_1_0 ;
  input \bbus_o[7]_INST_0_i_1_1 ;
  input \bbus_o[7]_INST_0_i_1_2 ;
  input \bbus_o[6]_INST_0_i_1 ;
  input \bbus_o[6]_INST_0_i_1_0 ;
  input \bbus_o[6]_INST_0_i_1_1 ;
  input \bbus_o[6]_INST_0_i_1_2 ;
  input \bbus_o[5]_INST_0_i_1 ;
  input \bbus_o[5]_INST_0_i_1_0 ;
  input \bbus_o[5]_INST_0_i_1_1 ;
  input \bbus_o[5]_INST_0_i_1_2 ;
  input \bbus_o[4]_INST_0_i_1 ;
  input \bbus_o[4]_INST_0_i_1_0 ;
  input \bbus_o[4]_INST_0_i_1_1 ;
  input \bbus_o[4]_INST_0_i_1_2 ;
  input \bbus_o[3]_INST_0_i_1 ;
  input \bbus_o[3]_INST_0_i_1_0 ;
  input \bbus_o[3]_INST_0_i_1_1 ;
  input \bbus_o[3]_INST_0_i_1_2 ;
  input \bbus_o[2]_INST_0_i_1 ;
  input \bbus_o[2]_INST_0_i_1_0 ;
  input \bbus_o[2]_INST_0_i_1_1 ;
  input \bbus_o[2]_INST_0_i_1_2 ;
  input \bbus_o[1]_INST_0_i_1 ;
  input \bbus_o[1]_INST_0_i_1_0 ;
  input \bbus_o[1]_INST_0_i_1_1 ;
  input \bbus_o[1]_INST_0_i_1_2 ;
  input \bbus_o[0]_INST_0_i_1 ;
  input \bbus_o[0]_INST_0_i_1_0 ;
  input \bbus_o[0]_INST_0_i_1_1 ;
  input \bbus_o[0]_INST_0_i_1_2 ;
  input [15:0]out;
  input [4:0]b0bus_sel_cr;
  input [15:0]\bdatw[15]_INST_0_i_1_3 ;
  input [0:0]O;
  input [15:0]\bdatw[15]_INST_0_i_11_0 ;
  input [15:0]\bdatw[15]_INST_0_i_11_1 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [4:0]b0bus_sel_cr;
  wire [15:0]b0bus_sr;
  wire \bbus_o[0]_INST_0_i_1 ;
  wire \bbus_o[0]_INST_0_i_17_n_0 ;
  wire \bbus_o[0]_INST_0_i_1_0 ;
  wire \bbus_o[0]_INST_0_i_1_1 ;
  wire \bbus_o[0]_INST_0_i_1_2 ;
  wire \bbus_o[1]_INST_0_i_1 ;
  wire \bbus_o[1]_INST_0_i_16_n_0 ;
  wire \bbus_o[1]_INST_0_i_1_0 ;
  wire \bbus_o[1]_INST_0_i_1_1 ;
  wire \bbus_o[1]_INST_0_i_1_2 ;
  wire \bbus_o[2]_INST_0_i_1 ;
  wire \bbus_o[2]_INST_0_i_17_n_0 ;
  wire \bbus_o[2]_INST_0_i_1_0 ;
  wire \bbus_o[2]_INST_0_i_1_1 ;
  wire \bbus_o[2]_INST_0_i_1_2 ;
  wire \bbus_o[3]_INST_0_i_1 ;
  wire \bbus_o[3]_INST_0_i_17_n_0 ;
  wire \bbus_o[3]_INST_0_i_1_0 ;
  wire \bbus_o[3]_INST_0_i_1_1 ;
  wire \bbus_o[3]_INST_0_i_1_2 ;
  wire \bbus_o[4]_INST_0_i_1 ;
  wire \bbus_o[4]_INST_0_i_19_n_0 ;
  wire \bbus_o[4]_INST_0_i_1_0 ;
  wire \bbus_o[4]_INST_0_i_1_1 ;
  wire \bbus_o[4]_INST_0_i_1_2 ;
  wire \bbus_o[5]_INST_0_i_1 ;
  wire \bbus_o[5]_INST_0_i_13_n_0 ;
  wire \bbus_o[5]_INST_0_i_1_0 ;
  wire \bbus_o[5]_INST_0_i_1_1 ;
  wire \bbus_o[5]_INST_0_i_1_2 ;
  wire \bbus_o[6]_INST_0_i_1 ;
  wire \bbus_o[6]_INST_0_i_13_n_0 ;
  wire \bbus_o[6]_INST_0_i_1_0 ;
  wire \bbus_o[6]_INST_0_i_1_1 ;
  wire \bbus_o[6]_INST_0_i_1_2 ;
  wire \bbus_o[7]_INST_0_i_1 ;
  wire \bbus_o[7]_INST_0_i_13_n_0 ;
  wire \bbus_o[7]_INST_0_i_1_0 ;
  wire \bbus_o[7]_INST_0_i_1_1 ;
  wire \bbus_o[7]_INST_0_i_1_2 ;
  wire \bdatw[10]_INST_0_i_1 ;
  wire \bdatw[10]_INST_0_i_1_0 ;
  wire \bdatw[10]_INST_0_i_1_1 ;
  wire \bdatw[10]_INST_0_i_1_2 ;
  wire \bdatw[10]_INST_0_i_23_n_0 ;
  wire \bdatw[11]_INST_0_i_1 ;
  wire \bdatw[11]_INST_0_i_1_0 ;
  wire \bdatw[11]_INST_0_i_1_1 ;
  wire \bdatw[11]_INST_0_i_1_2 ;
  wire \bdatw[11]_INST_0_i_22_n_0 ;
  wire \bdatw[12]_INST_0_i_1 ;
  wire \bdatw[12]_INST_0_i_1_0 ;
  wire \bdatw[12]_INST_0_i_1_1 ;
  wire \bdatw[12]_INST_0_i_1_2 ;
  wire \bdatw[12]_INST_0_i_22_n_0 ;
  wire \bdatw[13]_INST_0_i_1 ;
  wire \bdatw[13]_INST_0_i_1_0 ;
  wire \bdatw[13]_INST_0_i_1_1 ;
  wire \bdatw[13]_INST_0_i_1_2 ;
  wire \bdatw[13]_INST_0_i_22_n_0 ;
  wire \bdatw[14]_INST_0_i_1 ;
  wire \bdatw[14]_INST_0_i_1_0 ;
  wire \bdatw[14]_INST_0_i_1_1 ;
  wire \bdatw[14]_INST_0_i_1_2 ;
  wire \bdatw[14]_INST_0_i_23_n_0 ;
  wire \bdatw[15]_INST_0_i_1 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_11_1 ;
  wire \bdatw[15]_INST_0_i_1_0 ;
  wire \bdatw[15]_INST_0_i_1_1 ;
  wire \bdatw[15]_INST_0_i_1_2 ;
  wire [15:0]\bdatw[15]_INST_0_i_1_3 ;
  wire \bdatw[15]_INST_0_i_32_n_0 ;
  wire \bdatw[8]_INST_0_i_1 ;
  wire \bdatw[8]_INST_0_i_1_0 ;
  wire \bdatw[8]_INST_0_i_1_1 ;
  wire \bdatw[8]_INST_0_i_1_2 ;
  wire \bdatw[8]_INST_0_i_22_n_0 ;
  wire \bdatw[9]_INST_0_i_1 ;
  wire \bdatw[9]_INST_0_i_1_0 ;
  wire \bdatw[9]_INST_0_i_1_1 ;
  wire \bdatw[9]_INST_0_i_1_2 ;
  wire \bdatw[9]_INST_0_i_22_n_0 ;
  wire [14:0]data3;
  wire [15:0]out;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \tr_reg[0] ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[15] ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[0]_INST_0_i_17 
       (.I0(b0bus_sel_cr[4]),
        .I1(O),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [0]),
        .I4(\bdatw[15]_INST_0_i_11_1 [0]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[0]_INST_0_i_4 
       (.I0(out[0]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [0]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[0]_INST_0_i_7 
       (.I0(\bbus_o[0]_INST_0_i_17_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1 ),
        .I2(\bbus_o[0]_INST_0_i_1_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_1 ),
        .I4(\bbus_o[0]_INST_0_i_1_2 ),
        .I5(b0bus_sr[0]),
        .O(\sp_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[1]_INST_0_i_16 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[0]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [1]),
        .I4(\bdatw[15]_INST_0_i_11_1 [1]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[1]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[1]_INST_0_i_4 
       (.I0(out[1]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [1]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[1]_INST_0_i_7 
       (.I0(\bbus_o[1]_INST_0_i_16_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1 ),
        .I2(\bbus_o[1]_INST_0_i_1_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_1 ),
        .I4(\bbus_o[1]_INST_0_i_1_2 ),
        .I5(b0bus_sr[1]),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[2]_INST_0_i_17 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[1]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [2]),
        .I4(\bdatw[15]_INST_0_i_11_1 [2]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[2]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[2]_INST_0_i_4 
       (.I0(out[2]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [2]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[2]_INST_0_i_7 
       (.I0(\bbus_o[2]_INST_0_i_17_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1 ),
        .I2(\bbus_o[2]_INST_0_i_1_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_1 ),
        .I4(\bbus_o[2]_INST_0_i_1_2 ),
        .I5(b0bus_sr[2]),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[3]_INST_0_i_17 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[2]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [3]),
        .I4(\bdatw[15]_INST_0_i_11_1 [3]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[3]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[3]_INST_0_i_4 
       (.I0(out[3]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [3]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[3]_INST_0_i_7 
       (.I0(\bbus_o[3]_INST_0_i_17_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1 ),
        .I2(\bbus_o[3]_INST_0_i_1_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_1 ),
        .I4(\bbus_o[3]_INST_0_i_1_2 ),
        .I5(b0bus_sr[3]),
        .O(\sp_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[4]_INST_0_i_19 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[3]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [4]),
        .I4(\bdatw[15]_INST_0_i_11_1 [4]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[4]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[4]_INST_0_i_4 
       (.I0(out[4]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [4]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[4]_INST_0_i_7 
       (.I0(\bbus_o[4]_INST_0_i_19_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1 ),
        .I2(\bbus_o[4]_INST_0_i_1_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_1 ),
        .I4(\bbus_o[4]_INST_0_i_1_2 ),
        .I5(b0bus_sr[4]),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[5]_INST_0_i_13 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[4]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [5]),
        .I4(\bdatw[15]_INST_0_i_11_1 [5]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[5]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[5]_INST_0_i_4 
       (.I0(out[5]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [5]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[5]_INST_0_i_7 
       (.I0(\bbus_o[5]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1 ),
        .I2(\bbus_o[5]_INST_0_i_1_0 ),
        .I3(\bbus_o[5]_INST_0_i_1_1 ),
        .I4(\bbus_o[5]_INST_0_i_1_2 ),
        .I5(b0bus_sr[5]),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[6]_INST_0_i_13 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[5]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [6]),
        .I4(\bdatw[15]_INST_0_i_11_1 [6]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[6]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[6]_INST_0_i_4 
       (.I0(out[6]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [6]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[6]_INST_0_i_7 
       (.I0(\bbus_o[6]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[6]_INST_0_i_1 ),
        .I2(\bbus_o[6]_INST_0_i_1_0 ),
        .I3(\bbus_o[6]_INST_0_i_1_1 ),
        .I4(\bbus_o[6]_INST_0_i_1_2 ),
        .I5(b0bus_sr[6]),
        .O(\sp_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bbus_o[7]_INST_0_i_13 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[6]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [7]),
        .I4(\bdatw[15]_INST_0_i_11_1 [7]),
        .I5(b0bus_sel_cr[0]),
        .O(\bbus_o[7]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bbus_o[7]_INST_0_i_4 
       (.I0(out[7]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [7]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[7]_INST_0_i_7 
       (.I0(\bbus_o[7]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_1 ),
        .I2(\bbus_o[7]_INST_0_i_1_0 ),
        .I3(\bbus_o[7]_INST_0_i_1_1 ),
        .I4(\bbus_o[7]_INST_0_i_1_2 ),
        .I5(b0bus_sr[7]),
        .O(\sp_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_23 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[9]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [10]),
        .I4(\bdatw[15]_INST_0_i_11_1 [10]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[10]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[10]_INST_0_i_6 
       (.I0(out[10]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [10]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[10]_INST_0_i_9 
       (.I0(\bdatw[10]_INST_0_i_23_n_0 ),
        .I1(\bdatw[10]_INST_0_i_1 ),
        .I2(\bdatw[10]_INST_0_i_1_0 ),
        .I3(\bdatw[10]_INST_0_i_1_1 ),
        .I4(\bdatw[10]_INST_0_i_1_2 ),
        .I5(b0bus_sr[10]),
        .O(\sp_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_22 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[10]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [11]),
        .I4(\bdatw[15]_INST_0_i_11_1 [11]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[11]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[11]_INST_0_i_6 
       (.I0(out[11]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [11]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[11]_INST_0_i_9 
       (.I0(\bdatw[11]_INST_0_i_22_n_0 ),
        .I1(\bdatw[11]_INST_0_i_1 ),
        .I2(\bdatw[11]_INST_0_i_1_0 ),
        .I3(\bdatw[11]_INST_0_i_1_1 ),
        .I4(\bdatw[11]_INST_0_i_1_2 ),
        .I5(b0bus_sr[11]),
        .O(\sp_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_22 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[11]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [12]),
        .I4(\bdatw[15]_INST_0_i_11_1 [12]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[12]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[12]_INST_0_i_6 
       (.I0(out[12]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [12]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[12]_INST_0_i_9 
       (.I0(\bdatw[12]_INST_0_i_22_n_0 ),
        .I1(\bdatw[12]_INST_0_i_1 ),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\bdatw[12]_INST_0_i_1_1 ),
        .I4(\bdatw[12]_INST_0_i_1_2 ),
        .I5(b0bus_sr[12]),
        .O(\sp_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_22 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[12]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [13]),
        .I4(\bdatw[15]_INST_0_i_11_1 [13]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[13]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[13]_INST_0_i_6 
       (.I0(out[13]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [13]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_9 
       (.I0(\bdatw[13]_INST_0_i_22_n_0 ),
        .I1(\bdatw[13]_INST_0_i_1 ),
        .I2(\bdatw[13]_INST_0_i_1_0 ),
        .I3(\bdatw[13]_INST_0_i_1_1 ),
        .I4(\bdatw[13]_INST_0_i_1_2 ),
        .I5(b0bus_sr[13]),
        .O(\sp_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_23 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[13]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [14]),
        .I4(\bdatw[15]_INST_0_i_11_1 [14]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[14]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[14]_INST_0_i_6 
       (.I0(out[14]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [14]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[14]_INST_0_i_9 
       (.I0(\bdatw[14]_INST_0_i_23_n_0 ),
        .I1(\bdatw[14]_INST_0_i_1 ),
        .I2(\bdatw[14]_INST_0_i_1_0 ),
        .I3(\bdatw[14]_INST_0_i_1_1 ),
        .I4(\bdatw[14]_INST_0_i_1_2 ),
        .I5(b0bus_sr[14]),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_32_n_0 ),
        .I1(\bdatw[15]_INST_0_i_1 ),
        .I2(\bdatw[15]_INST_0_i_1_0 ),
        .I3(\bdatw[15]_INST_0_i_1_1 ),
        .I4(\bdatw[15]_INST_0_i_1_2 ),
        .I5(b0bus_sr[15]),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_32 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[14]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [15]),
        .I4(\bdatw[15]_INST_0_i_11_1 [15]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[15]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[15]_INST_0_i_8 
       (.I0(out[15]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [15]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_22 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[7]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [8]),
        .I4(\bdatw[15]_INST_0_i_11_1 [8]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[8]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[8]_INST_0_i_6 
       (.I0(out[8]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [8]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(\bdatw[8]_INST_0_i_22_n_0 ),
        .I1(\bdatw[8]_INST_0_i_1 ),
        .I2(\bdatw[8]_INST_0_i_1_0 ),
        .I3(\bdatw[8]_INST_0_i_1_1 ),
        .I4(\bdatw[8]_INST_0_i_1_2 ),
        .I5(b0bus_sr[8]),
        .O(\sp_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_22 
       (.I0(b0bus_sel_cr[4]),
        .I1(data3[8]),
        .I2(b0bus_sel_cr[1]),
        .I3(\bdatw[15]_INST_0_i_11_0 [9]),
        .I4(\bdatw[15]_INST_0_i_11_1 [9]),
        .I5(b0bus_sel_cr[0]),
        .O(\bdatw[9]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[9]_INST_0_i_6 
       (.I0(out[9]),
        .I1(b0bus_sel_cr[3]),
        .I2(\bdatw[15]_INST_0_i_1_3 [9]),
        .I3(b0bus_sel_cr[2]),
        .O(\tr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[9]_INST_0_i_9 
       (.I0(\bdatw[9]_INST_0_i_22_n_0 ),
        .I1(\bdatw[9]_INST_0_i_1 ),
        .I2(\bdatw[9]_INST_0_i_1_0 ),
        .I3(\bdatw[9]_INST_0_i_1_1 ),
        .I4(\bdatw[9]_INST_0_i_1_2 ),
        .I5(b0bus_sr[9]),
        .O(\sp_reg[9] ));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_bus" *) 
module mcss_rgf_bus_4
   (\iv_reg[15] ,
    \sr_reg[15] ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sr_reg[4] ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sr_reg[0] ,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \sp_reg[0] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \bdatw[15]_INST_0_i_2 ,
    \bdatw[15]_INST_0_i_2_0 ,
    b1bus_sel_cr,
    out,
    \bdatw[15]_INST_0_i_2_1 ,
    \bdatw[15]_INST_0_i_2_2 ,
    \bdatw[15]_INST_0_i_2_3 ,
    \bdatw[15]_INST_0_i_2_4 ,
    \bdatw[14]_INST_0_i_2 ,
    \bdatw[14]_INST_0_i_2_0 ,
    \bdatw[14]_INST_0_i_2_1 ,
    \bdatw[14]_INST_0_i_2_2 ,
    b1bus_sr,
    \bdatw[13]_INST_0_i_2 ,
    \bdatw[13]_INST_0_i_2_0 ,
    \bdatw[13]_INST_0_i_2_1 ,
    \bdatw[13]_INST_0_i_2_2 ,
    \bdatw[12]_INST_0_i_2 ,
    \bdatw[12]_INST_0_i_2_0 ,
    \bdatw[12]_INST_0_i_2_1 ,
    \bdatw[12]_INST_0_i_2_2 ,
    \bdatw[11]_INST_0_i_2 ,
    \bdatw[11]_INST_0_i_2_0 ,
    \bdatw[11]_INST_0_i_2_1 ,
    \bdatw[11]_INST_0_i_2_2 ,
    \bdatw[10]_INST_0_i_2 ,
    \bdatw[10]_INST_0_i_2_0 ,
    \bdatw[10]_INST_0_i_2_1 ,
    \bdatw[10]_INST_0_i_2_2 ,
    \bdatw[9]_INST_0_i_2 ,
    \bdatw[9]_INST_0_i_2_0 ,
    \bdatw[9]_INST_0_i_2_1 ,
    \bdatw[9]_INST_0_i_2_2 ,
    \bdatw[8]_INST_0_i_2 ,
    \bdatw[8]_INST_0_i_2_0 ,
    \bdatw[8]_INST_0_i_2_1 ,
    \bdatw[8]_INST_0_i_2_2 ,
    \bdatw[15]_INST_0_i_16 ,
    \bdatw[15]_INST_0_i_16_0 ,
    \bdatw[15]_INST_0_i_16_1 ,
    \bdatw[15]_INST_0_i_16_2 ,
    \bdatw[14]_INST_0_i_16 ,
    \bdatw[14]_INST_0_i_16_0 ,
    \bdatw[14]_INST_0_i_16_1 ,
    \bdatw[14]_INST_0_i_16_2 ,
    \bdatw[13]_INST_0_i_16 ,
    \bdatw[13]_INST_0_i_16_0 ,
    \bdatw[13]_INST_0_i_16_1 ,
    \bdatw[13]_INST_0_i_16_2 ,
    \bdatw[12]_INST_0_i_16 ,
    \bdatw[12]_INST_0_i_16_0 ,
    \bdatw[12]_INST_0_i_16_1 ,
    \bdatw[12]_INST_0_i_16_2 ,
    \bdatw[12]_INST_0_i_16_3 ,
    \bdatw[11]_INST_0_i_16 ,
    \bdatw[11]_INST_0_i_16_0 ,
    \bdatw[11]_INST_0_i_16_1 ,
    \bdatw[11]_INST_0_i_16_2 ,
    \bdatw[11]_INST_0_i_16_3 ,
    \bdatw[10]_INST_0_i_16 ,
    \bdatw[10]_INST_0_i_16_0 ,
    \bdatw[10]_INST_0_i_16_1 ,
    \bdatw[10]_INST_0_i_16_2 ,
    \bdatw[10]_INST_0_i_16_3 ,
    \bdatw[9]_INST_0_i_16 ,
    \bdatw[9]_INST_0_i_16_0 ,
    \bdatw[9]_INST_0_i_16_1 ,
    \bdatw[9]_INST_0_i_16_2 ,
    \bdatw[9]_INST_0_i_16_3 ,
    \bdatw[8]_INST_0_i_16 ,
    \bdatw[8]_INST_0_i_16_0 ,
    \bdatw[8]_INST_0_i_16_1 ,
    \bdatw[8]_INST_0_i_16_2 ,
    \bdatw[8]_INST_0_i_16_3 ,
    O,
    \bdatw[15]_INST_0_i_15_0 ,
    \bdatw[15]_INST_0_i_15_1 ,
    data3);
  output \iv_reg[15] ;
  output \sr_reg[15] ;
  output \sp_reg[14] ;
  output \sp_reg[13] ;
  output \sp_reg[12] ;
  output \sp_reg[11] ;
  output \sp_reg[10] ;
  output \sp_reg[9] ;
  output \sp_reg[8] ;
  output \sp_reg[7] ;
  output \sp_reg[6] ;
  output \sp_reg[5] ;
  output \sr_reg[4] ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sr_reg[0] ;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \sp_reg[0] ;
  output \sp_reg[1] ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  input \bdatw[15]_INST_0_i_2 ;
  input \bdatw[15]_INST_0_i_2_0 ;
  input [5:0]b1bus_sel_cr;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_2_1 ;
  input \bdatw[15]_INST_0_i_2_2 ;
  input \bdatw[15]_INST_0_i_2_3 ;
  input [0:0]\bdatw[15]_INST_0_i_2_4 ;
  input \bdatw[14]_INST_0_i_2 ;
  input \bdatw[14]_INST_0_i_2_0 ;
  input \bdatw[14]_INST_0_i_2_1 ;
  input \bdatw[14]_INST_0_i_2_2 ;
  input [14:0]b1bus_sr;
  input \bdatw[13]_INST_0_i_2 ;
  input \bdatw[13]_INST_0_i_2_0 ;
  input \bdatw[13]_INST_0_i_2_1 ;
  input \bdatw[13]_INST_0_i_2_2 ;
  input \bdatw[12]_INST_0_i_2 ;
  input \bdatw[12]_INST_0_i_2_0 ;
  input \bdatw[12]_INST_0_i_2_1 ;
  input \bdatw[12]_INST_0_i_2_2 ;
  input \bdatw[11]_INST_0_i_2 ;
  input \bdatw[11]_INST_0_i_2_0 ;
  input \bdatw[11]_INST_0_i_2_1 ;
  input \bdatw[11]_INST_0_i_2_2 ;
  input \bdatw[10]_INST_0_i_2 ;
  input \bdatw[10]_INST_0_i_2_0 ;
  input \bdatw[10]_INST_0_i_2_1 ;
  input \bdatw[10]_INST_0_i_2_2 ;
  input \bdatw[9]_INST_0_i_2 ;
  input \bdatw[9]_INST_0_i_2_0 ;
  input \bdatw[9]_INST_0_i_2_1 ;
  input \bdatw[9]_INST_0_i_2_2 ;
  input \bdatw[8]_INST_0_i_2 ;
  input \bdatw[8]_INST_0_i_2_0 ;
  input \bdatw[8]_INST_0_i_2_1 ;
  input \bdatw[8]_INST_0_i_2_2 ;
  input \bdatw[15]_INST_0_i_16 ;
  input \bdatw[15]_INST_0_i_16_0 ;
  input \bdatw[15]_INST_0_i_16_1 ;
  input \bdatw[15]_INST_0_i_16_2 ;
  input \bdatw[14]_INST_0_i_16 ;
  input \bdatw[14]_INST_0_i_16_0 ;
  input \bdatw[14]_INST_0_i_16_1 ;
  input \bdatw[14]_INST_0_i_16_2 ;
  input \bdatw[13]_INST_0_i_16 ;
  input \bdatw[13]_INST_0_i_16_0 ;
  input \bdatw[13]_INST_0_i_16_1 ;
  input \bdatw[13]_INST_0_i_16_2 ;
  input \bdatw[12]_INST_0_i_16 ;
  input \bdatw[12]_INST_0_i_16_0 ;
  input \bdatw[12]_INST_0_i_16_1 ;
  input \bdatw[12]_INST_0_i_16_2 ;
  input \bdatw[12]_INST_0_i_16_3 ;
  input \bdatw[11]_INST_0_i_16 ;
  input \bdatw[11]_INST_0_i_16_0 ;
  input \bdatw[11]_INST_0_i_16_1 ;
  input \bdatw[11]_INST_0_i_16_2 ;
  input \bdatw[11]_INST_0_i_16_3 ;
  input \bdatw[10]_INST_0_i_16 ;
  input \bdatw[10]_INST_0_i_16_0 ;
  input \bdatw[10]_INST_0_i_16_1 ;
  input \bdatw[10]_INST_0_i_16_2 ;
  input \bdatw[10]_INST_0_i_16_3 ;
  input \bdatw[9]_INST_0_i_16 ;
  input \bdatw[9]_INST_0_i_16_0 ;
  input \bdatw[9]_INST_0_i_16_1 ;
  input \bdatw[9]_INST_0_i_16_2 ;
  input \bdatw[9]_INST_0_i_16_3 ;
  input \bdatw[8]_INST_0_i_16 ;
  input \bdatw[8]_INST_0_i_16_0 ;
  input \bdatw[8]_INST_0_i_16_1 ;
  input \bdatw[8]_INST_0_i_16_2 ;
  input \bdatw[8]_INST_0_i_16_3 ;
  input [0:0]O;
  input [15:0]\bdatw[15]_INST_0_i_15_0 ;
  input [15:0]\bdatw[15]_INST_0_i_15_1 ;
  input [14:0]data3;

  wire [0:0]O;
  wire [5:0]b1bus_sel_cr;
  wire [14:0]b1bus_sr;
  wire \bdatw[10]_INST_0_i_16 ;
  wire \bdatw[10]_INST_0_i_16_0 ;
  wire \bdatw[10]_INST_0_i_16_1 ;
  wire \bdatw[10]_INST_0_i_16_2 ;
  wire \bdatw[10]_INST_0_i_16_3 ;
  wire \bdatw[10]_INST_0_i_2 ;
  wire \bdatw[10]_INST_0_i_2_0 ;
  wire \bdatw[10]_INST_0_i_2_1 ;
  wire \bdatw[10]_INST_0_i_2_2 ;
  wire \bdatw[10]_INST_0_i_34_n_0 ;
  wire \bdatw[11]_INST_0_i_16 ;
  wire \bdatw[11]_INST_0_i_16_0 ;
  wire \bdatw[11]_INST_0_i_16_1 ;
  wire \bdatw[11]_INST_0_i_16_2 ;
  wire \bdatw[11]_INST_0_i_16_3 ;
  wire \bdatw[11]_INST_0_i_2 ;
  wire \bdatw[11]_INST_0_i_2_0 ;
  wire \bdatw[11]_INST_0_i_2_1 ;
  wire \bdatw[11]_INST_0_i_2_2 ;
  wire \bdatw[11]_INST_0_i_34_n_0 ;
  wire \bdatw[12]_INST_0_i_16 ;
  wire \bdatw[12]_INST_0_i_16_0 ;
  wire \bdatw[12]_INST_0_i_16_1 ;
  wire \bdatw[12]_INST_0_i_16_2 ;
  wire \bdatw[12]_INST_0_i_16_3 ;
  wire \bdatw[12]_INST_0_i_2 ;
  wire \bdatw[12]_INST_0_i_2_0 ;
  wire \bdatw[12]_INST_0_i_2_1 ;
  wire \bdatw[12]_INST_0_i_2_2 ;
  wire \bdatw[12]_INST_0_i_32_n_0 ;
  wire \bdatw[13]_INST_0_i_16 ;
  wire \bdatw[13]_INST_0_i_16_0 ;
  wire \bdatw[13]_INST_0_i_16_1 ;
  wire \bdatw[13]_INST_0_i_16_2 ;
  wire \bdatw[13]_INST_0_i_2 ;
  wire \bdatw[13]_INST_0_i_2_0 ;
  wire \bdatw[13]_INST_0_i_2_1 ;
  wire \bdatw[13]_INST_0_i_2_2 ;
  wire \bdatw[13]_INST_0_i_34_n_0 ;
  wire \bdatw[13]_INST_0_i_63_n_0 ;
  wire \bdatw[14]_INST_0_i_16 ;
  wire \bdatw[14]_INST_0_i_16_0 ;
  wire \bdatw[14]_INST_0_i_16_1 ;
  wire \bdatw[14]_INST_0_i_16_2 ;
  wire \bdatw[14]_INST_0_i_2 ;
  wire \bdatw[14]_INST_0_i_2_0 ;
  wire \bdatw[14]_INST_0_i_2_1 ;
  wire \bdatw[14]_INST_0_i_2_2 ;
  wire \bdatw[14]_INST_0_i_39_n_0 ;
  wire \bdatw[14]_INST_0_i_82_n_0 ;
  wire \bdatw[15]_INST_0_i_134_n_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_15_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_15_1 ;
  wire \bdatw[15]_INST_0_i_16 ;
  wire \bdatw[15]_INST_0_i_16_0 ;
  wire \bdatw[15]_INST_0_i_16_1 ;
  wire \bdatw[15]_INST_0_i_16_2 ;
  wire \bdatw[15]_INST_0_i_2 ;
  wire \bdatw[15]_INST_0_i_2_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_2_1 ;
  wire \bdatw[15]_INST_0_i_2_2 ;
  wire \bdatw[15]_INST_0_i_2_3 ;
  wire [0:0]\bdatw[15]_INST_0_i_2_4 ;
  wire \bdatw[15]_INST_0_i_47_n_0 ;
  wire \bdatw[8]_INST_0_i_16 ;
  wire \bdatw[8]_INST_0_i_16_0 ;
  wire \bdatw[8]_INST_0_i_16_1 ;
  wire \bdatw[8]_INST_0_i_16_2 ;
  wire \bdatw[8]_INST_0_i_16_3 ;
  wire \bdatw[8]_INST_0_i_2 ;
  wire \bdatw[8]_INST_0_i_2_0 ;
  wire \bdatw[8]_INST_0_i_2_1 ;
  wire \bdatw[8]_INST_0_i_2_2 ;
  wire \bdatw[8]_INST_0_i_33_n_0 ;
  wire \bdatw[9]_INST_0_i_16 ;
  wire \bdatw[9]_INST_0_i_16_0 ;
  wire \bdatw[9]_INST_0_i_16_1 ;
  wire \bdatw[9]_INST_0_i_16_2 ;
  wire \bdatw[9]_INST_0_i_16_3 ;
  wire \bdatw[9]_INST_0_i_2 ;
  wire \bdatw[9]_INST_0_i_2_0 ;
  wire \bdatw[9]_INST_0_i_2_1 ;
  wire \bdatw[9]_INST_0_i_2_2 ;
  wire \bdatw[9]_INST_0_i_33_n_0 ;
  wire [14:0]data3;
  wire \iv_reg[15] ;
  wire [15:0]out;
  wire \sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[1] ;
  wire \sp_reg[2] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr_reg[0] ;
  wire \sr_reg[15] ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \tr_reg[0] ;
  wire \tr_reg[10] ;
  wire \tr_reg[11] ;
  wire \tr_reg[12] ;
  wire \tr_reg[13] ;
  wire \tr_reg[14] ;
  wire \tr_reg[1] ;
  wire \tr_reg[2] ;
  wire \tr_reg[3] ;
  wire \tr_reg[4] ;
  wire \tr_reg[5] ;
  wire \tr_reg[6] ;
  wire \tr_reg[7] ;
  wire \tr_reg[8] ;
  wire \tr_reg[9] ;

  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[10]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_2_1 [10]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[10]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[10]_INST_0_i_15 
       (.I0(\bdatw[10]_INST_0_i_34_n_0 ),
        .I1(\bdatw[10]_INST_0_i_2 ),
        .I2(\bdatw[10]_INST_0_i_2_0 ),
        .I3(\bdatw[10]_INST_0_i_2_1 ),
        .I4(\bdatw[10]_INST_0_i_2_2 ),
        .I5(b1bus_sr[10]),
        .O(\sp_reg[10] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_34 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[9]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [10]),
        .I4(\bdatw[15]_INST_0_i_15_1 [10]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[10]_INST_0_i_41 
       (.I0(\bdatw[15]_INST_0_i_2_1 [2]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[2]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[10]_INST_0_i_43 
       (.I0(b1bus_sr[2]),
        .I1(\bdatw[10]_INST_0_i_16 ),
        .I2(\bdatw[10]_INST_0_i_16_0 ),
        .I3(\bdatw[10]_INST_0_i_16_1 ),
        .I4(\bdatw[10]_INST_0_i_16_2 ),
        .I5(\bdatw[10]_INST_0_i_16_3 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_44 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[1]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [2]),
        .I4(\bdatw[15]_INST_0_i_15_1 [2]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[11]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_2_1 [11]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[11]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[11]_INST_0_i_15 
       (.I0(\bdatw[11]_INST_0_i_34_n_0 ),
        .I1(\bdatw[11]_INST_0_i_2 ),
        .I2(\bdatw[11]_INST_0_i_2_0 ),
        .I3(\bdatw[11]_INST_0_i_2_1 ),
        .I4(\bdatw[11]_INST_0_i_2_2 ),
        .I5(b1bus_sr[11]),
        .O(\sp_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_34 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[10]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [11]),
        .I4(\bdatw[15]_INST_0_i_15_1 [11]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[11]_INST_0_i_42 
       (.I0(\bdatw[15]_INST_0_i_2_1 [3]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[3]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[11]_INST_0_i_44 
       (.I0(b1bus_sr[3]),
        .I1(\bdatw[11]_INST_0_i_16 ),
        .I2(\bdatw[11]_INST_0_i_16_0 ),
        .I3(\bdatw[11]_INST_0_i_16_1 ),
        .I4(\bdatw[11]_INST_0_i_16_2 ),
        .I5(\bdatw[11]_INST_0_i_16_3 ),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_45 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[2]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [3]),
        .I4(\bdatw[15]_INST_0_i_15_1 [3]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[3] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[12]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_2_1 [12]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[12]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[12]_INST_0_i_15 
       (.I0(\bdatw[12]_INST_0_i_32_n_0 ),
        .I1(\bdatw[12]_INST_0_i_2 ),
        .I2(\bdatw[12]_INST_0_i_2_0 ),
        .I3(\bdatw[12]_INST_0_i_2_1 ),
        .I4(\bdatw[12]_INST_0_i_2_2 ),
        .I5(b1bus_sr[12]),
        .O(\sp_reg[12] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_32 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[11]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [12]),
        .I4(\bdatw[15]_INST_0_i_15_1 [12]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[12]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[12]_INST_0_i_40 
       (.I0(\bdatw[15]_INST_0_i_2_1 [4]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[4]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[12]_INST_0_i_42 
       (.I0(b1bus_sr[4]),
        .I1(\bdatw[12]_INST_0_i_16 ),
        .I2(\bdatw[12]_INST_0_i_16_0 ),
        .I3(\bdatw[12]_INST_0_i_16_1 ),
        .I4(\bdatw[12]_INST_0_i_16_2 ),
        .I5(\bdatw[12]_INST_0_i_16_3 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_43 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[3]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [4]),
        .I4(\bdatw[15]_INST_0_i_15_1 [4]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[13]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_2_1 [13]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[13]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_15 
       (.I0(\bdatw[13]_INST_0_i_34_n_0 ),
        .I1(\bdatw[13]_INST_0_i_2 ),
        .I2(\bdatw[13]_INST_0_i_2_0 ),
        .I3(\bdatw[13]_INST_0_i_2_1 ),
        .I4(\bdatw[13]_INST_0_i_2_2 ),
        .I5(b1bus_sr[13]),
        .O(\sp_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_34 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[12]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [13]),
        .I4(\bdatw[15]_INST_0_i_15_1 [13]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[13]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[13]_INST_0_i_42 
       (.I0(\bdatw[15]_INST_0_i_2_1 [5]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[5]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_45 
       (.I0(\bdatw[13]_INST_0_i_63_n_0 ),
        .I1(\bdatw[13]_INST_0_i_16 ),
        .I2(\bdatw[13]_INST_0_i_16_0 ),
        .I3(\bdatw[13]_INST_0_i_16_1 ),
        .I4(\bdatw[13]_INST_0_i_16_2 ),
        .I5(b1bus_sr[5]),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_63 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[4]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [5]),
        .I4(\bdatw[15]_INST_0_i_15_1 [5]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[13]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[14]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_2_1 [14]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[14]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[14]_INST_0_i_15 
       (.I0(\bdatw[14]_INST_0_i_39_n_0 ),
        .I1(\bdatw[14]_INST_0_i_2 ),
        .I2(\bdatw[14]_INST_0_i_2_0 ),
        .I3(\bdatw[14]_INST_0_i_2_1 ),
        .I4(\bdatw[14]_INST_0_i_2_2 ),
        .I5(b1bus_sr[14]),
        .O(\sp_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_39 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[13]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [14]),
        .I4(\bdatw[15]_INST_0_i_15_1 [14]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[14]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[14]_INST_0_i_47 
       (.I0(\bdatw[15]_INST_0_i_2_1 [6]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[6]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[14]_INST_0_i_50 
       (.I0(\bdatw[14]_INST_0_i_82_n_0 ),
        .I1(\bdatw[14]_INST_0_i_16 ),
        .I2(\bdatw[14]_INST_0_i_16_0 ),
        .I3(\bdatw[14]_INST_0_i_16_1 ),
        .I4(\bdatw[14]_INST_0_i_16_2 ),
        .I5(b1bus_sr[6]),
        .O(\sp_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_82 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[5]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [6]),
        .I4(\bdatw[15]_INST_0_i_15_1 [6]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[14]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_134 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[6]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [7]),
        .I4(\bdatw[15]_INST_0_i_15_1 [7]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[15]_INST_0_i_134_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[15]_INST_0_i_14 
       (.I0(\bdatw[15]_INST_0_i_2 ),
        .I1(\bdatw[15]_INST_0_i_2_0 ),
        .I2(b1bus_sel_cr[3]),
        .I3(out[15]),
        .I4(b1bus_sel_cr[4]),
        .I5(\bdatw[15]_INST_0_i_2_1 [15]),
        .O(\iv_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[15]_INST_0_i_15 
       (.I0(\bdatw[15]_INST_0_i_47_n_0 ),
        .I1(\bdatw[15]_INST_0_i_2_2 ),
        .I2(\bdatw[15]_INST_0_i_2_3 ),
        .I3(b1bus_sel_cr[0]),
        .I4(\bdatw[15]_INST_0_i_2_4 ),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_47 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[14]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [15]),
        .I4(\bdatw[15]_INST_0_i_15_1 [15]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[15]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[15]_INST_0_i_53 
       (.I0(\bdatw[15]_INST_0_i_2_1 [7]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[7]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_56 
       (.I0(\bdatw[15]_INST_0_i_134_n_0 ),
        .I1(\bdatw[15]_INST_0_i_16 ),
        .I2(\bdatw[15]_INST_0_i_16_0 ),
        .I3(\bdatw[15]_INST_0_i_16_1 ),
        .I4(\bdatw[15]_INST_0_i_16_2 ),
        .I5(b1bus_sr[7]),
        .O(\sp_reg[7] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[8]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_2_1 [8]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[8]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_15 
       (.I0(\bdatw[8]_INST_0_i_33_n_0 ),
        .I1(\bdatw[8]_INST_0_i_2 ),
        .I2(\bdatw[8]_INST_0_i_2_0 ),
        .I3(\bdatw[8]_INST_0_i_2_1 ),
        .I4(\bdatw[8]_INST_0_i_2_2 ),
        .I5(b1bus_sr[8]),
        .O(\sp_reg[8] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_33 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[7]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [8]),
        .I4(\bdatw[15]_INST_0_i_15_1 [8]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[8]_INST_0_i_41 
       (.I0(\bdatw[15]_INST_0_i_2_1 [0]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[0]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_43 
       (.I0(b1bus_sr[0]),
        .I1(\bdatw[8]_INST_0_i_16 ),
        .I2(\bdatw[8]_INST_0_i_16_0 ),
        .I3(\bdatw[8]_INST_0_i_16_1 ),
        .I4(\bdatw[8]_INST_0_i_16_2 ),
        .I5(\bdatw[8]_INST_0_i_16_3 ),
        .O(\sr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_44 
       (.I0(b1bus_sel_cr[5]),
        .I1(O),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [0]),
        .I4(\bdatw[15]_INST_0_i_15_1 [0]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[9]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_2_1 [9]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[9]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[9]_INST_0_i_15 
       (.I0(\bdatw[9]_INST_0_i_33_n_0 ),
        .I1(\bdatw[9]_INST_0_i_2 ),
        .I2(\bdatw[9]_INST_0_i_2_0 ),
        .I3(\bdatw[9]_INST_0_i_2_1 ),
        .I4(\bdatw[9]_INST_0_i_2_2 ),
        .I5(b1bus_sr[9]),
        .O(\sp_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_33 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[8]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [9]),
        .I4(\bdatw[15]_INST_0_i_15_1 [9]),
        .I5(b1bus_sel_cr[1]),
        .O(\bdatw[9]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[9]_INST_0_i_40 
       (.I0(\bdatw[15]_INST_0_i_2_1 [1]),
        .I1(b1bus_sel_cr[4]),
        .I2(out[1]),
        .I3(b1bus_sel_cr[3]),
        .O(\tr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[9]_INST_0_i_42 
       (.I0(b1bus_sr[1]),
        .I1(\bdatw[9]_INST_0_i_16 ),
        .I2(\bdatw[9]_INST_0_i_16_0 ),
        .I3(\bdatw[9]_INST_0_i_16_1 ),
        .I4(\bdatw[9]_INST_0_i_16_2 ),
        .I5(\bdatw[9]_INST_0_i_16_3 ),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_43 
       (.I0(b1bus_sel_cr[5]),
        .I1(data3[0]),
        .I2(b1bus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_15_0 [1]),
        .I4(\bdatw[15]_INST_0_i_15_1 [1]),
        .I5(b1bus_sel_cr[1]),
        .O(\sp_reg[1] ));
endmodule

module mcss_rgf_ctl
   (rgf_selc0_stat,
    rgf_selc1_stat,
    bank_sel,
    \sr_reg[0] ,
    \rgf_selc0_rn_wb_reg[2]_0 ,
    \rgf_selc0_wb_reg[1]_0 ,
    \rgf_selc1_rn_wb_reg[2]_0 ,
    \rgf_selc1_wb_reg[1]_0 ,
    \rgf_c0bus_wb_reg[15]_0 ,
    \rgf_c1bus_wb_reg[15]_0 ,
    E,
    p_2_in,
    clk,
    \rgf_selc1_wb_reg[0]_0 ,
    rgf_selc1_stat_reg_0,
    \rgf_c1bus_wb_reg[0]_0 ,
    rst_n,
    out,
    \rgf_selc0_rn_wb_reg[2]_1 ,
    \rgf_selc0_wb_reg[1]_1 ,
    \rgf_selc1_rn_wb_reg[2]_1 ,
    \rgf_selc1_wb_reg[1]_1 ,
    \rgf_c0bus_wb_reg[15]_1 ,
    \rgf_c1bus_wb_reg[15]_1 );
  output rgf_selc0_stat;
  output rgf_selc1_stat;
  output [0:0]bank_sel;
  output [0:0]\sr_reg[0] ;
  output [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc0_wb_reg[1]_0 ;
  output [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  output [1:0]\rgf_selc1_wb_reg[1]_0 ;
  output [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  output [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  input [0:0]E;
  input p_2_in;
  input clk;
  input [0:0]\rgf_selc1_wb_reg[0]_0 ;
  input rgf_selc1_stat_reg_0;
  input \rgf_c1bus_wb_reg[0]_0 ;
  input rst_n;
  input [1:0]out;
  input [2:0]\rgf_selc0_rn_wb_reg[2]_1 ;
  input [1:0]\rgf_selc0_wb_reg[1]_1 ;
  input [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  input [1:0]\rgf_selc1_wb_reg[1]_1 ;
  input [15:0]\rgf_c0bus_wb_reg[15]_1 ;
  input [15:0]\rgf_c1bus_wb_reg[15]_1 ;

  wire [0:0]E;
  wire [0:0]bank_sel;
  wire clk;
  wire [1:0]out;
  wire p_2_in;
  wire [15:0]\rgf_c0bus_wb_reg[15]_0 ;
  wire [15:0]\rgf_c0bus_wb_reg[15]_1 ;
  wire \rgf_c1bus_wb_reg[0]_0 ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_0 ;
  wire [15:0]\rgf_c1bus_wb_reg[15]_1 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_0 ;
  wire [2:0]\rgf_selc0_rn_wb_reg[2]_1 ;
  wire rgf_selc0_stat;
  wire rgf_selc0_stat_i_1_n_0;
  wire [1:0]\rgf_selc0_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc0_wb_reg[1]_1 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_0 ;
  wire [2:0]\rgf_selc1_rn_wb_reg[2]_1 ;
  wire rgf_selc1_stat;
  wire rgf_selc1_stat_reg_0;
  wire [0:0]\rgf_selc1_wb_reg[0]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_0 ;
  wire [1:0]\rgf_selc1_wb_reg[1]_1 ;
  wire rst_n;
  wire [0:0]\sr_reg[0] ;

  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_186 
       (.I0(out[0]),
        .I1(out[1]),
        .O(\sr_reg[0] ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[15]_INST_0_i_74 
       (.I0(out[0]),
        .I1(out[1]),
        .O(bank_sel));
  FDRE \rgf_c0bus_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [0]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[10] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [10]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[11] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [11]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[12] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [12]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[13] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [13]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[14] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [14]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[15] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [15]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [1]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [2]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[3] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [3]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[4] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [4]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[5] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [5]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[6] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [6]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[7] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [7]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[8] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [8]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c0bus_wb_reg[9] 
       (.C(clk),
        .CE(E),
        .D(\rgf_c0bus_wb_reg[15]_1 [9]),
        .Q(\rgf_c0bus_wb_reg[15]_0 [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [0]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[10] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [10]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[11] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [11]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[12] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [12]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[13] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [13]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[14] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [14]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[15] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [15]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [1]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [2]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[3] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [3]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[4] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [4]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[5] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [5]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[6] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [6]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[7] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [7]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[8] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [8]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_c1bus_wb_reg[9] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_c1bus_wb_reg[15]_1 [9]),
        .Q(\rgf_c1bus_wb_reg[15]_0 [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [0]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [1]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_rn_wb_reg[2] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_rn_wb_reg[2]_1 [2]),
        .Q(\rgf_selc0_rn_wb_reg[2]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    rgf_selc0_stat_i_1
       (.I0(\rgf_c1bus_wb_reg[0]_0 ),
        .I1(rst_n),
        .O(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc0_stat_reg
       (.C(clk),
        .CE(E),
        .D(p_2_in),
        .Q(rgf_selc0_stat),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[0] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [0]),
        .Q(\rgf_selc0_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc0_wb_reg[1] 
       (.C(clk),
        .CE(E),
        .D(\rgf_selc0_wb_reg[1]_1 [1]),
        .Q(\rgf_selc0_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [0]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [1]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_rn_wb_reg[2] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_rn_wb_reg[2]_1 [2]),
        .Q(\rgf_selc1_rn_wb_reg[2]_0 [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE rgf_selc1_stat_reg
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(rgf_selc1_stat_reg_0),
        .Q(rgf_selc1_stat),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[0] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [0]),
        .Q(\rgf_selc1_wb_reg[1]_0 [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf_selc1_wb_reg[1] 
       (.C(clk),
        .CE(\rgf_selc1_wb_reg[0]_0 ),
        .D(\rgf_selc1_wb_reg[1]_1 [1]),
        .Q(\rgf_selc1_wb_reg[1]_0 [1]),
        .R(rgf_selc0_stat_i_1_n_0));
endmodule

module mcss_rgf_grn
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_13
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_14
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_15
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_16
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_17
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_18
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_19
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_20
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_21
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_22
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_23
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_24
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_25
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_26
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_27
   (SR,
    \rgf_c1bus_wb[14]_i_28 ,
    \tr_reg[1] ,
    \tr_reg[14] ,
    \fdatx[15] ,
    .fdat_12_sp_1(fdat_12_sn_1),
    \fdat[15] ,
    Q,
    rst_n,
    \rgf_c1bus_wb[4]_i_4 ,
    \rgf_c1bus_wb[4]_i_4_0 ,
    \rgf_c1bus_wb[4]_i_4_1 ,
    \rgf_c1bus_wb[4]_i_4_2 ,
    \rgf_c1bus_wb[4]_i_4_3 ,
    \rgf_c1bus_wb[4]_i_4_4 ,
    \rgf_c1bus_wb[4]_i_13 ,
    \rgf_c1bus_wb[4]_i_11 ,
    \rgf_c1bus_wb[4]_i_13_0 ,
    \rgf_c1bus_wb[4]_i_11_0 ,
    \rgf_c1bus_wb[4]_i_13_1 ,
    \rgf_c1bus_wb[4]_i_13_2 ,
    \rgf_c1bus_wb[4]_i_11_1 ,
    \rgf_c1bus_wb[4]_i_11_2 ,
    \rgf_c1bus_wb[4]_i_11_3 ,
    \rgf_c1bus_wb[4]_i_11_4 ,
    fdatx,
    \ir0_id_fl[20]_i_4_0 ,
    fdat,
    \nir_id_reg[20] ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [0:0]SR;
  output \rgf_c1bus_wb[14]_i_28 ;
  output \tr_reg[1] ;
  output \tr_reg[14] ;
  output \fdatx[15] ;
  output [0:0]\fdat[15] ;
  output [15:0]Q;
  input rst_n;
  input \rgf_c1bus_wb[4]_i_4 ;
  input \rgf_c1bus_wb[4]_i_4_0 ;
  input \rgf_c1bus_wb[4]_i_4_1 ;
  input \rgf_c1bus_wb[4]_i_4_2 ;
  input \rgf_c1bus_wb[4]_i_4_3 ;
  input \rgf_c1bus_wb[4]_i_4_4 ;
  input \rgf_c1bus_wb[4]_i_13 ;
  input [1:0]\rgf_c1bus_wb[4]_i_11 ;
  input \rgf_c1bus_wb[4]_i_13_0 ;
  input \rgf_c1bus_wb[4]_i_11_0 ;
  input \rgf_c1bus_wb[4]_i_13_1 ;
  input \rgf_c1bus_wb[4]_i_13_2 ;
  input \rgf_c1bus_wb[4]_i_11_1 ;
  input \rgf_c1bus_wb[4]_i_11_2 ;
  input \rgf_c1bus_wb[4]_i_11_3 ;
  input \rgf_c1bus_wb[4]_i_11_4 ;
  input [13:0]fdatx;
  input \ir0_id_fl[20]_i_4_0 ;
  input [13:0]fdat;
  input \nir_id_reg[20] ;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;
  output fdat_12_sn_1;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [13:0]fdat;
  wire [0:0]\fdat[15] ;
  wire fdat_12_sn_1;
  wire [13:0]fdatx;
  wire \fdatx[15] ;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire \ir0_id_fl[20]_i_4_0 ;
  wire \ir0_id_fl[20]_i_4_n_0 ;
  wire \ir0_id_fl[20]_i_5_n_0 ;
  wire \ir0_id_fl[20]_i_6_n_0 ;
  wire \ir0_id_fl[20]_i_7_n_0 ;
  wire \nir_id[20]_i_2_n_0 ;
  wire \nir_id[20]_i_3_n_0 ;
  wire \nir_id[20]_i_4_n_0 ;
  wire \nir_id_reg[20] ;
  wire \rgf_c1bus_wb[14]_i_28 ;
  wire [1:0]\rgf_c1bus_wb[4]_i_11 ;
  wire \rgf_c1bus_wb[4]_i_11_0 ;
  wire \rgf_c1bus_wb[4]_i_11_1 ;
  wire \rgf_c1bus_wb[4]_i_11_2 ;
  wire \rgf_c1bus_wb[4]_i_11_3 ;
  wire \rgf_c1bus_wb[4]_i_11_4 ;
  wire \rgf_c1bus_wb[4]_i_13 ;
  wire \rgf_c1bus_wb[4]_i_13_0 ;
  wire \rgf_c1bus_wb[4]_i_13_1 ;
  wire \rgf_c1bus_wb[4]_i_13_2 ;
  wire \rgf_c1bus_wb[4]_i_4 ;
  wire \rgf_c1bus_wb[4]_i_4_0 ;
  wire \rgf_c1bus_wb[4]_i_4_1 ;
  wire \rgf_c1bus_wb[4]_i_4_2 ;
  wire \rgf_c1bus_wb[4]_i_4_3 ;
  wire \rgf_c1bus_wb[4]_i_4_4 ;
  wire rst_n;
  wire \tr_reg[14] ;
  wire \tr_reg[1] ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT6 #(
    .INIT(64'hABAAABABABABABAB)) 
    \ir0_id_fl[20]_i_3 
       (.I0(fdatx[13]),
        .I1(\ir0_id_fl[20]_i_4_n_0 ),
        .I2(\ir0_id_fl[20]_i_5_n_0 ),
        .I3(\ir0_id_fl[20]_i_6_n_0 ),
        .I4(fdatx[10]),
        .I5(fdatx[8]),
        .O(\fdatx[15] ));
  LUT6 #(
    .INIT(64'h0000000301020002)) 
    \ir0_id_fl[20]_i_4 
       (.I0(fdatx[1]),
        .I1(\ir0_id_fl[20]_i_7_n_0 ),
        .I2(fdatx[11]),
        .I3(fdatx[3]),
        .I4(fdatx[2]),
        .I5(fdatx[0]),
        .O(\ir0_id_fl[20]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h7776)) 
    \ir0_id_fl[20]_i_5 
       (.I0(fdatx[11]),
        .I1(fdatx[12]),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .O(\ir0_id_fl[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hA2AABBBBFFFFAAAA)) 
    \ir0_id_fl[20]_i_6 
       (.I0(fdatx[7]),
        .I1(fdatx[5]),
        .I2(fdatx[4]),
        .I3(\ir0_id_fl[20]_i_4_0 ),
        .I4(fdatx[6]),
        .I5(fdatx[9]),
        .O(\ir0_id_fl[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \ir0_id_fl[20]_i_7 
       (.I0(\ir0_id_fl[20]_i_4_0 ),
        .I1(fdatx[6]),
        .I2(fdatx[7]),
        .I3(fdatx[8]),
        .I4(fdatx[4]),
        .I5(fdatx[5]),
        .O(\ir0_id_fl[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5455545454545454)) 
    \nir_id[20]_i_1 
       (.I0(fdat[13]),
        .I1(fdat_12_sn_1),
        .I2(\nir_id[20]_i_2_n_0 ),
        .I3(\nir_id[20]_i_3_n_0 ),
        .I4(fdat[10]),
        .I5(fdat[8]),
        .O(\fdat[15] ));
  LUT6 #(
    .INIT(64'h0000000301020002)) 
    \nir_id[20]_i_2 
       (.I0(fdat[1]),
        .I1(\nir_id[20]_i_4_n_0 ),
        .I2(fdat[11]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[0]),
        .O(\nir_id[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA2AABBBBFFFFAAAA)) 
    \nir_id[20]_i_3 
       (.I0(fdat[7]),
        .I1(fdat[5]),
        .I2(fdat[4]),
        .I3(\nir_id_reg[20] ),
        .I4(fdat[6]),
        .I5(fdat[9]),
        .O(\nir_id[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \nir_id[20]_i_4 
       (.I0(fdat[8]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[6]),
        .I4(fdat[7]),
        .I5(\nir_id_reg[20] ),
        .O(\nir_id[20]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0FFE)) 
    \nir_id[24]_i_9 
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .I2(fdat[11]),
        .I3(fdat[12]),
        .O(fdat_12_sn_1));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \rgf_c1bus_wb[4]_i_12 
       (.I0(\rgf_c1bus_wb[4]_i_4 ),
        .I1(\rgf_c1bus_wb[4]_i_4_0 ),
        .I2(\rgf_c1bus_wb[4]_i_4_1 ),
        .I3(\rgf_c1bus_wb[4]_i_4_2 ),
        .I4(\rgf_c1bus_wb[4]_i_4_3 ),
        .I5(\rgf_c1bus_wb[4]_i_4_4 ),
        .O(\rgf_c1bus_wb[14]_i_28 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_23 
       (.I0(\rgf_c1bus_wb[4]_i_11_1 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [1]),
        .I2(\rgf_c1bus_wb[4]_i_11_2 ),
        .I3(\rgf_c1bus_wb[4]_i_11_0 ),
        .I4(\rgf_c1bus_wb[4]_i_11_3 ),
        .I5(\rgf_c1bus_wb[4]_i_11_4 ),
        .O(\tr_reg[14] ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_29 
       (.I0(\rgf_c1bus_wb[4]_i_13 ),
        .I1(\rgf_c1bus_wb[4]_i_11 [0]),
        .I2(\rgf_c1bus_wb[4]_i_13_0 ),
        .I3(\rgf_c1bus_wb[4]_i_11_0 ),
        .I4(\rgf_c1bus_wb[4]_i_13_1 ),
        .I5(\rgf_c1bus_wb[4]_i_13_2 ),
        .O(\tr_reg[1] ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1 
       (.I0(rst_n),
        .O(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_36
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_37
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_38
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_39
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_40
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_41
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_42
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_43
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_44
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_45
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_46
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_47
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_48
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_49
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_50
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "mcss_rgf_grn" *) 
module mcss_rgf_grn_51
   (\stat_reg[2] ,
    \tr_reg[6] ,
    \badr[6]_INST_0_i_1 ,
    \stat_reg[2]_0 ,
    \tr_reg[5] ,
    \badr[5]_INST_0_i_1 ,
    \rgf_c1bus_wb[13]_i_9_0 ,
    \rgf_c1bus_wb[14]_i_30_0 ,
    \sr_reg[6] ,
    \badr[15]_INST_0_i_1 ,
    \badr[15]_INST_0_i_1_0 ,
    \sr_reg[6]_0 ,
    \badr[9]_INST_0_i_1 ,
    \sr_reg[6]_1 ,
    \rgf_c1bus_wb[11]_i_13_0 ,
    \badr[14]_INST_0_i_1 ,
    \sr_reg[6]_2 ,
    \rgf_c1bus_wb[12]_i_20 ,
    \rgf_c1bus_wb[11]_i_10 ,
    \rgf_c1bus_wb[14]_i_28 ,
    \rgf_c1bus_wb[7]_i_4 ,
    \badr[5]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[4]_i_9_0 ,
    \badr[12]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_28_0 ,
    \badr[0]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_28_1 ,
    \sr_reg[6]_3 ,
    \badr[3]_INST_0_i_1 ,
    \rgf_c1bus_wb[9]_i_17 ,
    \badr[10]_INST_0_i_1 ,
    \rgf_c1bus_wb[13]_i_16_0 ,
    \rgf_c1bus_wb[14]_i_28_2 ,
    \sr_reg[6]_4 ,
    \sr_reg[6]_5 ,
    \sr_reg[6]_6 ,
    \sr_reg[6]_7 ,
    \rgf_c1bus_wb[15]_i_14 ,
    \rgf_c1bus_wb[14]_i_28_3 ,
    \badr[9]_INST_0_i_1_0 ,
    \rgf_c1bus_wb[14]_i_32_0 ,
    \badr[13]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \rgf_c1bus_wb[14]_i_32_1 ,
    \sr_reg[6]_8 ,
    \badr[14]_INST_0_i_1_0 ,
    \sr_reg[6]_9 ,
    \rgf_c1bus_wb[1]_i_14 ,
    \sr_reg[6]_10 ,
    \badr[11]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1_0 ,
    \badr[2]_INST_0_i_1_0 ,
    \badr[10]_INST_0_i_1_0 ,
    \stat_reg[2]_1 ,
    \stat_reg[2]_2 ,
    \rgf_c0bus_wb[15]_i_18_0 ,
    \rgf_c0bus_wb[11]_i_3 ,
    \tr_reg[7] ,
    \rgf_c0bus_wb[11]_i_3_0 ,
    \badr[6]_INST_0_i_2 ,
    \tr_reg[6]_0 ,
    \tr_reg[5]_0 ,
    \sr_reg[6]_11 ,
    \sr_reg[6]_12 ,
    \badr[10]_INST_0_i_2 ,
    \badr[14]_INST_0_i_2 ,
    \rgf_c0bus_wb[13]_i_29_0 ,
    \badr[4]_INST_0_i_2 ,
    \badr[12]_INST_0_i_2 ,
    \badr[8]_INST_0_i_2 ,
    \rgf_c0bus_wb[7]_i_7 ,
    \badr[6]_INST_0_i_2_0 ,
    \badr[10]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[7]_i_7_0 ,
    \sr_reg[6]_13 ,
    \sr_reg[6]_14 ,
    \badr[14]_INST_0_i_2_0 ,
    \badr[1]_INST_0_i_2 ,
    \sr_reg[6]_15 ,
    \rgf_c0bus_wb[15]_i_26_0 ,
    \sr_reg[6]_16 ,
    \badr[3]_INST_0_i_2 ,
    \badr[11]_INST_0_i_2 ,
    \badr[7]_INST_0_i_2 ,
    \rgf_c0bus_wb[11]_i_22 ,
    \badr[6]_INST_0_i_2_1 ,
    \badr[2]_INST_0_i_2 ,
    \sr_reg[6]_17 ,
    \sr_reg[6]_18 ,
    \sr_reg[6]_19 ,
    \rgf_c0bus_wb[10]_i_8_0 ,
    \badr[5]_INST_0_i_2 ,
    \badr[5]_INST_0_i_2_0 ,
    \badr[1]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[11]_i_9 ,
    \rgf_c0bus_wb[13]_i_28_0 ,
    \badr[14]_INST_0_i_2_1 ,
    \sr_reg[6]_20 ,
    \sr_reg[6]_21 ,
    \badr[12]_INST_0_i_2_0 ,
    \rgf_c0bus_wb[11]_i_3_1 ,
    \rgf_c1bus_wb[7]_i_4_0 ,
    \sr_reg[6]_22 ,
    \rgf_c0bus_wb[15]_i_6 ,
    \rgf_c0bus_wb[15]_i_6_0 ,
    \rgf_c0bus_wb[15]_i_6_1 ,
    \rgf_c0bus_wb[11]_i_9_0 ,
    \rgf_c0bus_wb[11]_i_9_1 ,
    \rgf_c0bus_wb[11]_i_9_2 ,
    \rgf_c0bus_wb[11]_i_3_2 ,
    Q,
    \rgf_c1bus_wb[2]_i_7 ,
    \rgf_c1bus_wb_reg[5] ,
    \rgf_c1bus_wb[10]_i_14 ,
    \rgf_c1bus_wb[14]_i_3 ,
    \rgf_c1bus_wb[5]_i_10 ,
    \rgf_c1bus_wb[14]_i_11 ,
    \rgf_c1bus_wb[14]_i_11_0 ,
    \rgf_c1bus_wb[14]_i_11_1 ,
    \rgf_c1bus_wb[14]_i_11_2 ,
    \rgf_c1bus_wb[14]_i_11_3 ,
    \rgf_c1bus_wb[14]_i_11_4 ,
    \rgf_c1bus_wb[11]_i_11 ,
    \rgf_c1bus_wb[2]_i_7_0 ,
    tout__1_carry__0_i_7__0,
    tout__1_carry__0_i_7__0_0,
    tout__1_carry__0_i_7__0_1,
    tout__1_carry__0_i_7__0_2,
    tout__1_carry__0_i_7__0_3,
    tout__1_carry__0_i_7__0_4,
    \rgf_c1bus_wb_reg[5]_0 ,
    \rgf_c1bus_wb_reg[5]_1 ,
    \rgf_c1bus_wb[4]_i_7_0 ,
    \rgf_c1bus_wb[11]_i_11_0 ,
    \rgf_c1bus_wb_reg[7] ,
    \rgf_c1bus_wb[2]_i_7_1 ,
    \rgf_c0bus_wb[3]_i_7 ,
    \rgf_c1bus_wb[3]_i_4 ,
    \rgf_c1bus_wb[11]_i_11_1 ,
    \rgf_c1bus_wb[2]_i_7_2 ,
    \rgf_c1bus_wb[3]_i_4_0 ,
    \rgf_c1bus_wb[8]_i_3 ,
    \rgf_c1bus_wb_reg[3] ,
    \rgf_c1bus_wb[8]_i_3_0 ,
    \rgf_c1bus_wb[11]_i_11_2 ,
    \rgf_c1bus_wb[11]_i_11_3 ,
    \rgf_c1bus_wb[11]_i_11_4 ,
    \rgf_c1bus_wb[11]_i_11_5 ,
    \rgf_c1bus_wb_reg[4] ,
    \rgf_c1bus_wb[4]_i_3_0 ,
    \rgf_c1bus_wb[4]_i_3_1 ,
    \rgf_c1bus_wb[4]_i_3_2 ,
    \rgf_c1bus_wb[12]_i_2 ,
    \rgf_c1bus_wb[12]_i_2_0 ,
    \rgf_c1bus_wb[11]_i_8 ,
    \rgf_c1bus_wb[11]_i_11_6 ,
    \rgf_c1bus_wb[11]_i_8_0 ,
    \rgf_c1bus_wb[10]_i_14_0 ,
    \rgf_c1bus_wb[11]_i_8_1 ,
    \rgf_c1bus_wb[1]_i_3 ,
    \rgf_c1bus_wb_reg[1] ,
    \rgf_c1bus_wb_reg[10] ,
    \rgf_c1bus_wb_reg[1]_0 ,
    \rgf_c1bus_wb[4]_i_7_1 ,
    \rgf_c1bus_wb[4]_i_7_2 ,
    \rgf_c1bus_wb[4]_i_7_3 ,
    \rgf_c1bus_wb[4]_i_7_4 ,
    \rgf_c1bus_wb[4]_i_7_5 ,
    \rgf_c0bus_wb_reg[7]_i_11 ,
    \rgf_c0bus_wb[1]_i_3 ,
    \rgf_c0bus_wb[6]_i_11 ,
    \rgf_c0bus_wb[7]_i_15_0 ,
    \rgf_c0bus_wb[5]_i_8 ,
    \rgf_c0bus_wb[11]_i_17 ,
    \rgf_c0bus_wb[10]_i_26 ,
    \bbus_o[7] ,
    \bbus_o[7]_0 ,
    \bbus_o[7]_1 ,
    p_1_in3_in,
    p_0_in2_in,
    \bbus_o[7]_2 ,
    \sr[4]_i_144 ,
    \bbus_o[6] ,
    \bbus_o[6]_0 ,
    \bbus_o[6]_1 ,
    \bbus_o[6]_2 ,
    \bbus_o[5] ,
    \bbus_o[5]_0 ,
    \bbus_o[5]_1 ,
    \bbus_o[5]_2 ,
    \rgf_c0bus_wb_reg[10] ,
    \rgf_c0bus_wb_reg[10]_0 ,
    \rgf_c0bus_wb[13]_i_4 ,
    \rgf_c0bus_wb[10]_i_4 ,
    \rgf_c0bus_wb[5]_i_2 ,
    \sr[4]_i_56 ,
    \rgf_c0bus_wb_reg[10]_1 ,
    \sr[4]_i_144_0 ,
    \sr[4]_i_144_1 ,
    \rgf_c0bus_wb[11]_i_17_0 ,
    \rgf_c0bus_wb[11]_i_17_1 ,
    \rgf_c0bus_wb[10]_i_26_0 ,
    \rgf_c0bus_wb[11]_i_17_2 ,
    \rgf_c0bus_wb[11]_i_17_3 ,
    \rgf_c0bus_wb[7]_i_15_1 ,
    \rgf_c0bus_wb[11]_i_17_4 ,
    \rgf_c0bus_wb[5]_i_8_0 ,
    \rgf_c0bus_wb[5]_i_8_1 ,
    \rgf_c0bus_wb[0]_i_8 ,
    \rgf_c0bus_wb[5]_i_8_2 ,
    \rgf_c0bus_wb[10]_i_26_1 ,
    \rgf_c0bus_wb[4]_i_3 ,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output \stat_reg[2] ;
  output \tr_reg[6] ;
  output \badr[6]_INST_0_i_1 ;
  output \stat_reg[2]_0 ;
  output \tr_reg[5] ;
  output \badr[5]_INST_0_i_1 ;
  output \rgf_c1bus_wb[13]_i_9_0 ;
  output \rgf_c1bus_wb[14]_i_30_0 ;
  output \sr_reg[6] ;
  output \badr[15]_INST_0_i_1 ;
  output \badr[15]_INST_0_i_1_0 ;
  output \sr_reg[6]_0 ;
  output \badr[9]_INST_0_i_1 ;
  output \sr_reg[6]_1 ;
  output \rgf_c1bus_wb[11]_i_13_0 ;
  output \badr[14]_INST_0_i_1 ;
  output \sr_reg[6]_2 ;
  output \rgf_c1bus_wb[12]_i_20 ;
  output \rgf_c1bus_wb[11]_i_10 ;
  output \rgf_c1bus_wb[14]_i_28 ;
  output \rgf_c1bus_wb[7]_i_4 ;
  output \badr[5]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[4]_i_9_0 ;
  output \badr[12]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_28_0 ;
  output \badr[0]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_28_1 ;
  output \sr_reg[6]_3 ;
  output \badr[3]_INST_0_i_1 ;
  output \rgf_c1bus_wb[9]_i_17 ;
  output \badr[10]_INST_0_i_1 ;
  output \rgf_c1bus_wb[13]_i_16_0 ;
  output \rgf_c1bus_wb[14]_i_28_2 ;
  output \sr_reg[6]_4 ;
  output \sr_reg[6]_5 ;
  output \sr_reg[6]_6 ;
  output \sr_reg[6]_7 ;
  output \rgf_c1bus_wb[15]_i_14 ;
  output \rgf_c1bus_wb[14]_i_28_3 ;
  output \badr[9]_INST_0_i_1_0 ;
  output \rgf_c1bus_wb[14]_i_32_0 ;
  output \badr[13]_INST_0_i_1 ;
  output \badr[2]_INST_0_i_1 ;
  output \rgf_c1bus_wb[14]_i_32_1 ;
  output \sr_reg[6]_8 ;
  output \badr[14]_INST_0_i_1_0 ;
  output \sr_reg[6]_9 ;
  output \rgf_c1bus_wb[1]_i_14 ;
  output \sr_reg[6]_10 ;
  output \badr[11]_INST_0_i_1 ;
  output \badr[6]_INST_0_i_1_0 ;
  output \badr[2]_INST_0_i_1_0 ;
  output \badr[10]_INST_0_i_1_0 ;
  output \stat_reg[2]_1 ;
  output \stat_reg[2]_2 ;
  output \rgf_c0bus_wb[15]_i_18_0 ;
  output \rgf_c0bus_wb[11]_i_3 ;
  output \tr_reg[7] ;
  output \rgf_c0bus_wb[11]_i_3_0 ;
  output \badr[6]_INST_0_i_2 ;
  output \tr_reg[6]_0 ;
  output \tr_reg[5]_0 ;
  output \sr_reg[6]_11 ;
  output \sr_reg[6]_12 ;
  output \badr[10]_INST_0_i_2 ;
  output \badr[14]_INST_0_i_2 ;
  output \rgf_c0bus_wb[13]_i_29_0 ;
  output \badr[4]_INST_0_i_2 ;
  output \badr[12]_INST_0_i_2 ;
  output \badr[8]_INST_0_i_2 ;
  output \rgf_c0bus_wb[7]_i_7 ;
  output \badr[6]_INST_0_i_2_0 ;
  output \badr[10]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[7]_i_7_0 ;
  output \sr_reg[6]_13 ;
  output \sr_reg[6]_14 ;
  output \badr[14]_INST_0_i_2_0 ;
  output \badr[1]_INST_0_i_2 ;
  output \sr_reg[6]_15 ;
  output \rgf_c0bus_wb[15]_i_26_0 ;
  output \sr_reg[6]_16 ;
  output \badr[3]_INST_0_i_2 ;
  output \badr[11]_INST_0_i_2 ;
  output \badr[7]_INST_0_i_2 ;
  output \rgf_c0bus_wb[11]_i_22 ;
  output \badr[6]_INST_0_i_2_1 ;
  output \badr[2]_INST_0_i_2 ;
  output \sr_reg[6]_17 ;
  output \sr_reg[6]_18 ;
  output \sr_reg[6]_19 ;
  output \rgf_c0bus_wb[10]_i_8_0 ;
  output \badr[5]_INST_0_i_2 ;
  output \badr[5]_INST_0_i_2_0 ;
  output \badr[1]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[11]_i_9 ;
  output \rgf_c0bus_wb[13]_i_28_0 ;
  output \badr[14]_INST_0_i_2_1 ;
  output \sr_reg[6]_20 ;
  output \sr_reg[6]_21 ;
  output \badr[12]_INST_0_i_2_0 ;
  output \rgf_c0bus_wb[11]_i_3_1 ;
  output \rgf_c1bus_wb[7]_i_4_0 ;
  output \sr_reg[6]_22 ;
  output \rgf_c0bus_wb[15]_i_6 ;
  output \rgf_c0bus_wb[15]_i_6_0 ;
  output \rgf_c0bus_wb[15]_i_6_1 ;
  output \rgf_c0bus_wb[11]_i_9_0 ;
  output \rgf_c0bus_wb[11]_i_9_1 ;
  output \rgf_c0bus_wb[11]_i_9_2 ;
  output \rgf_c0bus_wb[11]_i_3_2 ;
  output [15:0]Q;
  input \rgf_c1bus_wb[2]_i_7 ;
  input \rgf_c1bus_wb_reg[5] ;
  input \rgf_c1bus_wb[10]_i_14 ;
  input \rgf_c1bus_wb[14]_i_3 ;
  input \rgf_c1bus_wb[5]_i_10 ;
  input \rgf_c1bus_wb[14]_i_11 ;
  input \rgf_c1bus_wb[14]_i_11_0 ;
  input \rgf_c1bus_wb[14]_i_11_1 ;
  input \rgf_c1bus_wb[14]_i_11_2 ;
  input \rgf_c1bus_wb[14]_i_11_3 ;
  input \rgf_c1bus_wb[14]_i_11_4 ;
  input \rgf_c1bus_wb[11]_i_11 ;
  input \rgf_c1bus_wb[2]_i_7_0 ;
  input tout__1_carry__0_i_7__0;
  input tout__1_carry__0_i_7__0_0;
  input tout__1_carry__0_i_7__0_1;
  input tout__1_carry__0_i_7__0_2;
  input tout__1_carry__0_i_7__0_3;
  input tout__1_carry__0_i_7__0_4;
  input \rgf_c1bus_wb_reg[5]_0 ;
  input \rgf_c1bus_wb_reg[5]_1 ;
  input \rgf_c1bus_wb[4]_i_7_0 ;
  input \rgf_c1bus_wb[11]_i_11_0 ;
  input \rgf_c1bus_wb_reg[7] ;
  input \rgf_c1bus_wb[2]_i_7_1 ;
  input [0:0]\rgf_c0bus_wb[3]_i_7 ;
  input \rgf_c1bus_wb[3]_i_4 ;
  input \rgf_c1bus_wb[11]_i_11_1 ;
  input \rgf_c1bus_wb[2]_i_7_2 ;
  input \rgf_c1bus_wb[3]_i_4_0 ;
  input \rgf_c1bus_wb[8]_i_3 ;
  input \rgf_c1bus_wb_reg[3] ;
  input \rgf_c1bus_wb[8]_i_3_0 ;
  input \rgf_c1bus_wb[11]_i_11_2 ;
  input \rgf_c1bus_wb[11]_i_11_3 ;
  input \rgf_c1bus_wb[11]_i_11_4 ;
  input \rgf_c1bus_wb[11]_i_11_5 ;
  input \rgf_c1bus_wb_reg[4] ;
  input \rgf_c1bus_wb[4]_i_3_0 ;
  input \rgf_c1bus_wb[4]_i_3_1 ;
  input \rgf_c1bus_wb[4]_i_3_2 ;
  input \rgf_c1bus_wb[12]_i_2 ;
  input \rgf_c1bus_wb[12]_i_2_0 ;
  input \rgf_c1bus_wb[11]_i_8 ;
  input \rgf_c1bus_wb[11]_i_11_6 ;
  input \rgf_c1bus_wb[11]_i_8_0 ;
  input \rgf_c1bus_wb[10]_i_14_0 ;
  input \rgf_c1bus_wb[11]_i_8_1 ;
  input \rgf_c1bus_wb[1]_i_3 ;
  input \rgf_c1bus_wb_reg[1] ;
  input \rgf_c1bus_wb_reg[10] ;
  input \rgf_c1bus_wb_reg[1]_0 ;
  input \rgf_c1bus_wb[4]_i_7_1 ;
  input \rgf_c1bus_wb[4]_i_7_2 ;
  input \rgf_c1bus_wb[4]_i_7_3 ;
  input \rgf_c1bus_wb[4]_i_7_4 ;
  input \rgf_c1bus_wb[4]_i_7_5 ;
  input \rgf_c0bus_wb_reg[7]_i_11 ;
  input \rgf_c0bus_wb[1]_i_3 ;
  input \rgf_c0bus_wb[6]_i_11 ;
  input \rgf_c0bus_wb[7]_i_15_0 ;
  input \rgf_c0bus_wb[5]_i_8 ;
  input \rgf_c0bus_wb[11]_i_17 ;
  input \rgf_c0bus_wb[10]_i_26 ;
  input \bbus_o[7] ;
  input \bbus_o[7]_0 ;
  input \bbus_o[7]_1 ;
  input [2:0]p_1_in3_in;
  input [2:0]p_0_in2_in;
  input \bbus_o[7]_2 ;
  input \sr[4]_i_144 ;
  input \bbus_o[6] ;
  input \bbus_o[6]_0 ;
  input \bbus_o[6]_1 ;
  input \bbus_o[6]_2 ;
  input \bbus_o[5] ;
  input \bbus_o[5]_0 ;
  input \bbus_o[5]_1 ;
  input \bbus_o[5]_2 ;
  input \rgf_c0bus_wb_reg[10] ;
  input \rgf_c0bus_wb_reg[10]_0 ;
  input \rgf_c0bus_wb[13]_i_4 ;
  input \rgf_c0bus_wb[10]_i_4 ;
  input \rgf_c0bus_wb[5]_i_2 ;
  input \sr[4]_i_56 ;
  input \rgf_c0bus_wb_reg[10]_1 ;
  input \sr[4]_i_144_0 ;
  input \sr[4]_i_144_1 ;
  input \rgf_c0bus_wb[11]_i_17_0 ;
  input \rgf_c0bus_wb[11]_i_17_1 ;
  input \rgf_c0bus_wb[10]_i_26_0 ;
  input \rgf_c0bus_wb[11]_i_17_2 ;
  input \rgf_c0bus_wb[11]_i_17_3 ;
  input \rgf_c0bus_wb[7]_i_15_1 ;
  input \rgf_c0bus_wb[11]_i_17_4 ;
  input \rgf_c0bus_wb[5]_i_8_0 ;
  input \rgf_c0bus_wb[5]_i_8_1 ;
  input \rgf_c0bus_wb[0]_i_8 ;
  input \rgf_c0bus_wb[5]_i_8_2 ;
  input \rgf_c0bus_wb[10]_i_26_1 ;
  input \rgf_c0bus_wb[4]_i_3 ;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1 ;
  wire \badr[10]_INST_0_i_1_0 ;
  wire \badr[10]_INST_0_i_2 ;
  wire \badr[10]_INST_0_i_2_0 ;
  wire \badr[11]_INST_0_i_1 ;
  wire \badr[11]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_1 ;
  wire \badr[12]_INST_0_i_2 ;
  wire \badr[12]_INST_0_i_2_0 ;
  wire \badr[13]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire \badr[14]_INST_0_i_2 ;
  wire \badr[14]_INST_0_i_2_0 ;
  wire \badr[14]_INST_0_i_2_1 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_1_0 ;
  wire \badr[1]_INST_0_i_2 ;
  wire \badr[1]_INST_0_i_2_0 ;
  wire \badr[2]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1_0 ;
  wire \badr[2]_INST_0_i_2 ;
  wire \badr[3]_INST_0_i_1 ;
  wire \badr[3]_INST_0_i_2 ;
  wire \badr[4]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_2 ;
  wire \badr[5]_INST_0_i_2_0 ;
  wire \badr[6]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1_0 ;
  wire \badr[6]_INST_0_i_2 ;
  wire \badr[6]_INST_0_i_2_0 ;
  wire \badr[6]_INST_0_i_2_1 ;
  wire \badr[7]_INST_0_i_2 ;
  wire \badr[8]_INST_0_i_2 ;
  wire \badr[9]_INST_0_i_1 ;
  wire \badr[9]_INST_0_i_1_0 ;
  wire \bbus_o[5] ;
  wire \bbus_o[5]_0 ;
  wire \bbus_o[5]_1 ;
  wire \bbus_o[5]_2 ;
  wire \bbus_o[6] ;
  wire \bbus_o[6]_0 ;
  wire \bbus_o[6]_1 ;
  wire \bbus_o[6]_2 ;
  wire \bbus_o[7] ;
  wire \bbus_o[7]_0 ;
  wire \bbus_o[7]_1 ;
  wire \bbus_o[7]_2 ;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire [2:0]p_0_in2_in;
  wire [2:0]p_1_in3_in;
  wire \rgf_c0bus_wb[0]_i_8 ;
  wire \rgf_c0bus_wb[10]_i_26 ;
  wire \rgf_c0bus_wb[10]_i_26_0 ;
  wire \rgf_c0bus_wb[10]_i_26_1 ;
  wire \rgf_c0bus_wb[10]_i_4 ;
  wire \rgf_c0bus_wb[10]_i_8_0 ;
  wire \rgf_c0bus_wb[11]_i_17 ;
  wire \rgf_c0bus_wb[11]_i_17_0 ;
  wire \rgf_c0bus_wb[11]_i_17_1 ;
  wire \rgf_c0bus_wb[11]_i_17_2 ;
  wire \rgf_c0bus_wb[11]_i_17_3 ;
  wire \rgf_c0bus_wb[11]_i_17_4 ;
  wire \rgf_c0bus_wb[11]_i_22 ;
  wire \rgf_c0bus_wb[11]_i_3 ;
  wire \rgf_c0bus_wb[11]_i_3_0 ;
  wire \rgf_c0bus_wb[11]_i_3_1 ;
  wire \rgf_c0bus_wb[11]_i_3_2 ;
  wire \rgf_c0bus_wb[11]_i_9 ;
  wire \rgf_c0bus_wb[11]_i_9_0 ;
  wire \rgf_c0bus_wb[11]_i_9_1 ;
  wire \rgf_c0bus_wb[11]_i_9_2 ;
  wire \rgf_c0bus_wb[13]_i_28_0 ;
  wire \rgf_c0bus_wb[13]_i_29_0 ;
  wire \rgf_c0bus_wb[13]_i_4 ;
  wire \rgf_c0bus_wb[15]_i_18_0 ;
  wire \rgf_c0bus_wb[15]_i_26_0 ;
  wire \rgf_c0bus_wb[15]_i_6 ;
  wire \rgf_c0bus_wb[15]_i_6_0 ;
  wire \rgf_c0bus_wb[15]_i_6_1 ;
  wire \rgf_c0bus_wb[1]_i_3 ;
  wire [0:0]\rgf_c0bus_wb[3]_i_7 ;
  wire \rgf_c0bus_wb[4]_i_3 ;
  wire \rgf_c0bus_wb[5]_i_2 ;
  wire \rgf_c0bus_wb[5]_i_8 ;
  wire \rgf_c0bus_wb[5]_i_8_0 ;
  wire \rgf_c0bus_wb[5]_i_8_1 ;
  wire \rgf_c0bus_wb[5]_i_8_2 ;
  wire \rgf_c0bus_wb[6]_i_11 ;
  wire \rgf_c0bus_wb[7]_i_15_0 ;
  wire \rgf_c0bus_wb[7]_i_15_1 ;
  wire \rgf_c0bus_wb[7]_i_16_n_0 ;
  wire \rgf_c0bus_wb[7]_i_17_n_0 ;
  wire \rgf_c0bus_wb[7]_i_18_n_0 ;
  wire \rgf_c0bus_wb[7]_i_7 ;
  wire \rgf_c0bus_wb[7]_i_7_0 ;
  wire \rgf_c0bus_wb_reg[10] ;
  wire \rgf_c0bus_wb_reg[10]_0 ;
  wire \rgf_c0bus_wb_reg[10]_1 ;
  wire \rgf_c0bus_wb_reg[7]_i_11 ;
  wire \rgf_c1bus_wb[10]_i_14 ;
  wire \rgf_c1bus_wb[10]_i_14_0 ;
  wire \rgf_c1bus_wb[10]_i_6_n_0 ;
  wire \rgf_c1bus_wb[11]_i_10 ;
  wire \rgf_c1bus_wb[11]_i_11 ;
  wire \rgf_c1bus_wb[11]_i_11_0 ;
  wire \rgf_c1bus_wb[11]_i_11_1 ;
  wire \rgf_c1bus_wb[11]_i_11_2 ;
  wire \rgf_c1bus_wb[11]_i_11_3 ;
  wire \rgf_c1bus_wb[11]_i_11_4 ;
  wire \rgf_c1bus_wb[11]_i_11_5 ;
  wire \rgf_c1bus_wb[11]_i_11_6 ;
  wire \rgf_c1bus_wb[11]_i_13_0 ;
  wire \rgf_c1bus_wb[11]_i_8 ;
  wire \rgf_c1bus_wb[11]_i_8_0 ;
  wire \rgf_c1bus_wb[11]_i_8_1 ;
  wire \rgf_c1bus_wb[12]_i_2 ;
  wire \rgf_c1bus_wb[12]_i_20 ;
  wire \rgf_c1bus_wb[12]_i_2_0 ;
  wire \rgf_c1bus_wb[13]_i_16_0 ;
  wire \rgf_c1bus_wb[13]_i_9_0 ;
  wire \rgf_c1bus_wb[14]_i_11 ;
  wire \rgf_c1bus_wb[14]_i_11_0 ;
  wire \rgf_c1bus_wb[14]_i_11_1 ;
  wire \rgf_c1bus_wb[14]_i_11_2 ;
  wire \rgf_c1bus_wb[14]_i_11_3 ;
  wire \rgf_c1bus_wb[14]_i_11_4 ;
  wire \rgf_c1bus_wb[14]_i_28 ;
  wire \rgf_c1bus_wb[14]_i_28_0 ;
  wire \rgf_c1bus_wb[14]_i_28_1 ;
  wire \rgf_c1bus_wb[14]_i_28_2 ;
  wire \rgf_c1bus_wb[14]_i_28_3 ;
  wire \rgf_c1bus_wb[14]_i_3 ;
  wire \rgf_c1bus_wb[14]_i_30_0 ;
  wire \rgf_c1bus_wb[14]_i_32_0 ;
  wire \rgf_c1bus_wb[14]_i_32_1 ;
  wire \rgf_c1bus_wb[15]_i_14 ;
  wire \rgf_c1bus_wb[1]_i_14 ;
  wire \rgf_c1bus_wb[1]_i_3 ;
  wire \rgf_c1bus_wb[2]_i_7 ;
  wire \rgf_c1bus_wb[2]_i_7_0 ;
  wire \rgf_c1bus_wb[2]_i_7_1 ;
  wire \rgf_c1bus_wb[2]_i_7_2 ;
  wire \rgf_c1bus_wb[3]_i_4 ;
  wire \rgf_c1bus_wb[3]_i_4_0 ;
  wire \rgf_c1bus_wb[4]_i_20_n_0 ;
  wire \rgf_c1bus_wb[4]_i_3_0 ;
  wire \rgf_c1bus_wb[4]_i_3_1 ;
  wire \rgf_c1bus_wb[4]_i_3_2 ;
  wire \rgf_c1bus_wb[4]_i_7_0 ;
  wire \rgf_c1bus_wb[4]_i_7_1 ;
  wire \rgf_c1bus_wb[4]_i_7_2 ;
  wire \rgf_c1bus_wb[4]_i_7_3 ;
  wire \rgf_c1bus_wb[4]_i_7_4 ;
  wire \rgf_c1bus_wb[4]_i_7_5 ;
  wire \rgf_c1bus_wb[4]_i_7_n_0 ;
  wire \rgf_c1bus_wb[4]_i_9_0 ;
  wire \rgf_c1bus_wb[5]_i_10 ;
  wire \rgf_c1bus_wb[7]_i_4 ;
  wire \rgf_c1bus_wb[7]_i_4_0 ;
  wire \rgf_c1bus_wb[8]_i_3 ;
  wire \rgf_c1bus_wb[8]_i_3_0 ;
  wire \rgf_c1bus_wb[9]_i_17 ;
  wire \rgf_c1bus_wb_reg[10] ;
  wire \rgf_c1bus_wb_reg[1] ;
  wire \rgf_c1bus_wb_reg[1]_0 ;
  wire \rgf_c1bus_wb_reg[3] ;
  wire \rgf_c1bus_wb_reg[4] ;
  wire \rgf_c1bus_wb_reg[5] ;
  wire \rgf_c1bus_wb_reg[5]_0 ;
  wire \rgf_c1bus_wb_reg[5]_1 ;
  wire \rgf_c1bus_wb_reg[7] ;
  wire \sr[4]_i_144 ;
  wire \sr[4]_i_144_0 ;
  wire \sr[4]_i_144_1 ;
  wire \sr[4]_i_56 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_11 ;
  wire \sr_reg[6]_12 ;
  wire \sr_reg[6]_13 ;
  wire \sr_reg[6]_14 ;
  wire \sr_reg[6]_15 ;
  wire \sr_reg[6]_16 ;
  wire \sr_reg[6]_17 ;
  wire \sr_reg[6]_18 ;
  wire \sr_reg[6]_19 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_20 ;
  wire \sr_reg[6]_21 ;
  wire \sr_reg[6]_22 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_7 ;
  wire \sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;
  wire \stat_reg[2] ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire tout__1_carry__0_i_7__0;
  wire tout__1_carry__0_i_7__0_0;
  wire tout__1_carry__0_i_7__0_1;
  wire tout__1_carry__0_i_7__0_2;
  wire tout__1_carry__0_i_7__0_3;
  wire tout__1_carry__0_i_7__0_4;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[7] ;

  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bbus_o[5]_INST_0_i_1 
       (.I0(\bbus_o[5] ),
        .I1(\bbus_o[5]_0 ),
        .I2(\bbus_o[5]_1 ),
        .I3(p_1_in3_in[0]),
        .I4(p_0_in2_in[0]),
        .I5(\bbus_o[5]_2 ),
        .O(\tr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bbus_o[6]_INST_0_i_1 
       (.I0(\bbus_o[6] ),
        .I1(\bbus_o[6]_0 ),
        .I2(\bbus_o[6]_1 ),
        .I3(p_1_in3_in[1]),
        .I4(p_0_in2_in[1]),
        .I5(\bbus_o[6]_2 ),
        .O(\tr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[7]_INST_0_i_1 
       (.I0(\bbus_o[7] ),
        .I1(\bbus_o[7]_0 ),
        .I2(\bbus_o[7]_1 ),
        .I3(p_1_in3_in[2]),
        .I4(p_0_in2_in[2]),
        .I5(\bbus_o[7]_2 ),
        .O(\tr_reg[7] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[13]_INST_0_i_16 
       (.I0(tout__1_carry__0_i_7__0),
        .I1(tout__1_carry__0_i_7__0_0),
        .I2(tout__1_carry__0_i_7__0_1),
        .I3(tout__1_carry__0_i_7__0_2),
        .I4(tout__1_carry__0_i_7__0_3),
        .I5(tout__1_carry__0_i_7__0_4),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_16 
       (.I0(\rgf_c1bus_wb[14]_i_11 ),
        .I1(\rgf_c1bus_wb[14]_i_11_0 ),
        .I2(\rgf_c1bus_wb[14]_i_11_1 ),
        .I3(\rgf_c1bus_wb[14]_i_11_2 ),
        .I4(\rgf_c1bus_wb[14]_i_11_3 ),
        .I5(\rgf_c1bus_wb[14]_i_11_4 ),
        .O(\tr_reg[6] ));
  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT4 #(
    .INIT(16'hFFE2)) 
    \rgf_c0bus_wb[10]_i_14 
       (.I0(\badr[14]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_0 ),
        .I2(\sr_reg[6]_14 ),
        .I3(\rgf_c0bus_wb[10]_i_4 ),
        .O(\sr_reg[6]_15 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[10]_i_19 
       (.I0(\rgf_c0bus_wb[7]_i_15_0 ),
        .I1(\sr[4]_i_144_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[5]_i_8_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\sr[4]_i_144 ),
        .O(\badr[6]_INST_0_i_2_1 ));
  LUT6 #(
    .INIT(64'hAACCFFFFF0FFFFFF)) 
    \rgf_c0bus_wb[10]_i_2 
       (.I0(\sr_reg[6]_14 ),
        .I1(\badr[14]_INST_0_i_2_0 ),
        .I2(\badr[1]_INST_0_i_2 ),
        .I3(\rgf_c0bus_wb_reg[10]_0 ),
        .I4(\rgf_c0bus_wb_reg[10] ),
        .I5(\rgf_c0bus_wb_reg[10]_1 ),
        .O(\sr_reg[6]_13 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[10]_i_20 
       (.I0(\rgf_c0bus_wb[5]_i_8 ),
        .I1(\rgf_c0bus_wb[5]_i_8_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[5]_i_8_2 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[10]_i_26_1 ),
        .O(\badr[2]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[10]_i_21 
       (.I0(\rgf_c0bus_wb[11]_i_17_3 ),
        .I1(\rgf_c0bus_wb[11]_i_17_2 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[10]_i_26_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[11]_i_17 ),
        .O(\badr[11]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[10]_i_22 
       (.I0(\rgf_c0bus_wb[3]_i_7 ),
        .I1(\rgf_c0bus_wb[0]_i_8 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[11]_i_17_4 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[7]_i_15_1 ),
        .O(\sr_reg[6]_17 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[10]_i_24 
       (.I0(\rgf_c0bus_wb[7]_i_15_1 ),
        .I1(\rgf_c0bus_wb[11]_i_17_0 ),
        .O(\rgf_c0bus_wb[11]_i_22 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[10]_i_27 
       (.I0(\rgf_c0bus_wb[10]_i_26_1 ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .O(\rgf_c0bus_wb[11]_i_3_2 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_c0bus_wb[10]_i_28 
       (.I0(\rgf_c0bus_wb[10]_i_26_0 ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .O(\rgf_c0bus_wb[11]_i_3_1 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[10]_i_6 
       (.I0(\rgf_c0bus_wb[0]_i_8 ),
        .I1(\rgf_c0bus_wb[3]_i_7 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[10]_i_26_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[5]_i_8_2 ),
        .O(\sr_reg[6]_14 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[10]_i_7 
       (.I0(\rgf_c0bus_wb[11]_i_17_2 ),
        .I1(\rgf_c0bus_wb[11]_i_17_3 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[7]_i_15_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[11]_i_17_4 ),
        .O(\badr[14]_INST_0_i_2_0 ));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    \rgf_c0bus_wb[10]_i_8 
       (.I0(\rgf_c0bus_wb[0]_i_8 ),
        .I1(\rgf_c0bus_wb[11]_i_17_0 ),
        .I2(\rgf_c0bus_wb[10]_i_26_1 ),
        .I3(\rgf_c0bus_wb[11]_i_17_1 ),
        .I4(\rgf_c0bus_wb[5]_i_8_2 ),
        .O(\badr[1]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[10]_i_9 
       (.I0(\rgf_c0bus_wb[5]_i_8_1 ),
        .I1(\rgf_c0bus_wb[5]_i_8 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\sr[4]_i_144 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[5]_i_8_0 ),
        .O(\badr[5]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c0bus_wb[11]_i_13 
       (.I0(\rgf_c0bus_wb[3]_i_7 ),
        .I1(\rgf_c0bus_wb[7]_i_15_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_4 ),
        .I3(\rgf_c0bus_wb[11]_i_17_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_2 ),
        .I5(\rgf_c0bus_wb[11]_i_17_0 ),
        .O(\sr_reg[6]_21 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[11]_i_23 
       (.I0(\rgf_c0bus_wb[5]_i_8_1 ),
        .I1(\rgf_c0bus_wb[5]_i_8_0 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[10]_i_26_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[5]_i_8 ),
        .O(\badr[3]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[11]_i_24 
       (.I0(\sr[4]_i_144_1 ),
        .I1(\sr[4]_i_144_0 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\sr[4]_i_144 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[7]_i_15_0 ),
        .O(\badr[7]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[11]_i_25 
       (.I0(\rgf_c0bus_wb[0]_i_8 ),
        .I1(\rgf_c0bus_wb[5]_i_8_2 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[7]_i_15_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[3]_i_7 ),
        .O(\sr_reg[6]_16 ));
  LUT5 #(
    .INIT(32'hA0AF3F30)) 
    \rgf_c0bus_wb[11]_i_26 
       (.I0(\tr_reg[7] ),
        .I1(\rgf_c0bus_wb[5]_i_8 ),
        .I2(\rgf_c0bus_wb[1]_i_3 ),
        .I3(\rgf_c0bus_wb[11]_i_17 ),
        .I4(\rgf_c0bus_wb[10]_i_26 ),
        .O(\rgf_c0bus_wb[11]_i_3_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[11]_i_8 
       (.I0(\rgf_c0bus_wb[11]_i_17_2 ),
        .I1(\rgf_c0bus_wb[11]_i_17_4 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[11]_i_17 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[11]_i_17_3 ),
        .O(\badr[12]_INST_0_i_2_0 ));
  LUT4 #(
    .INIT(16'h2EFF)) 
    \rgf_c0bus_wb[12]_i_14 
       (.I0(\rgf_c0bus_wb[5]_i_8_1 ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .I2(\tr_reg[7] ),
        .I3(\rgf_c0bus_wb[1]_i_3 ),
        .O(\rgf_c0bus_wb[15]_i_6 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[13]_i_14 
       (.I0(\badr[4]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb[13]_i_4 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\badr[12]_INST_0_i_2 ),
        .I4(\rgf_c0bus_wb_reg[10]_0 ),
        .I5(\badr[8]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[13]_i_29_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[13]_i_19 
       (.I0(\rgf_c0bus_wb[10]_i_26_1 ),
        .I1(\rgf_c0bus_wb[5]_i_8 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[5]_i_8_2 ),
        .O(\badr[1]_INST_0_i_2_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[13]_i_20 
       (.I0(\rgf_c0bus_wb[7]_i_15_1 ),
        .I1(\rgf_c0bus_wb[3]_i_7 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[11]_i_17_2 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[11]_i_17_4 ),
        .O(\sr_reg[6]_12 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[13]_i_22 
       (.I0(\sr[4]_i_144 ),
        .I1(\rgf_c0bus_wb[7]_i_15_0 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[5]_i_8_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[5]_i_8_0 ),
        .O(\badr[5]_INST_0_i_2_0 ));
  LUT6 #(
    .INIT(64'hB8BBB888AAAAAAAA)) 
    \rgf_c0bus_wb[13]_i_24 
       (.I0(\rgf_c0bus_wb[7]_i_15_1 ),
        .I1(\rgf_c0bus_wb[11]_i_17_0 ),
        .I2(\rgf_c0bus_wb[11]_i_17_2 ),
        .I3(\rgf_c0bus_wb[11]_i_17_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_4 ),
        .I5(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_9 ));
  LUT6 #(
    .INIT(64'h331DFF1DFFFFFFFF)) 
    \rgf_c0bus_wb[13]_i_26 
       (.I0(\rgf_c0bus_wb[11]_i_17_4 ),
        .I1(\rgf_c0bus_wb[11]_i_17_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_2 ),
        .I3(\rgf_c0bus_wb[11]_i_17_0 ),
        .I4(\rgf_c0bus_wb[7]_i_15_1 ),
        .I5(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_9_1 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[13]_i_28 
       (.I0(\rgf_c0bus_wb[5]_i_8 ),
        .I1(\rgf_c0bus_wb[10]_i_26_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[5]_i_8_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[5]_i_8_1 ),
        .O(\badr[4]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[13]_i_29 
       (.I0(\rgf_c0bus_wb[7]_i_15_0 ),
        .I1(\sr[4]_i_144 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\sr[4]_i_144_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\sr[4]_i_144_1 ),
        .O(\badr[8]_INST_0_i_2 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[15]_i_18 
       (.I0(\tr_reg[7] ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .O(\rgf_c0bus_wb[11]_i_3 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[15]_i_26 
       (.I0(\sr[4]_i_144_0 ),
        .I1(\sr[4]_i_144_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[11]_i_17 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[10]_i_26_0 ),
        .O(\badr[10]_INST_0_i_2_0 ));
  LUT6 #(
    .INIT(64'h00F0101000F0D0D0)) 
    \rgf_c0bus_wb[1]_i_6 
       (.I0(\sr_reg[6]_12 ),
        .I1(\rgf_c0bus_wb[1]_i_3 ),
        .I2(\rgf_c0bus_wb_reg[10] ),
        .I3(\badr[10]_INST_0_i_2 ),
        .I4(\rgf_c0bus_wb_reg[10]_0 ),
        .I5(\badr[14]_INST_0_i_2 ),
        .O(\sr_reg[6]_11 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c0bus_wb[2]_i_5 
       (.I0(\badr[6]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_0 ),
        .I2(\badr[10]_INST_0_i_2_0 ),
        .I3(\rgf_c0bus_wb[10]_i_4 ),
        .O(\rgf_c0bus_wb[7]_i_7 ));
  LUT6 #(
    .INIT(64'h331DFF1DFFFFFFFF)) 
    \rgf_c0bus_wb[2]_i_7 
       (.I0(\rgf_c0bus_wb[5]_i_8_2 ),
        .I1(\rgf_c0bus_wb[11]_i_17_1 ),
        .I2(\rgf_c0bus_wb[10]_i_26_1 ),
        .I3(\rgf_c0bus_wb[11]_i_17_0 ),
        .I4(\rgf_c0bus_wb[0]_i_8 ),
        .I5(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_9_0 ));
  LUT6 #(
    .INIT(64'hFF1D001DFFFFFFFF)) 
    \rgf_c0bus_wb[4]_i_12 
       (.I0(\rgf_c0bus_wb[11]_i_17_2 ),
        .I1(\rgf_c0bus_wb[11]_i_17_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_3 ),
        .I3(\rgf_c0bus_wb[11]_i_17_0 ),
        .I4(\rgf_c0bus_wb[4]_i_3 ),
        .I5(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\rgf_c0bus_wb[11]_i_9_2 ));
  LUT4 #(
    .INIT(16'h001D)) 
    \rgf_c0bus_wb[5]_i_7 
       (.I0(\rgf_c0bus_wb[5]_i_2 ),
        .I1(\rgf_c0bus_wb_reg[10]_0 ),
        .I2(\sr[4]_i_56 ),
        .I3(\rgf_c0bus_wb[10]_i_4 ),
        .O(\rgf_c0bus_wb[7]_i_7_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c0bus_wb[6]_i_14 
       (.I0(\tr_reg[6]_0 ),
        .I1(\rgf_c0bus_wb[6]_i_11 ),
        .I2(\sr[4]_i_144 ),
        .O(\badr[6]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[6]_i_5 
       (.I0(\badr[5]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb_reg[10]_0 ),
        .I2(\badr[1]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[10]_i_8_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[6]_i_6 
       (.I0(\badr[14]_INST_0_i_2_0 ),
        .I1(\rgf_c0bus_wb_reg[10]_0 ),
        .I2(\badr[10]_INST_0_i_2_0 ),
        .O(\rgf_c0bus_wb[15]_i_26_0 ));
  LUT6 #(
    .INIT(64'h0074007400743374)) 
    \rgf_c0bus_wb[7]_i_15 
       (.I0(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_11 ),
        .I2(\rgf_c0bus_wb[7]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_3 ),
        .I4(\rgf_c0bus_wb[7]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_3 ),
        .O(\rgf_c0bus_wb[15]_i_18_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c0bus_wb[7]_i_16 
       (.I0(\tr_reg[7] ),
        .I1(\rgf_c0bus_wb[6]_i_11 ),
        .I2(\rgf_c0bus_wb[7]_i_15_0 ),
        .O(\rgf_c0bus_wb[7]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_c0bus_wb[7]_i_17 
       (.I0(\rgf_c0bus_wb[7]_i_15_0 ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .O(\rgf_c0bus_wb[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[7]_i_18 
       (.I0(\rgf_c0bus_wb[7]_i_15_1 ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .O(\rgf_c0bus_wb[7]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[7]_i_6 
       (.I0(\rgf_c0bus_wb[5]_i_8_0 ),
        .I1(\rgf_c0bus_wb[5]_i_8_1 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[7]_i_15_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\sr[4]_i_144 ),
        .O(\badr[6]_INST_0_i_2_0 ));
  LUT4 #(
    .INIT(16'h74FF)) 
    \rgf_c0bus_wb[8]_i_17 
       (.I0(\tr_reg[7] ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .I2(\rgf_c0bus_wb[0]_i_8 ),
        .I3(\rgf_c0bus_wb[1]_i_3 ),
        .O(\rgf_c0bus_wb[15]_i_6_1 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[8]_i_8 
       (.I0(\rgf_c0bus_wb[11]_i_17 ),
        .I1(\rgf_c0bus_wb[10]_i_26_0 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[11]_i_17_2 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[11]_i_17_3 ),
        .O(\badr[12]_INST_0_i_2 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[8]_i_9 
       (.I0(\rgf_c0bus_wb[7]_i_15_1 ),
        .I1(\rgf_c0bus_wb[11]_i_17_4 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[0]_i_8 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[3]_i_7 ),
        .O(\sr_reg[6]_20 ));
  LUT4 #(
    .INIT(16'h2EFF)) 
    \rgf_c0bus_wb[9]_i_17 
       (.I0(\rgf_c0bus_wb[5]_i_8_2 ),
        .I1(\rgf_c0bus_wb[10]_i_26 ),
        .I2(\tr_reg[7] ),
        .I3(\rgf_c0bus_wb[1]_i_3 ),
        .O(\rgf_c0bus_wb[15]_i_6_0 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c0bus_wb[9]_i_19 
       (.I0(\rgf_c0bus_wb[5]_i_8_2 ),
        .I1(\rgf_c0bus_wb[0]_i_8 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\rgf_c0bus_wb[3]_i_7 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[7]_i_15_1 ),
        .O(\sr_reg[6]_19 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c0bus_wb[9]_i_21 
       (.I0(\rgf_c0bus_wb[11]_i_17 ),
        .I1(\rgf_c0bus_wb[11]_i_17_3 ),
        .I2(\rgf_c0bus_wb[11]_i_17_0 ),
        .I3(\sr[4]_i_144_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_1 ),
        .I5(\rgf_c0bus_wb[10]_i_26_0 ),
        .O(\badr[10]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h47444777)) 
    \rgf_c0bus_wb[9]_i_22 
       (.I0(\rgf_c0bus_wb[7]_i_15_1 ),
        .I1(\rgf_c0bus_wb[11]_i_17_0 ),
        .I2(\rgf_c0bus_wb[11]_i_17_2 ),
        .I3(\rgf_c0bus_wb[11]_i_17_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_4 ),
        .O(\badr[14]_INST_0_i_2 ));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    \rgf_c0bus_wb[9]_i_23 
       (.I0(\rgf_c0bus_wb[7]_i_15_1 ),
        .I1(\rgf_c0bus_wb[11]_i_17_0 ),
        .I2(\rgf_c0bus_wb[11]_i_17_2 ),
        .I3(\rgf_c0bus_wb[11]_i_17_1 ),
        .I4(\rgf_c0bus_wb[11]_i_17_4 ),
        .O(\badr[14]_INST_0_i_2_1 ));
  LUT3 #(
    .INIT(8'h5C)) 
    \rgf_c0bus_wb[9]_i_6 
       (.I0(\sr_reg[6]_19 ),
        .I1(\sr[4]_i_56 ),
        .I2(\rgf_c0bus_wb_reg[10]_0 ),
        .O(\sr_reg[6]_18 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_7 
       (.I0(\badr[8]_INST_0_i_2 ),
        .I1(\rgf_c0bus_wb_reg[10]_0 ),
        .I2(\badr[4]_INST_0_i_2 ),
        .O(\rgf_c0bus_wb[13]_i_28_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c1bus_wb[0]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_28_2 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb[14]_i_28_0 ),
        .I3(\rgf_c1bus_wb_reg[3] ),
        .O(\rgf_c1bus_wb[7]_i_4_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[10]_i_11 
       (.I0(\rgf_c1bus_wb[2]_i_7_2 ),
        .I1(\rgf_c1bus_wb[2]_i_7_0 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[11]_i_11_2 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_1 ),
        .O(\badr[11]_INST_0_i_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[10]_i_15 
       (.I0(\rgf_c1bus_wb[10]_i_14_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14 ),
        .O(\stat_reg[2]_2 ));
  LUT6 #(
    .INIT(64'h000CCC0C88888888)) 
    \rgf_c1bus_wb[10]_i_2 
       (.I0(\rgf_c1bus_wb[10]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb_reg[10] ),
        .I2(\rgf_c1bus_wb[14]_i_28_3 ),
        .I3(\rgf_c1bus_wb_reg[7] ),
        .I4(\badr[9]_INST_0_i_1_0 ),
        .I5(\rgf_c1bus_wb_reg[5]_1 ),
        .O(\rgf_c1bus_wb[15]_i_14 ));
  LUT5 #(
    .INIT(32'hAFA0CFCF)) 
    \rgf_c1bus_wb[10]_i_6 
       (.I0(\sr_reg[6]_8 ),
        .I1(\badr[14]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb_reg[4] ),
        .I3(\badr[2]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \rgf_c1bus_wb[10]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_11_6 ),
        .I1(\rgf_c1bus_wb[11]_i_8_1 ),
        .I2(\rgf_c1bus_wb[14]_i_3 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_3 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[10]_i_8 
       (.I0(\rgf_c1bus_wb[11]_i_11_4 ),
        .I1(\rgf_c1bus_wb[11]_i_11_5 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[11]_i_11_2 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_3 ),
        .O(\badr[9]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c1bus_wb[11]_i_13 
       (.I0(\rgf_c1bus_wb[11]_i_11_1 ),
        .I1(\rgf_c1bus_wb[2]_i_7_2 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[2]_i_7_0 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[2]_i_7 ),
        .O(\badr[14]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[11]_i_14 
       (.I0(\rgf_c1bus_wb[11]_i_8_0 ),
        .I1(\rgf_c1bus_wb[11]_i_8 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[11]_i_8_1 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[10]_i_14_0 ),
        .O(\badr[2]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000CCAACCAA)) 
    \rgf_c1bus_wb[11]_i_9 
       (.I0(\rgf_c1bus_wb[2]_i_7_1 ),
        .I1(\rgf_c0bus_wb[3]_i_7 ),
        .I2(\rgf_c1bus_wb[2]_i_7 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[2]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\sr_reg[6]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[12]_i_11 
       (.I0(\rgf_c1bus_wb[3]_i_4_0 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb[3]_i_4 ),
        .O(\rgf_c1bus_wb[12]_i_20 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[12]_i_18 
       (.I0(\rgf_c1bus_wb[2]_i_7_1 ),
        .I1(\rgf_c1bus_wb[2]_i_7 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c0bus_wb[3]_i_7 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_8 ),
        .O(\sr_reg[6]_9 ));
  LUT4 #(
    .INIT(16'h7477)) 
    \rgf_c1bus_wb[12]_i_7 
       (.I0(\rgf_c1bus_wb[12]_i_2 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb[12]_i_2_0 ),
        .I3(\rgf_c1bus_wb[11]_i_8 ),
        .O(\badr[0]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[13]_i_10 
       (.I0(\sr_reg[6]_3 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\badr[3]_INST_0_i_1 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \rgf_c1bus_wb[13]_i_16 
       (.I0(\rgf_c1bus_wb[11]_i_8_1 ),
        .I1(\rgf_c1bus_wb[10]_i_14_0 ),
        .I2(\rgf_c1bus_wb[11]_i_11 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11_6 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_2 ));
  LUT6 #(
    .INIT(64'hFFF000F0AACCAACC)) 
    \rgf_c1bus_wb[13]_i_18 
       (.I0(\rgf_c1bus_wb[11]_i_8_0 ),
        .I1(\rgf_c1bus_wb[11]_i_8 ),
        .I2(\rgf_c1bus_wb[2]_i_7_1 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c0bus_wb[3]_i_7 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\sr_reg[6]_5 ));
  LUT6 #(
    .INIT(64'h303F5050303F5F5F)) 
    \rgf_c1bus_wb[13]_i_19 
       (.I0(\rgf_c0bus_wb[3]_i_7 ),
        .I1(\rgf_c1bus_wb[2]_i_7_1 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[2]_i_7_0 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[2]_i_7 ),
        .O(\sr_reg[6]_3 ));
  LUT6 #(
    .INIT(64'h05F5030305F5F3F3)) 
    \rgf_c1bus_wb[13]_i_20 
       (.I0(\rgf_c1bus_wb[11]_i_8 ),
        .I1(\rgf_c1bus_wb[11]_i_8_0 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[10]_i_14_0 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_8_1 ),
        .O(\badr[3]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c1bus_wb[13]_i_21 
       (.I0(\rgf_c1bus_wb[11]_i_11_6 ),
        .I1(\rgf_c1bus_wb[11]_i_11 ),
        .I2(\rgf_c1bus_wb[14]_i_3 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11_5 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_1 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c1bus_wb[13]_i_22 
       (.I0(\rgf_c1bus_wb[11]_i_11_4 ),
        .I1(\rgf_c1bus_wb[11]_i_11_3 ),
        .I2(\rgf_c1bus_wb[11]_i_11_2 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11_1 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\rgf_c1bus_wb[14]_i_28 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[13]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_28_2 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\sr_reg[6]_5 ),
        .O(\sr_reg[6]_4 ));
  LUT6 #(
    .INIT(64'hFFB8FFFF00B80000)) 
    \rgf_c1bus_wb[13]_i_9 
       (.I0(\rgf_c1bus_wb[2]_i_7_0 ),
        .I1(\rgf_c1bus_wb[4]_i_7_0 ),
        .I2(\rgf_c1bus_wb[2]_i_7 ),
        .I3(\rgf_c1bus_wb[11]_i_11_0 ),
        .I4(\rgf_c1bus_wb_reg[7] ),
        .I5(\rgf_c1bus_wb[2]_i_7_1 ),
        .O(\badr[15]_INST_0_i_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[14]_i_10 
       (.I0(\rgf_c1bus_wb[14]_i_3 ),
        .I1(\rgf_c1bus_wb[10]_i_14 ),
        .O(\stat_reg[2]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_17 
       (.I0(\sr_reg[6]_7 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb_reg[1] ),
        .O(\sr_reg[6]_6 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_18 
       (.I0(\rgf_c1bus_wb_reg[1]_0 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\badr[10]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[14]_i_30_0 ));
  LUT6 #(
    .INIT(64'h505F3F3F505F3030)) 
    \rgf_c1bus_wb[14]_i_20 
       (.I0(\badr[13]_INST_0_i_1 ),
        .I1(\badr[9]_INST_0_i_1_0 ),
        .I2(\rgf_c1bus_wb_reg[5]_1 ),
        .I3(\rgf_c1bus_wb[14]_i_28_3 ),
        .I4(\rgf_c1bus_wb_reg[7] ),
        .I5(\badr[2]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[14]_i_32_0 ));
  LUT6 #(
    .INIT(64'h000FFF0F55335533)) 
    \rgf_c1bus_wb[14]_i_29 
       (.I0(\rgf_c1bus_wb[2]_i_7 ),
        .I1(\rgf_c1bus_wb[2]_i_7_1 ),
        .I2(\rgf_c1bus_wb[11]_i_8 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c0bus_wb[3]_i_7 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\sr_reg[6]_7 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[14]_i_30 
       (.I0(\rgf_c1bus_wb[11]_i_11_1 ),
        .I1(\rgf_c1bus_wb[2]_i_7_2 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[11]_i_11_3 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_2 ),
        .O(\badr[10]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[14]_i_31 
       (.I0(\rgf_c1bus_wb[2]_i_7_2 ),
        .I1(\rgf_c1bus_wb[11]_i_11_1 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[2]_i_7 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[2]_i_7_0 ),
        .O(\badr[13]_INST_0_i_1 ));
  LUT5 #(
    .INIT(32'h44CF77CF)) 
    \rgf_c1bus_wb[14]_i_32 
       (.I0(\rgf_c1bus_wb[11]_i_8 ),
        .I1(\rgf_c1bus_wb[11]_i_11_0 ),
        .I2(\rgf_c1bus_wb[11]_i_8_0 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[10]_i_14_0 ),
        .O(\badr[2]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h030305F5F3F305F5)) 
    \rgf_c1bus_wb[14]_i_33 
       (.I0(\rgf_c1bus_wb[11]_i_8_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_0 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c0bus_wb[3]_i_7 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_8 ),
        .O(\sr_reg[6]_8 ));
  LUT6 #(
    .INIT(64'h5050303F5F5F303F)) 
    \rgf_c1bus_wb[15]_i_20 
       (.I0(\rgf_c1bus_wb[11]_i_8 ),
        .I1(\rgf_c1bus_wb[11]_i_8_0 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c0bus_wb[3]_i_7 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[2]_i_7_1 ),
        .O(\sr_reg[6]_10 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[15]_i_25 
       (.I0(\rgf_c1bus_wb[2]_i_7_0 ),
        .I1(\rgf_c1bus_wb[2]_i_7_2 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[2]_i_7_1 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[2]_i_7 ),
        .O(\badr[14]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_26 
       (.I0(\rgf_c1bus_wb[11]_i_11_3 ),
        .I1(\rgf_c1bus_wb[11]_i_11_4 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[11]_i_11_1 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_2 ),
        .O(\badr[10]_INST_0_i_1_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[1]_i_11 
       (.I0(\badr[10]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb[1]_i_3 ),
        .O(\rgf_c1bus_wb[9]_i_17 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[1]_i_4 
       (.I0(\rgf_c1bus_wb_reg[1] ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb_reg[1]_0 ),
        .O(\rgf_c1bus_wb[1]_i_14 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[3]_i_2 
       (.I0(\badr[5]_INST_0_i_1_0 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\badr[9]_INST_0_i_1 ),
        .I3(\rgf_c1bus_wb_reg[3] ),
        .O(\rgf_c1bus_wb[7]_i_4 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c1bus_wb[3]_i_6 
       (.I0(\rgf_c1bus_wb[11]_i_11_4 ),
        .I1(\rgf_c1bus_wb[11]_i_11_5 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[14]_i_3 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11 ),
        .O(\badr[5]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[4]_i_20 
       (.I0(\rgf_c1bus_wb[4]_i_7_1 ),
        .I1(\rgf_c1bus_wb[4]_i_7_2 ),
        .I2(\rgf_c1bus_wb[4]_i_7_3 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[4]_i_7_4 ),
        .I5(\rgf_c1bus_wb[4]_i_7_5 ),
        .O(\rgf_c1bus_wb[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h4C404C4C4C404040)) 
    \rgf_c1bus_wb[4]_i_3 
       (.I0(\rgf_c1bus_wb[4]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[4] ),
        .I2(\rgf_c1bus_wb_reg[5]_1 ),
        .I3(\badr[12]_INST_0_i_1 ),
        .I4(\rgf_c1bus_wb_reg[7] ),
        .I5(\rgf_c1bus_wb[14]_i_28_0 ),
        .O(\rgf_c1bus_wb[4]_i_9_0 ));
  LUT6 #(
    .INIT(64'hC0CFA0A0C0CFAFAF)) 
    \rgf_c1bus_wb[4]_i_7 
       (.I0(\rgf_c1bus_wb[4]_i_3_0 ),
        .I1(\rgf_c1bus_wb[4]_i_3_1 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .I3(\rgf_c1bus_wb[4]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11_0 ),
        .I5(\rgf_c1bus_wb[4]_i_3_2 ),
        .O(\rgf_c1bus_wb[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[4]_i_8 
       (.I0(\rgf_c1bus_wb[11]_i_11_1 ),
        .I1(\rgf_c1bus_wb[11]_i_11_2 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[2]_i_7_0 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[2]_i_7_2 ),
        .O(\badr[12]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \rgf_c1bus_wb[4]_i_9 
       (.I0(\rgf_c1bus_wb[11]_i_11_5 ),
        .I1(\rgf_c1bus_wb[14]_i_3 ),
        .I2(\rgf_c1bus_wb[11]_i_11_3 ),
        .I3(\rgf_c1bus_wb[4]_i_7_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11_4 ),
        .I5(\rgf_c1bus_wb[11]_i_11_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c1bus_wb[5]_i_13 
       (.I0(\tr_reg[5] ),
        .I1(\rgf_c1bus_wb[5]_i_10 ),
        .I2(\rgf_c1bus_wb[11]_i_11 ),
        .O(\badr[5]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hFCCCFCFFDDEEDDEE)) 
    \rgf_c1bus_wb[5]_i_14 
       (.I0(\rgf_c1bus_wb[11]_i_11 ),
        .I1(\rgf_c1bus_wb[5]_i_10 ),
        .I2(\tr_reg[5] ),
        .I3(\rgf_c1bus_wb[10]_i_14 ),
        .I4(\rgf_c1bus_wb[2]_i_7_0 ),
        .I5(\rgf_c1bus_wb_reg[5] ),
        .O(\stat_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hDFDCDFDFDCDCDCDF)) 
    \rgf_c1bus_wb[5]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_30_0 ),
        .I1(\rgf_c1bus_wb_reg[5]_0 ),
        .I2(\rgf_c1bus_wb_reg[5]_1 ),
        .I3(\rgf_c1bus_wb_reg[5] ),
        .I4(\sr_reg[6] ),
        .I5(\badr[15]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[13]_i_9_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c1bus_wb[6]_i_17 
       (.I0(\tr_reg[6] ),
        .I1(\rgf_c1bus_wb[5]_i_10 ),
        .I2(\rgf_c1bus_wb[14]_i_3 ),
        .O(\badr[6]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h000000005FC050CF)) 
    \rgf_c1bus_wb[6]_i_18 
       (.I0(\tr_reg[6] ),
        .I1(\rgf_c1bus_wb[2]_i_7 ),
        .I2(\rgf_c1bus_wb_reg[5] ),
        .I3(\rgf_c1bus_wb[10]_i_14 ),
        .I4(\rgf_c1bus_wb[14]_i_3 ),
        .I5(\rgf_c1bus_wb[5]_i_10 ),
        .O(\stat_reg[2] ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c1bus_wb[6]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_28_3 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\badr[2]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[14]_i_32_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[7]_i_10 
       (.I0(\rgf_c1bus_wb[3]_i_4 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\badr[14]_INST_0_i_1 ),
        .O(\rgf_c1bus_wb[11]_i_13_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[7]_i_3 
       (.I0(\badr[9]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\sr_reg[6]_1 ),
        .O(\sr_reg[6]_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[7]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_11 ),
        .I1(\rgf_c1bus_wb[11]_i_11_6 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[11]_i_11_5 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[14]_i_3 ),
        .O(\badr[6]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c1bus_wb[7]_i_8 
       (.I0(\rgf_c1bus_wb[2]_i_7_2 ),
        .I1(\rgf_c1bus_wb[11]_i_11_1 ),
        .I2(\rgf_c1bus_wb[11]_i_11_0 ),
        .I3(\rgf_c1bus_wb[11]_i_11_2 ),
        .I4(\rgf_c1bus_wb[4]_i_7_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_3 ),
        .O(\badr[9]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[8]_i_10 
       (.I0(\rgf_c1bus_wb[8]_i_3_0 ),
        .I1(\rgf_c1bus_wb[14]_i_28 ),
        .I2(\rgf_c1bus_wb_reg[7] ),
        .O(\rgf_c1bus_wb[11]_i_10 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[8]_i_11 
       (.I0(\rgf_c1bus_wb[3]_i_4_0 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb[8]_i_3 ),
        .I3(\rgf_c1bus_wb_reg[3] ),
        .O(\sr_reg[6]_2 ));
  LUT4 #(
    .INIT(16'h2EFF)) 
    \rgf_c1bus_wb[8]_i_8 
       (.I0(\badr[12]_INST_0_i_1 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\sr_reg[6]_9 ),
        .I3(\rgf_c1bus_wb_reg[3] ),
        .O(\sr_reg[6]_22 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \rgf_c1bus_wb[9]_i_16 
       (.I0(\rgf_c1bus_wb[2]_i_7_0 ),
        .I1(\rgf_c1bus_wb[4]_i_7_0 ),
        .I2(\rgf_c1bus_wb[2]_i_7 ),
        .I3(\rgf_c1bus_wb[11]_i_11_0 ),
        .I4(\rgf_c1bus_wb[2]_i_7_1 ),
        .O(\badr[15]_INST_0_i_1_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c1bus_wb[9]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_28_0 ),
        .I1(\rgf_c1bus_wb_reg[7] ),
        .I2(\rgf_c1bus_wb[14]_i_28_2 ),
        .O(\rgf_c1bus_wb[13]_i_16_0 ));
endmodule

module mcss_rgf_ivec
   (.out({iv[15],iv[14],iv[13],iv[12],iv[11],iv[10],iv[9],iv[8],iv[7],iv[6],iv[5],iv[4],iv[3],iv[2],iv[1],iv[0]}),
    SR,
    \iv_reg[15]_0 ,
    clk);
  input [0:0]SR;
  input [15:0]\iv_reg[15]_0 ;
  input clk;
     output [15:0]iv;

  wire \<const1> ;
  wire [0:0]SR;
  wire clk;
  (* DONT_TOUCH *) wire [15:0]iv;
  wire [15:0]\iv_reg[15]_0 ;

  VCC VCC
       (.P(\<const1> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [0]),
        .Q(iv[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [10]),
        .Q(iv[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [11]),
        .Q(iv[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [12]),
        .Q(iv[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [13]),
        .Q(iv[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [14]),
        .Q(iv[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [15]),
        .Q(iv[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [1]),
        .Q(iv[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [2]),
        .Q(iv[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [3]),
        .Q(iv[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [4]),
        .Q(iv[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [5]),
        .Q(iv[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [6]),
        .Q(iv[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [7]),
        .Q(iv[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [8]),
        .Q(iv[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\iv_reg[15]_0 [9]),
        .Q(iv[9]),
        .R(SR));
endmodule

module mcss_rgf_pcnt
   (.out({pc[15],pc[14],pc[13],pc[12],pc[11],pc[10],pc[9],pc[8],pc[7],pc[6],pc[5],pc[4],pc[3],pc[2],pc[1],pc[0]}),
    \pc_reg[15]_0 ,
    D,
    \pc_reg[14]_0 ,
    \pc_reg[13]_0 ,
    fadr,
    S,
    \pc_reg[1]_0 ,
    \pc_reg[15]_1 ,
    \pc_reg[13]_1 ,
    \pc0_reg[15] ,
    \fadr[15] ,
    O,
    \fadr[15]_0 ,
    \pc0_reg[15]_0 ,
    \pc0_reg[15]_1 ,
    \pc0_reg[15]_2 ,
    SR,
    \pc_reg[15]_2 ,
    clk);
  output \pc_reg[15]_0 ;
  output [2:0]D;
  output \pc_reg[14]_0 ;
  output \pc_reg[13]_0 ;
  output [2:0]fadr;
  output [0:0]S;
  output [0:0]\pc_reg[1]_0 ;
  output [2:0]\pc_reg[15]_1 ;
  input \pc_reg[13]_1 ;
  input [2:0]\pc0_reg[15] ;
  input \fadr[15] ;
  input [2:0]O;
  input \fadr[15]_0 ;
  input \pc0_reg[15]_0 ;
  input \pc0_reg[15]_1 ;
  input \pc0_reg[15]_2 ;
  input [0:0]SR;
  input [15:0]\pc_reg[15]_2 ;
  input clk;
     output [15:0]pc;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]O;
  wire [0:0]S;
  wire [0:0]SR;
  wire clk;
  wire [2:0]fadr;
  wire \fadr[15] ;
  wire \fadr[15]_0 ;
  (* DONT_TOUCH *) wire [15:0]pc;
  wire [2:0]\pc0_reg[15] ;
  wire \pc0_reg[15]_0 ;
  wire \pc0_reg[15]_1 ;
  wire \pc0_reg[15]_2 ;
  wire \pc_reg[13]_0 ;
  wire \pc_reg[13]_1 ;
  wire \pc_reg[14]_0 ;
  wire \pc_reg[15]_0 ;
  wire [2:0]\pc_reg[15]_1 ;
  wire [15:0]\pc_reg[15]_2 ;
  wire [0:0]\pc_reg[1]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[13]_INST_0 
       (.I0(\pc0_reg[15] [0]),
        .I1(\fadr[15] ),
        .I2(O[0]),
        .I3(\fadr[15]_0 ),
        .I4(pc[13]),
        .O(fadr[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[14]_INST_0 
       (.I0(\pc0_reg[15] [1]),
        .I1(\fadr[15] ),
        .I2(O[1]),
        .I3(\fadr[15]_0 ),
        .I4(pc[14]),
        .O(fadr[1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[15]_INST_0 
       (.I0(\pc0_reg[15] [2]),
        .I1(\fadr[15] ),
        .I2(O[2]),
        .I3(\fadr[15]_0 ),
        .I4(pc[15]),
        .O(fadr[2]));
  LUT1 #(
    .INIT(2'h1)) 
    fch_pc_nx2_carry_i_1
       (.I0(pc[1]),
        .O(\pc_reg[1]_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    fch_pc_nx4_carry_i_1
       (.I0(pc[2]),
        .O(S));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[13]_i_1 
       (.I0(\pc0_reg[15]_0 ),
        .I1(pc[13]),
        .I2(\pc0_reg[15]_1 ),
        .I3(\pc0_reg[15] [0]),
        .I4(\pc0_reg[15]_2 ),
        .I5(O[0]),
        .O(D[0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[14]_i_1 
       (.I0(\pc0_reg[15]_0 ),
        .I1(pc[14]),
        .I2(\pc0_reg[15]_1 ),
        .I3(\pc0_reg[15] [1]),
        .I4(\pc0_reg[15]_2 ),
        .I5(O[1]),
        .O(D[1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[15]_i_1 
       (.I0(\pc0_reg[15]_0 ),
        .I1(pc[15]),
        .I2(\pc0_reg[15]_1 ),
        .I3(\pc0_reg[15] [2]),
        .I4(\pc0_reg[15]_2 ),
        .I5(O[2]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_1
       (.I0(\pc0_reg[15]_0 ),
        .I1(pc[15]),
        .I2(\pc0_reg[15]_1 ),
        .I3(\pc0_reg[15] [2]),
        .I4(\pc0_reg[15]_2 ),
        .I5(O[2]),
        .O(\pc_reg[15]_1 [2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_2
       (.I0(\pc0_reg[15]_0 ),
        .I1(pc[14]),
        .I2(\pc0_reg[15]_1 ),
        .I3(\pc0_reg[15] [1]),
        .I4(\pc0_reg[15]_2 ),
        .I5(O[1]),
        .O(\pc_reg[15]_1 [1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_3
       (.I0(\pc0_reg[15]_0 ),
        .I1(pc[13]),
        .I2(\pc0_reg[15]_1 ),
        .I3(\pc0_reg[15] [0]),
        .I4(\pc0_reg[15]_2 ),
        .I5(O[0]),
        .O(\pc_reg[15]_1 [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[13]_i_4 
       (.I0(D[0]),
        .I1(\pc_reg[13]_1 ),
        .I2(pc[13]),
        .O(\pc_reg[13]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[14]_i_4 
       (.I0(D[1]),
        .I1(\pc_reg[13]_1 ),
        .I2(pc[14]),
        .O(\pc_reg[14]_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[15]_i_6 
       (.I0(D[2]),
        .I1(\pc_reg[13]_1 ),
        .I2(pc[15]),
        .O(\pc_reg[15]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [0]),
        .Q(pc[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [10]),
        .Q(pc[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [11]),
        .Q(pc[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [12]),
        .Q(pc[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [13]),
        .Q(pc[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [14]),
        .Q(pc[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [15]),
        .Q(pc[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [1]),
        .Q(pc[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [2]),
        .Q(pc[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [3]),
        .Q(pc[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [4]),
        .Q(pc[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [5]),
        .Q(pc[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [6]),
        .Q(pc[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [7]),
        .Q(pc[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [8]),
        .Q(pc[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_2 [9]),
        .Q(pc[9]),
        .R(SR));
endmodule

module mcss_rgf_sptr
   (.out({sp[15],sp[14],sp[13],sp[12],sp[11],sp[10],sp[9],sp[8],sp[7],sp[6],sp[5],sp[4],sp[3],sp[2],sp[1],sp[0]}),
    O,
    data3,
    \sp_reg[15]_0 ,
    \sp_reg[1]_0 ,
    \sp_reg[2]_0 ,
    \sp_reg[3]_0 ,
    \sp_reg[4]_0 ,
    \sp_reg[5]_0 ,
    \sp_reg[6]_0 ,
    \sp_reg[7]_0 ,
    \sp_reg[8]_0 ,
    \sp_reg[9]_0 ,
    \sp_reg[10]_0 ,
    \sp_reg[11]_0 ,
    \sp_reg[12]_0 ,
    \sp_reg[13]_0 ,
    \sp_reg[14]_0 ,
    \sp_reg[14]_1 ,
    \sp_reg[14]_2 ,
    SR,
    \sp_reg[15]_1 ,
    clk);
  output [0:0]O;
  output [14:0]data3;
  output \sp_reg[15]_0 ;
  output \sp_reg[1]_0 ;
  output \sp_reg[2]_0 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[4]_0 ;
  output \sp_reg[5]_0 ;
  output \sp_reg[6]_0 ;
  output \sp_reg[7]_0 ;
  output \sp_reg[8]_0 ;
  output \sp_reg[9]_0 ;
  output \sp_reg[10]_0 ;
  output \sp_reg[11]_0 ;
  output \sp_reg[12]_0 ;
  output \sp_reg[13]_0 ;
  output \sp_reg[14]_0 ;
  input \sp_reg[14]_1 ;
  input \sp_reg[14]_2 ;
  input [0:0]SR;
  input [15:0]\sp_reg[15]_1 ;
  input clk;
     output [15:0]sp;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]O;
  wire [0:0]SR;
  wire \badr[0]_INST_0_i_24_n_0 ;
  wire \badr[0]_INST_0_i_24_n_1 ;
  wire \badr[0]_INST_0_i_24_n_2 ;
  wire \badr[0]_INST_0_i_24_n_3 ;
  wire \badr[0]_INST_0_i_37_n_0 ;
  wire \badr[11]_INST_0_i_24_n_0 ;
  wire \badr[11]_INST_0_i_24_n_1 ;
  wire \badr[11]_INST_0_i_24_n_2 ;
  wire \badr[11]_INST_0_i_24_n_3 ;
  wire \badr[11]_INST_0_i_37_n_0 ;
  wire \badr[11]_INST_0_i_38_n_0 ;
  wire \badr[11]_INST_0_i_39_n_0 ;
  wire \badr[11]_INST_0_i_40_n_0 ;
  wire \badr[15]_INST_0_i_103_n_0 ;
  wire \badr[15]_INST_0_i_104_n_0 ;
  wire \badr[15]_INST_0_i_105_n_0 ;
  wire \badr[15]_INST_0_i_106_n_0 ;
  wire \badr[15]_INST_0_i_36_n_1 ;
  wire \badr[15]_INST_0_i_36_n_2 ;
  wire \badr[15]_INST_0_i_36_n_3 ;
  wire \badr[3]_INST_0_i_24_n_0 ;
  wire \badr[3]_INST_0_i_24_n_1 ;
  wire \badr[3]_INST_0_i_24_n_2 ;
  wire \badr[3]_INST_0_i_24_n_3 ;
  wire \badr[3]_INST_0_i_37_n_0 ;
  wire \badr[3]_INST_0_i_38_n_0 ;
  wire \badr[3]_INST_0_i_39_n_0 ;
  wire \badr[7]_INST_0_i_24_n_0 ;
  wire \badr[7]_INST_0_i_24_n_1 ;
  wire \badr[7]_INST_0_i_24_n_2 ;
  wire \badr[7]_INST_0_i_24_n_3 ;
  wire \badr[7]_INST_0_i_37_n_0 ;
  wire \badr[7]_INST_0_i_38_n_0 ;
  wire \badr[7]_INST_0_i_39_n_0 ;
  wire \badr[7]_INST_0_i_40_n_0 ;
  wire clk;
  wire [15:1]data2;
  wire [14:0]data3;
  (* DONT_TOUCH *) wire [15:0]sp;
  wire \sp_reg[10]_0 ;
  wire \sp_reg[11]_0 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[12]_0 ;
  wire \sp_reg[13]_0 ;
  wire \sp_reg[14]_0 ;
  wire \sp_reg[14]_1 ;
  wire \sp_reg[14]_2 ;
  wire \sp_reg[15]_0 ;
  wire [15:0]\sp_reg[15]_1 ;
  wire \sp_reg[15]_i_7_n_1 ;
  wire \sp_reg[15]_i_7_n_2 ;
  wire \sp_reg[15]_i_7_n_3 ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[5]_0 ;
  wire \sp_reg[6]_0 ;
  wire \sp_reg[7]_0 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sp_reg[8]_0 ;
  wire \sp_reg[9]_0 ;
  wire [3:0]\NLW_badr[3]_INST_0_i_24_O_UNCONNECTED ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[0]_INST_0_i_24 
       (.CI(\<const0> ),
        .CO({\badr[0]_INST_0_i_24_n_0 ,\badr[0]_INST_0_i_24_n_1 ,\badr[0]_INST_0_i_24_n_2 ,\badr[0]_INST_0_i_24_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,sp[1],\<const0> }),
        .O({data2[3:1],O}),
        .S({sp[3:2],\badr[0]_INST_0_i_37_n_0 ,sp[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[0]_INST_0_i_37 
       (.I0(sp[1]),
        .O(\badr[0]_INST_0_i_37_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[11]_INST_0_i_24 
       (.CI(\badr[7]_INST_0_i_24_n_0 ),
        .CO({\badr[11]_INST_0_i_24_n_0 ,\badr[11]_INST_0_i_24_n_1 ,\badr[11]_INST_0_i_24_n_2 ,\badr[11]_INST_0_i_24_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[11:8]),
        .O(data3[10:7]),
        .S({\badr[11]_INST_0_i_37_n_0 ,\badr[11]_INST_0_i_38_n_0 ,\badr[11]_INST_0_i_39_n_0 ,\badr[11]_INST_0_i_40_n_0 }));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_37 
       (.I0(sp[11]),
        .O(\badr[11]_INST_0_i_37_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_38 
       (.I0(sp[10]),
        .O(\badr[11]_INST_0_i_38_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_39 
       (.I0(sp[9]),
        .O(\badr[11]_INST_0_i_39_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_40 
       (.I0(sp[8]),
        .O(\badr[11]_INST_0_i_40_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_103 
       (.I0(sp[15]),
        .O(\badr[15]_INST_0_i_103_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_104 
       (.I0(sp[14]),
        .O(\badr[15]_INST_0_i_104_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_105 
       (.I0(sp[13]),
        .O(\badr[15]_INST_0_i_105_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_106 
       (.I0(sp[12]),
        .O(\badr[15]_INST_0_i_106_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[15]_INST_0_i_36 
       (.CI(\badr[11]_INST_0_i_24_n_0 ),
        .CO({\badr[15]_INST_0_i_36_n_1 ,\badr[15]_INST_0_i_36_n_2 ,\badr[15]_INST_0_i_36_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,sp[14:12]}),
        .O(data3[14:11]),
        .S({\badr[15]_INST_0_i_103_n_0 ,\badr[15]_INST_0_i_104_n_0 ,\badr[15]_INST_0_i_105_n_0 ,\badr[15]_INST_0_i_106_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[3]_INST_0_i_24 
       (.CI(\<const0> ),
        .CO({\badr[3]_INST_0_i_24_n_0 ,\badr[3]_INST_0_i_24_n_1 ,\badr[3]_INST_0_i_24_n_2 ,\badr[3]_INST_0_i_24_n_3 }),
        .CYINIT(\<const0> ),
        .DI({sp[3:1],\<const0> }),
        .O({data3[2:0],\NLW_badr[3]_INST_0_i_24_O_UNCONNECTED [0]}),
        .S({\badr[3]_INST_0_i_37_n_0 ,\badr[3]_INST_0_i_38_n_0 ,\badr[3]_INST_0_i_39_n_0 ,sp[0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_37 
       (.I0(sp[3]),
        .O(\badr[3]_INST_0_i_37_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_38 
       (.I0(sp[2]),
        .O(\badr[3]_INST_0_i_38_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_39 
       (.I0(sp[1]),
        .O(\badr[3]_INST_0_i_39_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[7]_INST_0_i_24 
       (.CI(\badr[3]_INST_0_i_24_n_0 ),
        .CO({\badr[7]_INST_0_i_24_n_0 ,\badr[7]_INST_0_i_24_n_1 ,\badr[7]_INST_0_i_24_n_2 ,\badr[7]_INST_0_i_24_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[7:4]),
        .O(data3[6:3]),
        .S({\badr[7]_INST_0_i_37_n_0 ,\badr[7]_INST_0_i_38_n_0 ,\badr[7]_INST_0_i_39_n_0 ,\badr[7]_INST_0_i_40_n_0 }));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_37 
       (.I0(sp[7]),
        .O(\badr[7]_INST_0_i_37_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_38 
       (.I0(sp[6]),
        .O(\badr[7]_INST_0_i_38_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_39 
       (.I0(sp[5]),
        .O(\badr[7]_INST_0_i_39_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_40 
       (.I0(sp[4]),
        .O(\badr[7]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[10]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[9]),
        .I2(sp[10]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[10]),
        .O(\sp_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[11]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[10]),
        .I2(sp[11]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[11]),
        .O(\sp_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[12]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[11]),
        .I2(sp[12]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[12]),
        .O(\sp_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[13]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[12]),
        .I2(sp[13]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[13]),
        .O(\sp_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[14]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[13]),
        .I2(sp[14]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[14]),
        .O(\sp_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[15]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[14]),
        .I2(sp[15]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[15]),
        .O(\sp_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[1]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[0]),
        .I2(sp[1]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[1]),
        .O(\sp_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[2]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[1]),
        .I2(sp[2]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[2]),
        .O(\sp_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[3]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[2]),
        .I2(sp[3]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[3]),
        .O(\sp_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[4]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[3]),
        .I2(sp[4]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[4]),
        .O(\sp_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[5]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[4]),
        .I2(sp[5]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[5]),
        .O(\sp_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[6]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[5]),
        .I2(sp[6]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[6]),
        .O(\sp_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[7]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[6]),
        .I2(sp[7]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[7]),
        .O(\sp_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[8]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[7]),
        .I2(sp[8]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[8]),
        .O(\sp_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[9]_i_2 
       (.I0(\sp_reg[14]_1 ),
        .I1(data3[8]),
        .I2(sp[9]),
        .I3(\sp_reg[14]_2 ),
        .I4(data2[9]),
        .O(\sp_reg[9]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [0]),
        .Q(sp[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [10]),
        .Q(sp[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [11]),
        .Q(sp[11]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[11:8]),
        .S(sp[11:8]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [12]),
        .Q(sp[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [13]),
        .Q(sp[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [14]),
        .Q(sp[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [15]),
        .Q(sp[15]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_7 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_7_n_1 ,\sp_reg[15]_i_7_n_2 ,\sp_reg[15]_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[15:12]),
        .S(sp[15:12]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [1]),
        .Q(sp[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [2]),
        .Q(sp[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [3]),
        .Q(sp[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [4]),
        .Q(sp[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [5]),
        .Q(sp[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [6]),
        .Q(sp[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [7]),
        .Q(sp[7]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\badr[0]_INST_0_i_24_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(data2[7:4]),
        .S(sp[7:4]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [8]),
        .Q(sp[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[15]_1 [9]),
        .Q(sp[9]),
        .R(SR));
endmodule

module mcss_rgf_sreg
   (.\sr_reg[15]_0 ({sr[15],sr[14],sr[13],sr[12],sr[11],sr[10],sr[9],sr[8],sr[7],sr[6],sr[5],sr[4],sr[3],sr[2],sr[1],sr[0]}),
    \sr_reg[4]_0 ,
    \sr_reg[5]_0 ,
    \sr_reg[6]_0 ,
    \sr_reg[6]_1 ,
    \sr_reg[6]_2 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    \sr_reg[4]_1 ,
    \sr_reg[5]_1 ,
    \sr_reg[7]_0 ,
    \sr_reg[5]_2 ,
    \sr_reg[6]_5 ,
    \sr_reg[5]_3 ,
    \sr_reg[6]_6 ,
    irq_0,
    fch_irq_req,
    \sr_reg[10]_0 ,
    \sr_reg[4]_2 ,
    \sr_reg[0]_0 ,
    \sr_reg[0]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[0]_5 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[0]_11 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[0]_17 ,
    \sr_reg[0]_18 ,
    \sr_reg[0]_19 ,
    \sr_reg[0]_20 ,
    \sr_reg[1]_0 ,
    \sr_reg[1]_1 ,
    \sr_reg[1]_2 ,
    \sr_reg[1]_3 ,
    \sr_reg[1]_4 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[0]_23 ,
    \sr_reg[0]_24 ,
    \sr_reg[0]_25 ,
    \sr_reg[0]_26 ,
    \sr_reg[0]_27 ,
    \sr_reg[0]_28 ,
    \sr_reg[0]_29 ,
    \sr_reg[0]_30 ,
    \sr_reg[0]_31 ,
    \sr_reg[0]_32 ,
    \sr_reg[0]_33 ,
    \sr_reg[0]_34 ,
    \sr_reg[0]_35 ,
    \sr_reg[0]_36 ,
    \sr_reg[1]_5 ,
    \sr_reg[1]_6 ,
    \sr_reg[1]_7 ,
    \sr_reg[1]_8 ,
    \sr_reg[1]_9 ,
    \sr_reg[1]_10 ,
    \sr_reg[1]_11 ,
    \sr_reg[1]_12 ,
    \sr_reg[1]_13 ,
    \sr_reg[1]_14 ,
    \sr_reg[1]_15 ,
    \sr_reg[1]_16 ,
    \sr_reg[1]_17 ,
    \sr_reg[1]_18 ,
    \sr_reg[1]_19 ,
    \sr_reg[5]_4 ,
    \sr_reg[5]_5 ,
    \sr_reg[5]_6 ,
    \sr_reg[0]_37 ,
    \sr_reg[1]_20 ,
    \sr_reg[1]_21 ,
    \sr_reg[1]_22 ,
    \sr_reg[1]_23 ,
    \sr_reg[1]_24 ,
    \sr_reg[1]_25 ,
    \sr_reg[1]_26 ,
    \sr_reg[1]_27 ,
    \sr_reg[1]_28 ,
    \sr_reg[1]_29 ,
    \sr_reg[1]_30 ,
    \sr_reg[1]_31 ,
    \sr_reg[1]_32 ,
    \sr_reg[1]_33 ,
    \sr_reg[1]_34 ,
    \sr_reg[1]_35 ,
    \sr_reg[1]_36 ,
    \sr_reg[0]_38 ,
    \sr_reg[0]_39 ,
    \sr_reg[0]_40 ,
    \sr_reg[0]_41 ,
    \sr_reg[0]_42 ,
    \sr_reg[0]_43 ,
    \sr_reg[0]_44 ,
    \sr_reg[0]_45 ,
    \sr_reg[0]_46 ,
    \sr_reg[0]_47 ,
    \sr_reg[0]_48 ,
    \sr_reg[0]_49 ,
    \sr_reg[0]_50 ,
    \sr_reg[0]_51 ,
    \sr_reg[0]_52 ,
    \sr_reg[0]_53 ,
    \sr_reg[1]_37 ,
    \sr_reg[1]_38 ,
    \sr_reg[1]_39 ,
    \sr_reg[1]_40 ,
    \sr_reg[1]_41 ,
    \sr_reg[1]_42 ,
    \sr_reg[1]_43 ,
    \sr_reg[1]_44 ,
    \sr_reg[1]_45 ,
    \sr_reg[1]_46 ,
    \sr_reg[1]_47 ,
    \sr_reg[1]_48 ,
    \sr_reg[1]_49 ,
    \sr_reg[1]_50 ,
    \sr_reg[1]_51 ,
    \sr_reg[1]_52 ,
    \sr_reg[1]_53 ,
    \sr_reg[1]_54 ,
    \sr_reg[1]_55 ,
    \sr_reg[1]_56 ,
    \sr_reg[1]_57 ,
    \sr_reg[1]_58 ,
    \sr_reg[1]_59 ,
    \sr_reg[1]_60 ,
    \sr_reg[1]_61 ,
    \sr_reg[1]_62 ,
    \sr_reg[1]_63 ,
    \sr_reg[1]_64 ,
    \sr_reg[1]_65 ,
    \sr_reg[1]_66 ,
    \sr_reg[1]_67 ,
    \sr_reg[1]_68 ,
    \sr_reg[5]_7 ,
    \sr[4]_i_160 ,
    \sr[4]_i_160_0 ,
    \sr[4]_i_160_1 ,
    \sr[4]_i_160_2 ,
    \sr[4]_i_160_3 ,
    \sr[4]_i_172 ,
    \sr[4]_i_172_0 ,
    \sr[4]_i_172_1 ,
    \sr[4]_i_172_2 ,
    \sr[4]_i_188 ,
    \sr[4]_i_188_0 ,
    \sr[4]_i_188_1 ,
    \sr[4]_i_188_2 ,
    \rgf_c0bus_wb[4]_i_10 ,
    \rgf_c0bus_wb[4]_i_10_0 ,
    \rgf_c0bus_wb[4]_i_10_1 ,
    \rgf_c0bus_wb[0]_i_5 ,
    \badr[15]_INST_0_i_208 ,
    \rgf_selc1_wb[1]_i_16 ,
    irq,
    irq_lev,
    Q,
    ctl_fetch1_fl_i_15,
    b0bus_sel_0,
    \i_/bbus_o[4]_INST_0_i_5 ,
    a1bus_sel_0,
    \badr[15]_INST_0_i_7 ,
    \i_/bbus_o[4]_INST_0_i_6 ,
    \rgf_c1bus_wb[4]_i_45 ,
    \rgf_c1bus_wb[4]_i_39 ,
    \rgf_c1bus_wb[4]_i_47 ,
    \rgf_c1bus_wb[4]_i_47_0 ,
    \rgf_c1bus_wb[4]_i_39_0 ,
    gr6_bus1,
    \rgf_c1bus_wb[4]_i_45_0 ,
    gr6_bus1_0,
    \badr[15]_INST_0_i_7_0 ,
    gr6_bus1_1,
    \sr_reg[15]_1 ,
    clk);
  output \sr_reg[4]_0 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[6]_4 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[5]_1 ;
  output \sr_reg[7]_0 ;
  output \sr_reg[5]_2 ;
  output \sr_reg[6]_5 ;
  output \sr_reg[5]_3 ;
  output \sr_reg[6]_6 ;
  output irq_0;
  output fch_irq_req;
  output \sr_reg[10]_0 ;
  output \sr_reg[4]_2 ;
  output \sr_reg[0]_0 ;
  output \sr_reg[0]_1 ;
  output \sr_reg[0]_2 ;
  output \sr_reg[0]_3 ;
  output \sr_reg[0]_4 ;
  output \sr_reg[0]_5 ;
  output \sr_reg[0]_6 ;
  output \sr_reg[0]_7 ;
  output \sr_reg[0]_8 ;
  output \sr_reg[0]_9 ;
  output \sr_reg[0]_10 ;
  output \sr_reg[0]_11 ;
  output \sr_reg[0]_12 ;
  output \sr_reg[0]_13 ;
  output \sr_reg[0]_14 ;
  output \sr_reg[0]_15 ;
  output \sr_reg[0]_16 ;
  output \sr_reg[0]_17 ;
  output \sr_reg[0]_18 ;
  output \sr_reg[0]_19 ;
  output \sr_reg[0]_20 ;
  output \sr_reg[1]_0 ;
  output \sr_reg[1]_1 ;
  output \sr_reg[1]_2 ;
  output \sr_reg[1]_3 ;
  output \sr_reg[1]_4 ;
  output \sr_reg[0]_21 ;
  output \sr_reg[0]_22 ;
  output \sr_reg[0]_23 ;
  output \sr_reg[0]_24 ;
  output \sr_reg[0]_25 ;
  output \sr_reg[0]_26 ;
  output \sr_reg[0]_27 ;
  output \sr_reg[0]_28 ;
  output \sr_reg[0]_29 ;
  output \sr_reg[0]_30 ;
  output \sr_reg[0]_31 ;
  output \sr_reg[0]_32 ;
  output \sr_reg[0]_33 ;
  output \sr_reg[0]_34 ;
  output \sr_reg[0]_35 ;
  output \sr_reg[0]_36 ;
  output \sr_reg[1]_5 ;
  output \sr_reg[1]_6 ;
  output \sr_reg[1]_7 ;
  output \sr_reg[1]_8 ;
  output \sr_reg[1]_9 ;
  output \sr_reg[1]_10 ;
  output \sr_reg[1]_11 ;
  output \sr_reg[1]_12 ;
  output \sr_reg[1]_13 ;
  output \sr_reg[1]_14 ;
  output \sr_reg[1]_15 ;
  output \sr_reg[1]_16 ;
  output \sr_reg[1]_17 ;
  output \sr_reg[1]_18 ;
  output \sr_reg[1]_19 ;
  output \sr_reg[5]_4 ;
  output \sr_reg[5]_5 ;
  output \sr_reg[5]_6 ;
  output \sr_reg[0]_37 ;
  output \sr_reg[1]_20 ;
  output \sr_reg[1]_21 ;
  output \sr_reg[1]_22 ;
  output \sr_reg[1]_23 ;
  output \sr_reg[1]_24 ;
  output \sr_reg[1]_25 ;
  output \sr_reg[1]_26 ;
  output \sr_reg[1]_27 ;
  output \sr_reg[1]_28 ;
  output \sr_reg[1]_29 ;
  output \sr_reg[1]_30 ;
  output \sr_reg[1]_31 ;
  output \sr_reg[1]_32 ;
  output \sr_reg[1]_33 ;
  output \sr_reg[1]_34 ;
  output \sr_reg[1]_35 ;
  output \sr_reg[1]_36 ;
  output \sr_reg[0]_38 ;
  output \sr_reg[0]_39 ;
  output \sr_reg[0]_40 ;
  output \sr_reg[0]_41 ;
  output \sr_reg[0]_42 ;
  output \sr_reg[0]_43 ;
  output \sr_reg[0]_44 ;
  output \sr_reg[0]_45 ;
  output \sr_reg[0]_46 ;
  output \sr_reg[0]_47 ;
  output \sr_reg[0]_48 ;
  output \sr_reg[0]_49 ;
  output \sr_reg[0]_50 ;
  output \sr_reg[0]_51 ;
  output \sr_reg[0]_52 ;
  output \sr_reg[0]_53 ;
  output \sr_reg[1]_37 ;
  output \sr_reg[1]_38 ;
  output \sr_reg[1]_39 ;
  output \sr_reg[1]_40 ;
  output \sr_reg[1]_41 ;
  output \sr_reg[1]_42 ;
  output \sr_reg[1]_43 ;
  output \sr_reg[1]_44 ;
  output \sr_reg[1]_45 ;
  output \sr_reg[1]_46 ;
  output \sr_reg[1]_47 ;
  output \sr_reg[1]_48 ;
  output \sr_reg[1]_49 ;
  output \sr_reg[1]_50 ;
  output \sr_reg[1]_51 ;
  output \sr_reg[1]_52 ;
  output \sr_reg[1]_53 ;
  output \sr_reg[1]_54 ;
  output \sr_reg[1]_55 ;
  output \sr_reg[1]_56 ;
  output \sr_reg[1]_57 ;
  output \sr_reg[1]_58 ;
  output \sr_reg[1]_59 ;
  output \sr_reg[1]_60 ;
  output \sr_reg[1]_61 ;
  output \sr_reg[1]_62 ;
  output \sr_reg[1]_63 ;
  output \sr_reg[1]_64 ;
  output \sr_reg[1]_65 ;
  output \sr_reg[1]_66 ;
  output \sr_reg[1]_67 ;
  output \sr_reg[1]_68 ;
  input \sr_reg[5]_7 ;
  input \sr[4]_i_160 ;
  input \sr[4]_i_160_0 ;
  input [0:0]\sr[4]_i_160_1 ;
  input \sr[4]_i_160_2 ;
  input \sr[4]_i_160_3 ;
  input \sr[4]_i_172 ;
  input [0:0]\sr[4]_i_172_0 ;
  input \sr[4]_i_172_1 ;
  input \sr[4]_i_172_2 ;
  input \sr[4]_i_188 ;
  input \sr[4]_i_188_0 ;
  input \sr[4]_i_188_1 ;
  input \sr[4]_i_188_2 ;
  input \rgf_c0bus_wb[4]_i_10 ;
  input \rgf_c0bus_wb[4]_i_10_0 ;
  input \rgf_c0bus_wb[4]_i_10_1 ;
  input \rgf_c0bus_wb[0]_i_5 ;
  input [4:0]\badr[15]_INST_0_i_208 ;
  input [3:0]\rgf_selc1_wb[1]_i_16 ;
  input irq;
  input [1:0]irq_lev;
  input [0:0]Q;
  input ctl_fetch1_fl_i_15;
  input [0:0]b0bus_sel_0;
  input [4:0]\i_/bbus_o[4]_INST_0_i_5 ;
  input [1:0]a1bus_sel_0;
  input [15:0]\badr[15]_INST_0_i_7 ;
  input [4:0]\i_/bbus_o[4]_INST_0_i_6 ;
  input [15:0]\rgf_c1bus_wb[4]_i_45 ;
  input [15:0]\rgf_c1bus_wb[4]_i_39 ;
  input [15:0]\rgf_c1bus_wb[4]_i_47 ;
  input [15:0]\rgf_c1bus_wb[4]_i_47_0 ;
  input [15:0]\rgf_c1bus_wb[4]_i_39_0 ;
  input gr6_bus1;
  input [15:0]\rgf_c1bus_wb[4]_i_45_0 ;
  input gr6_bus1_0;
  input [15:0]\badr[15]_INST_0_i_7_0 ;
  input gr6_bus1_1;
  input [15:0]\sr_reg[15]_1 ;
  input clk;
     output [15:0]sr;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]Q;
  wire [1:0]a1bus_sel_0;
  wire [0:0]b0bus_sel_0;
  wire [4:0]\badr[15]_INST_0_i_208 ;
  wire [15:0]\badr[15]_INST_0_i_7 ;
  wire [15:0]\badr[15]_INST_0_i_7_0 ;
  wire clk;
  wire ctl_fetch1_fl_i_15;
  wire ctl_fetch1_fl_i_38_n_0;
  wire fch_irq_req;
  wire gr6_bus1;
  wire gr6_bus1_0;
  wire gr6_bus1_1;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_5 ;
  wire [4:0]\i_/bbus_o[4]_INST_0_i_6 ;
  wire irq;
  wire irq_0;
  wire [1:0]irq_lev;
  wire \rgf_c0bus_wb[0]_i_5 ;
  wire \rgf_c0bus_wb[4]_i_10 ;
  wire \rgf_c0bus_wb[4]_i_10_0 ;
  wire \rgf_c0bus_wb[4]_i_10_1 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_39 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_39_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_45_0 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_47 ;
  wire [15:0]\rgf_c1bus_wb[4]_i_47_0 ;
  wire [3:0]\rgf_selc1_wb[1]_i_16 ;
  (* DONT_TOUCH *) wire [15:0]sr;
  wire \sr[4]_i_160 ;
  wire \sr[4]_i_160_0 ;
  wire [0:0]\sr[4]_i_160_1 ;
  wire \sr[4]_i_160_2 ;
  wire \sr[4]_i_160_3 ;
  wire \sr[4]_i_172 ;
  wire [0:0]\sr[4]_i_172_0 ;
  wire \sr[4]_i_172_1 ;
  wire \sr[4]_i_172_2 ;
  wire \sr[4]_i_188 ;
  wire \sr[4]_i_188_0 ;
  wire \sr[4]_i_188_1 ;
  wire \sr[4]_i_188_2 ;
  wire \sr_reg[0]_0 ;
  wire \sr_reg[0]_1 ;
  wire \sr_reg[0]_10 ;
  wire \sr_reg[0]_11 ;
  wire \sr_reg[0]_12 ;
  wire \sr_reg[0]_13 ;
  wire \sr_reg[0]_14 ;
  wire \sr_reg[0]_15 ;
  wire \sr_reg[0]_16 ;
  wire \sr_reg[0]_17 ;
  wire \sr_reg[0]_18 ;
  wire \sr_reg[0]_19 ;
  wire \sr_reg[0]_2 ;
  wire \sr_reg[0]_20 ;
  wire \sr_reg[0]_21 ;
  wire \sr_reg[0]_22 ;
  wire \sr_reg[0]_23 ;
  wire \sr_reg[0]_24 ;
  wire \sr_reg[0]_25 ;
  wire \sr_reg[0]_26 ;
  wire \sr_reg[0]_27 ;
  wire \sr_reg[0]_28 ;
  wire \sr_reg[0]_29 ;
  wire \sr_reg[0]_3 ;
  wire \sr_reg[0]_30 ;
  wire \sr_reg[0]_31 ;
  wire \sr_reg[0]_32 ;
  wire \sr_reg[0]_33 ;
  wire \sr_reg[0]_34 ;
  wire \sr_reg[0]_35 ;
  wire \sr_reg[0]_36 ;
  wire \sr_reg[0]_37 ;
  wire \sr_reg[0]_38 ;
  wire \sr_reg[0]_39 ;
  wire \sr_reg[0]_4 ;
  wire \sr_reg[0]_40 ;
  wire \sr_reg[0]_41 ;
  wire \sr_reg[0]_42 ;
  wire \sr_reg[0]_43 ;
  wire \sr_reg[0]_44 ;
  wire \sr_reg[0]_45 ;
  wire \sr_reg[0]_46 ;
  wire \sr_reg[0]_47 ;
  wire \sr_reg[0]_48 ;
  wire \sr_reg[0]_49 ;
  wire \sr_reg[0]_5 ;
  wire \sr_reg[0]_50 ;
  wire \sr_reg[0]_51 ;
  wire \sr_reg[0]_52 ;
  wire \sr_reg[0]_53 ;
  wire \sr_reg[0]_6 ;
  wire \sr_reg[0]_7 ;
  wire \sr_reg[0]_8 ;
  wire \sr_reg[0]_9 ;
  wire \sr_reg[10]_0 ;
  wire [15:0]\sr_reg[15]_1 ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[1]_1 ;
  wire \sr_reg[1]_10 ;
  wire \sr_reg[1]_11 ;
  wire \sr_reg[1]_12 ;
  wire \sr_reg[1]_13 ;
  wire \sr_reg[1]_14 ;
  wire \sr_reg[1]_15 ;
  wire \sr_reg[1]_16 ;
  wire \sr_reg[1]_17 ;
  wire \sr_reg[1]_18 ;
  wire \sr_reg[1]_19 ;
  wire \sr_reg[1]_2 ;
  wire \sr_reg[1]_20 ;
  wire \sr_reg[1]_21 ;
  wire \sr_reg[1]_22 ;
  wire \sr_reg[1]_23 ;
  wire \sr_reg[1]_24 ;
  wire \sr_reg[1]_25 ;
  wire \sr_reg[1]_26 ;
  wire \sr_reg[1]_27 ;
  wire \sr_reg[1]_28 ;
  wire \sr_reg[1]_29 ;
  wire \sr_reg[1]_3 ;
  wire \sr_reg[1]_30 ;
  wire \sr_reg[1]_31 ;
  wire \sr_reg[1]_32 ;
  wire \sr_reg[1]_33 ;
  wire \sr_reg[1]_34 ;
  wire \sr_reg[1]_35 ;
  wire \sr_reg[1]_36 ;
  wire \sr_reg[1]_37 ;
  wire \sr_reg[1]_38 ;
  wire \sr_reg[1]_39 ;
  wire \sr_reg[1]_4 ;
  wire \sr_reg[1]_40 ;
  wire \sr_reg[1]_41 ;
  wire \sr_reg[1]_42 ;
  wire \sr_reg[1]_43 ;
  wire \sr_reg[1]_44 ;
  wire \sr_reg[1]_45 ;
  wire \sr_reg[1]_46 ;
  wire \sr_reg[1]_47 ;
  wire \sr_reg[1]_48 ;
  wire \sr_reg[1]_49 ;
  wire \sr_reg[1]_5 ;
  wire \sr_reg[1]_50 ;
  wire \sr_reg[1]_51 ;
  wire \sr_reg[1]_52 ;
  wire \sr_reg[1]_53 ;
  wire \sr_reg[1]_54 ;
  wire \sr_reg[1]_55 ;
  wire \sr_reg[1]_56 ;
  wire \sr_reg[1]_57 ;
  wire \sr_reg[1]_58 ;
  wire \sr_reg[1]_59 ;
  wire \sr_reg[1]_6 ;
  wire \sr_reg[1]_60 ;
  wire \sr_reg[1]_61 ;
  wire \sr_reg[1]_62 ;
  wire \sr_reg[1]_63 ;
  wire \sr_reg[1]_64 ;
  wire \sr_reg[1]_65 ;
  wire \sr_reg[1]_66 ;
  wire \sr_reg[1]_67 ;
  wire \sr_reg[1]_68 ;
  wire \sr_reg[1]_7 ;
  wire \sr_reg[1]_8 ;
  wire \sr_reg[1]_9 ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[5]_3 ;
  wire \sr_reg[5]_4 ;
  wire \sr_reg[5]_5 ;
  wire \sr_reg[5]_6 ;
  wire \sr_reg[5]_7 ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[7]_0 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[0]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [0]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [0]),
        .O(\sr_reg[1]_36 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[0]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [0]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [0]),
        .O(\sr_reg[0]_38 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[0]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [0]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [0]),
        .O(\sr_reg[1]_37 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[0]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [0]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [0]),
        .O(\sr_reg[1]_53 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[10]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [10]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [10]),
        .O(\sr_reg[1]_26 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[10]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [10]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [10]),
        .O(\sr_reg[0]_48 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[10]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [10]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [10]),
        .O(\sr_reg[1]_47 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[10]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [10]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [10]),
        .O(\sr_reg[1]_63 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[11]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [11]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [11]),
        .O(\sr_reg[1]_25 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[11]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [11]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [11]),
        .O(\sr_reg[0]_49 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[11]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [11]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [11]),
        .O(\sr_reg[1]_48 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[11]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [11]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [11]),
        .O(\sr_reg[1]_64 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[12]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [12]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [12]),
        .O(\sr_reg[1]_24 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[12]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [12]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [12]),
        .O(\sr_reg[0]_50 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[12]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [12]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [12]),
        .O(\sr_reg[1]_49 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[12]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [12]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [12]),
        .O(\sr_reg[1]_65 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[13]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [13]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [13]),
        .O(\sr_reg[1]_23 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[13]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [13]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [13]),
        .O(\sr_reg[0]_51 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[13]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [13]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [13]),
        .O(\sr_reg[1]_50 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[13]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [13]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [13]),
        .O(\sr_reg[1]_66 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[14]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [14]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [14]),
        .O(\sr_reg[1]_22 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[14]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [14]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [14]),
        .O(\sr_reg[0]_52 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[14]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [14]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [14]),
        .O(\sr_reg[1]_51 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[14]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [14]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [14]),
        .O(\sr_reg[1]_67 ));
  LUT4 #(
    .INIT(16'h6F60)) 
    \badr[15]_INST_0_i_145 
       (.I0(sr[5]),
        .I1(sr[7]),
        .I2(\rgf_selc1_wb[1]_i_16 [3]),
        .I3(sr[4]),
        .O(\sr_reg[5]_1 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[15]_INST_0_i_16 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [15]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [15]),
        .O(\sr_reg[1]_21 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_185 
       (.I0(sr[0]),
        .I1(sr[1]),
        .O(\sr_reg[0]_37 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[15]_INST_0_i_20 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [15]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [15]),
        .O(\sr_reg[0]_53 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA0305F30)) 
    \badr[15]_INST_0_i_295 
       (.I0(sr[7]),
        .I1(sr[4]),
        .I2(\badr[15]_INST_0_i_208 [1]),
        .I3(\badr[15]_INST_0_i_208 [3]),
        .I4(sr[5]),
        .I5(\badr[15]_INST_0_i_208 [4]),
        .O(\sr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[15]_INST_0_i_31 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [15]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [15]),
        .O(\sr_reg[1]_52 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[15]_INST_0_i_34 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [15]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [15]),
        .O(\sr_reg[1]_68 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[1]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [1]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [1]),
        .O(\sr_reg[1]_35 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[1]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [1]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [1]),
        .O(\sr_reg[0]_39 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[1]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [1]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [1]),
        .O(\sr_reg[1]_38 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[1]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [1]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [1]),
        .O(\sr_reg[1]_54 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[2]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [2]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [2]),
        .O(\sr_reg[1]_34 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[2]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [2]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [2]),
        .O(\sr_reg[0]_40 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[2]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [2]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [2]),
        .O(\sr_reg[1]_39 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[2]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [2]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [2]),
        .O(\sr_reg[1]_55 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[3]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [3]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [3]),
        .O(\sr_reg[1]_33 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[3]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [3]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [3]),
        .O(\sr_reg[0]_41 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[3]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [3]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [3]),
        .O(\sr_reg[1]_40 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[3]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [3]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [3]),
        .O(\sr_reg[1]_56 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[4]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [4]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [4]),
        .O(\sr_reg[1]_32 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[4]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [4]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [4]),
        .O(\sr_reg[0]_42 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[4]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [4]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [4]),
        .O(\sr_reg[1]_41 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[4]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [4]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [4]),
        .O(\sr_reg[1]_57 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[5]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [5]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [5]),
        .O(\sr_reg[1]_31 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[5]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [5]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [5]),
        .O(\sr_reg[0]_43 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[5]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [5]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [5]),
        .O(\sr_reg[1]_42 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[5]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [5]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [5]),
        .O(\sr_reg[1]_58 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[6]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [6]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [6]),
        .O(\sr_reg[1]_30 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[6]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [6]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [6]),
        .O(\sr_reg[0]_44 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[6]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [6]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [6]),
        .O(\sr_reg[1]_43 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[6]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [6]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [6]),
        .O(\sr_reg[1]_59 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[7]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [7]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [7]),
        .O(\sr_reg[1]_29 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[7]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [7]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [7]),
        .O(\sr_reg[0]_45 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[7]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [7]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [7]),
        .O(\sr_reg[1]_44 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[7]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [7]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [7]),
        .O(\sr_reg[1]_60 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[8]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [8]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [8]),
        .O(\sr_reg[1]_28 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[8]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [8]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [8]),
        .O(\sr_reg[0]_46 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[8]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [8]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [8]),
        .O(\sr_reg[1]_45 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[8]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [8]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [8]),
        .O(\sr_reg[1]_61 ));
  LUT6 #(
    .INIT(64'h1110101011000000)) 
    \badr[9]_INST_0_i_14 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(a1bus_sel_0[1]),
        .I4(\rgf_c1bus_wb[4]_i_47 [9]),
        .I5(\rgf_c1bus_wb[4]_i_47_0 [9]),
        .O(\sr_reg[1]_27 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[9]_INST_0_i_16 
       (.I0(sr[0]),
        .I1(sr[1]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_39_0 [9]),
        .I4(gr6_bus1),
        .I5(\rgf_c1bus_wb[4]_i_39 [9]),
        .O(\sr_reg[0]_47 ));
  LUT6 #(
    .INIT(64'hFF404040FF000000)) 
    \badr[9]_INST_0_i_20 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\rgf_c1bus_wb[4]_i_45_0 [9]),
        .I4(gr6_bus1_0),
        .I5(\rgf_c1bus_wb[4]_i_45 [9]),
        .O(\sr_reg[1]_46 ));
  LUT6 #(
    .INIT(64'hFF808080FF000000)) 
    \badr[9]_INST_0_i_23 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(a1bus_sel_0[0]),
        .I3(\badr[15]_INST_0_i_7_0 [9]),
        .I4(gr6_bus1_1),
        .I5(\badr[15]_INST_0_i_7 [9]),
        .O(\sr_reg[1]_62 ));
  LUT4 #(
    .INIT(16'h0200)) 
    \bbus_o[0]_INST_0_i_11 
       (.I0(b0bus_sel_0),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\i_/bbus_o[4]_INST_0_i_5 [0]),
        .O(\sr_reg[0]_4 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bbus_o[0]_INST_0_i_15 
       (.I0(b0bus_sel_0),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\i_/bbus_o[4]_INST_0_i_6 [0]),
        .O(\sr_reg[1]_4 ));
  LUT4 #(
    .INIT(16'h0200)) 
    \bbus_o[1]_INST_0_i_10 
       (.I0(b0bus_sel_0),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\i_/bbus_o[4]_INST_0_i_5 [1]),
        .O(\sr_reg[0]_3 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bbus_o[1]_INST_0_i_14 
       (.I0(b0bus_sel_0),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\i_/bbus_o[4]_INST_0_i_6 [1]),
        .O(\sr_reg[1]_3 ));
  LUT4 #(
    .INIT(16'h0200)) 
    \bbus_o[2]_INST_0_i_11 
       (.I0(b0bus_sel_0),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\i_/bbus_o[4]_INST_0_i_5 [2]),
        .O(\sr_reg[0]_2 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bbus_o[2]_INST_0_i_15 
       (.I0(b0bus_sel_0),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\i_/bbus_o[4]_INST_0_i_6 [2]),
        .O(\sr_reg[1]_2 ));
  LUT4 #(
    .INIT(16'h0200)) 
    \bbus_o[3]_INST_0_i_11 
       (.I0(b0bus_sel_0),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\i_/bbus_o[4]_INST_0_i_5 [3]),
        .O(\sr_reg[0]_1 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bbus_o[3]_INST_0_i_15 
       (.I0(b0bus_sel_0),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\i_/bbus_o[4]_INST_0_i_6 [3]),
        .O(\sr_reg[1]_1 ));
  LUT4 #(
    .INIT(16'h0200)) 
    \bbus_o[4]_INST_0_i_12 
       (.I0(b0bus_sel_0),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\i_/bbus_o[4]_INST_0_i_5 [4]),
        .O(\sr_reg[0]_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bbus_o[4]_INST_0_i_17 
       (.I0(b0bus_sel_0),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\i_/bbus_o[4]_INST_0_i_6 [4]),
        .O(\sr_reg[1]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_81 
       (.I0(sr[1]),
        .I1(sr[0]),
        .O(\sr_reg[1]_20 ));
  LUT4 #(
    .INIT(16'h6F60)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(sr[5]),
        .I1(sr[7]),
        .I2(\badr[15]_INST_0_i_208 [3]),
        .I3(sr[4]),
        .O(\sr_reg[5]_2 ));
  LUT5 #(
    .INIT(32'h10000010)) 
    ctl_fetch0_fl_i_10
       (.I0(\badr[15]_INST_0_i_208 [3]),
        .I1(\badr[15]_INST_0_i_208 [2]),
        .I2(sr[4]),
        .I3(sr[5]),
        .I4(sr[7]),
        .O(\sr_reg[4]_1 ));
  LUT5 #(
    .INIT(32'h8A8A088A)) 
    ctl_fetch0_fl_i_42
       (.I0(irq),
        .I1(irq_lev[1]),
        .I2(sr[3]),
        .I3(sr[2]),
        .I4(irq_lev[0]),
        .O(irq_0));
  LUT6 #(
    .INIT(64'h0303999F00000000)) 
    ctl_fetch0_fl_i_7
       (.I0(sr[5]),
        .I1(sr[7]),
        .I2(\badr[15]_INST_0_i_208 [3]),
        .I3(sr[4]),
        .I4(\badr[15]_INST_0_i_208 [2]),
        .I5(\badr[15]_INST_0_i_208 [1]),
        .O(\sr_reg[5]_6 ));
  LUT3 #(
    .INIT(8'h37)) 
    ctl_fetch1_fl_i_23
       (.I0(sr[10]),
        .I1(Q),
        .I2(ctl_fetch1_fl_i_15),
        .O(\sr_reg[10]_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch1_fl_i_26
       (.I0(sr[5]),
        .I1(sr[7]),
        .O(\sr_reg[5]_3 ));
  LUT6 #(
    .INIT(64'h8B88BBBB8B888B88)) 
    ctl_fetch1_fl_i_33
       (.I0(ctl_fetch1_fl_i_38_n_0),
        .I1(\rgf_selc1_wb[1]_i_16 [1]),
        .I2(sr[6]),
        .I3(\rgf_selc1_wb[1]_i_16 [2]),
        .I4(sr[5]),
        .I5(\rgf_selc1_wb[1]_i_16 [3]),
        .O(\sr_reg[6]_5 ));
  LUT5 #(
    .INIT(32'h41634177)) 
    ctl_fetch1_fl_i_38
       (.I0(\rgf_selc1_wb[1]_i_16 [2]),
        .I1(sr[7]),
        .I2(sr[5]),
        .I3(\rgf_selc1_wb[1]_i_16 [3]),
        .I4(sr[4]),
        .O(ctl_fetch1_fl_i_38_n_0));
  LUT5 #(
    .INIT(32'h2020A220)) 
    fch_irq_req_fl_i_1
       (.I0(irq),
        .I1(irq_lev[1]),
        .I2(sr[3]),
        .I3(sr[2]),
        .I4(irq_lev[0]),
        .O(fch_irq_req));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[0]_i_13 
       (.I0(sr[6]),
        .I1(\rgf_c0bus_wb[0]_i_5 ),
        .O(\sr_reg[6]_4 ));
  LUT5 #(
    .INIT(32'h44444447)) 
    \rgf_c0bus_wb[13]_i_33 
       (.I0(sr[6]),
        .I1(\sr[4]_i_188 ),
        .I2(\sr[4]_i_188_0 ),
        .I3(\sr[4]_i_188_1 ),
        .I4(\sr[4]_i_188_2 ),
        .O(\sr_reg[6]_2 ));
  LUT5 #(
    .INIT(32'h44444447)) 
    \rgf_c0bus_wb[4]_i_28 
       (.I0(sr[6]),
        .I1(\sr[4]_i_188 ),
        .I2(\rgf_c0bus_wb[4]_i_10 ),
        .I3(\rgf_c0bus_wb[4]_i_10_0 ),
        .I4(\rgf_c0bus_wb[4]_i_10_1 ),
        .O(\sr_reg[6]_3 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_136 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [4]),
        .O(\sr_reg[0]_32 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_138 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [4]),
        .O(\sr_reg[0]_16 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_140 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [3]),
        .O(\sr_reg[1]_16 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_142 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [3]),
        .O(\sr_reg[0]_33 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_144 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [3]),
        .O(\sr_reg[0]_17 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_146 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [2]),
        .O(\sr_reg[0]_34 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_148 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [2]),
        .O(\sr_reg[0]_18 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_150 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [1]),
        .O(\sr_reg[1]_18 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_152 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [1]),
        .O(\sr_reg[0]_35 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_154 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [1]),
        .O(\sr_reg[0]_19 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_156 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [15]),
        .O(\sr_reg[0]_21 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_158 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [15]),
        .O(\sr_reg[0]_5 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_160 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [14]),
        .O(\sr_reg[1]_6 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_162 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [14]),
        .O(\sr_reg[0]_22 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_164 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [14]),
        .O(\sr_reg[0]_6 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_166 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [0]),
        .O(\sr_reg[0]_20 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_168 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [15]),
        .O(\sr_reg[1]_5 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_170 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [12]),
        .O(\sr_reg[0]_24 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_172 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [12]),
        .O(\sr_reg[0]_8 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_174 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [13]),
        .O(\sr_reg[0]_23 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_176 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [13]),
        .O(\sr_reg[0]_7 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_178 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [13]),
        .O(\sr_reg[1]_7 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_180 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [5]),
        .O(\sr_reg[0]_31 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_182 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [5]),
        .O(\sr_reg[0]_15 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_184 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [5]),
        .O(\sr_reg[1]_14 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_186 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [6]),
        .O(\sr_reg[0]_30 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_188 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [6]),
        .O(\sr_reg[0]_14 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_190 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [7]),
        .O(\sr_reg[0]_29 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_192 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [7]),
        .O(\sr_reg[0]_13 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_194 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [7]),
        .O(\sr_reg[1]_12 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_196 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [8]),
        .O(\sr_reg[0]_28 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_198 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [8]),
        .O(\sr_reg[0]_12 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_200 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [9]),
        .O(\sr_reg[0]_27 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_202 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [9]),
        .O(\sr_reg[0]_11 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_204 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [9]),
        .O(\sr_reg[1]_11 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_206 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [10]),
        .O(\sr_reg[0]_26 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_208 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [10]),
        .O(\sr_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h111111111111111D)) 
    \rgf_c1bus_wb[4]_i_21 
       (.I0(sr[6]),
        .I1(\sr[4]_i_160 ),
        .I2(\sr[4]_i_172 ),
        .I3(\sr[4]_i_172_0 ),
        .I4(\sr[4]_i_172_1 ),
        .I5(\sr[4]_i_172_2 ),
        .O(\sr_reg[6]_1 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_210 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [11]),
        .O(\sr_reg[0]_25 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[4]_i_212 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\badr[15]_INST_0_i_7 [11]),
        .O(\sr_reg[0]_9 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_214 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [11]),
        .O(\sr_reg[1]_9 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[4]_i_216 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [2]),
        .O(\sr_reg[1]_17 ));
  LUT6 #(
    .INIT(64'h6F60909FFFFFFFFF)) 
    \rgf_selc0_wb[1]_i_25 
       (.I0(sr[5]),
        .I1(sr[7]),
        .I2(\badr[15]_INST_0_i_208 [3]),
        .I3(sr[4]),
        .I4(\badr[15]_INST_0_i_208 [0]),
        .I5(\badr[15]_INST_0_i_208 [1]),
        .O(\sr_reg[5]_5 ));
  LUT6 #(
    .INIT(64'h6F60909FFFFFFFFF)) 
    \rgf_selc1_wb[1]_i_25 
       (.I0(sr[5]),
        .I1(sr[7]),
        .I2(\rgf_selc1_wb[1]_i_16 [3]),
        .I3(sr[4]),
        .I4(\rgf_selc1_wb[1]_i_16 [0]),
        .I5(\rgf_selc1_wb[1]_i_16 [1]),
        .O(\sr_reg[5]_4 ));
  LUT6 #(
    .INIT(64'h111111111111111D)) 
    \sr[4]_i_212 
       (.I0(sr[6]),
        .I1(\sr[4]_i_160 ),
        .I2(\sr[4]_i_160_0 ),
        .I3(\sr[4]_i_160_1 ),
        .I4(\sr[4]_i_160_2 ),
        .I5(\sr[4]_i_160_3 ),
        .O(\sr_reg[6]_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \sr[4]_i_259 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [12]),
        .O(\sr_reg[1]_8 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \sr[4]_i_261 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [10]),
        .O(\sr_reg[1]_10 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \sr[4]_i_263 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[0]),
        .I2(sr[1]),
        .I3(\rgf_c1bus_wb[4]_i_45 [0]),
        .O(\sr_reg[0]_36 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \sr[4]_i_265 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [0]),
        .O(\sr_reg[1]_19 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \sr[4]_i_267 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [4]),
        .O(\sr_reg[1]_15 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \sr[4]_i_269 
       (.I0(a1bus_sel_0[0]),
        .I1(sr[1]),
        .I2(sr[0]),
        .I3(\rgf_c1bus_wb[4]_i_39 [6]),
        .O(\sr_reg[1]_13 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_5 
       (.I0(sr[4]),
        .I1(\sr_reg[5]_7 ),
        .O(\sr_reg[4]_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[5]_i_5 
       (.I0(sr[5]),
        .I1(\sr_reg[5]_7 ),
        .O(\sr_reg[5]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [0]),
        .Q(sr[0]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [10]),
        .Q(sr[10]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [11]),
        .Q(sr[11]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [12]),
        .Q(sr[12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [13]),
        .Q(sr[13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [14]),
        .Q(sr[14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [15]),
        .Q(sr[15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [1]),
        .Q(sr[1]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [2]),
        .Q(sr[2]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [3]),
        .Q(sr[3]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [4]),
        .Q(sr[4]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [5]),
        .Q(sr[5]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [6]),
        .Q(sr[6]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [7]),
        .Q(sr[7]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [8]),
        .Q(sr[8]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[15]_1 [9]),
        .Q(sr[9]),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h3C333CCCEEFFEEFF)) 
    \stat[2]_i_17 
       (.I0(sr[4]),
        .I1(\rgf_selc1_wb[1]_i_16 [0]),
        .I2(sr[7]),
        .I3(\rgf_selc1_wb[1]_i_16 [1]),
        .I4(sr[6]),
        .I5(\rgf_selc1_wb[1]_i_16 [2]),
        .O(\sr_reg[4]_2 ));
  LUT6 #(
    .INIT(64'h37F7FB3B37F7CB0B)) 
    \stat[2]_i_7 
       (.I0(sr[6]),
        .I1(\badr[15]_INST_0_i_208 [2]),
        .I2(\badr[15]_INST_0_i_208 [1]),
        .I3(sr[7]),
        .I4(\badr[15]_INST_0_i_208 [0]),
        .I5(sr[4]),
        .O(\sr_reg[6]_6 ));
endmodule

module mcss_rgf_treg
   (.out({tr[15],tr[14],tr[13],tr[12],tr[11],tr[10],tr[9],tr[8],tr[7],tr[6],tr[5],tr[4],tr[3],tr[2],tr[1],tr[0]}),
    \sr_reg[6] ,
    \sr_reg[6]_0 ,
    badrx,
    \rgf_c1bus_wb[4]_i_13 ,
    \rgf_c1bus_wb[4]_i_13_0 ,
    \rgf_c1bus_wb[4]_i_13_1 ,
    \rgf_c1bus_wb[4]_i_13_2 ,
    \rgf_c1bus_wb[4]_i_13_3 ,
    \rgf_c1bus_wb[4]_i_13_4 ,
    \sr[4]_i_167 ,
    \sr[4]_i_167_0 ,
    \sr[4]_i_167_1 ,
    \sr[4]_i_167_2 ,
    .badrx_15_sp_1(badrx_15_sn_1),
    SR,
    \tr_reg[15]_0 ,
    clk);
  output \sr_reg[6] ;
  output \sr_reg[6]_0 ;
  output [15:0]badrx;
  input \rgf_c1bus_wb[4]_i_13 ;
  input [0:0]\rgf_c1bus_wb[4]_i_13_0 ;
  input \rgf_c1bus_wb[4]_i_13_1 ;
  input \rgf_c1bus_wb[4]_i_13_2 ;
  input \rgf_c1bus_wb[4]_i_13_3 ;
  input [0:0]\rgf_c1bus_wb[4]_i_13_4 ;
  input \sr[4]_i_167 ;
  input [0:0]\sr[4]_i_167_0 ;
  input \sr[4]_i_167_1 ;
  input \sr[4]_i_167_2 ;
  input [0:0]SR;
  input [15:0]\tr_reg[15]_0 ;
  input clk;
     output [15:0]tr;
  input badrx_15_sn_1;

  wire \<const1> ;
  wire [0:0]SR;
  wire [15:0]badrx;
  wire badrx_15_sn_1;
  wire clk;
  wire \rgf_c1bus_wb[4]_i_13 ;
  wire [0:0]\rgf_c1bus_wb[4]_i_13_0 ;
  wire \rgf_c1bus_wb[4]_i_13_1 ;
  wire \rgf_c1bus_wb[4]_i_13_2 ;
  wire \rgf_c1bus_wb[4]_i_13_3 ;
  wire [0:0]\rgf_c1bus_wb[4]_i_13_4 ;
  wire \sr[4]_i_167 ;
  wire [0:0]\sr[4]_i_167_0 ;
  wire \sr[4]_i_167_1 ;
  wire \sr[4]_i_167_2 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  (* DONT_TOUCH *) wire [15:0]tr;
  wire [15:0]\tr_reg[15]_0 ;

  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[0]_INST_0 
       (.I0(tr[0]),
        .I1(badrx_15_sn_1),
        .O(badrx[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[10]_INST_0 
       (.I0(tr[10]),
        .I1(badrx_15_sn_1),
        .O(badrx[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[11]_INST_0 
       (.I0(tr[11]),
        .I1(badrx_15_sn_1),
        .O(badrx[11]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[12]_INST_0 
       (.I0(tr[12]),
        .I1(badrx_15_sn_1),
        .O(badrx[12]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[13]_INST_0 
       (.I0(tr[13]),
        .I1(badrx_15_sn_1),
        .O(badrx[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[14]_INST_0 
       (.I0(tr[14]),
        .I1(badrx_15_sn_1),
        .O(badrx[14]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[15]_INST_0 
       (.I0(tr[15]),
        .I1(badrx_15_sn_1),
        .O(badrx[15]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[1]_INST_0 
       (.I0(tr[1]),
        .I1(badrx_15_sn_1),
        .O(badrx[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[2]_INST_0 
       (.I0(tr[2]),
        .I1(badrx_15_sn_1),
        .O(badrx[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[3]_INST_0 
       (.I0(tr[3]),
        .I1(badrx_15_sn_1),
        .O(badrx[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[4]_INST_0 
       (.I0(tr[4]),
        .I1(badrx_15_sn_1),
        .O(badrx[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[5]_INST_0 
       (.I0(tr[5]),
        .I1(badrx_15_sn_1),
        .O(badrx[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[6]_INST_0 
       (.I0(tr[6]),
        .I1(badrx_15_sn_1),
        .O(badrx[6]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[7]_INST_0 
       (.I0(tr[7]),
        .I1(badrx_15_sn_1),
        .O(badrx[7]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[8]_INST_0 
       (.I0(tr[8]),
        .I1(badrx_15_sn_1),
        .O(badrx[8]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[9]_INST_0 
       (.I0(tr[9]),
        .I1(badrx_15_sn_1),
        .O(badrx[9]));
  LUT6 #(
    .INIT(64'h00000001FFFF0001)) 
    \rgf_c1bus_wb[4]_i_30 
       (.I0(\rgf_c1bus_wb[4]_i_13 ),
        .I1(\rgf_c1bus_wb[4]_i_13_0 ),
        .I2(\rgf_c1bus_wb[4]_i_13_1 ),
        .I3(\rgf_c1bus_wb[4]_i_13_2 ),
        .I4(\rgf_c1bus_wb[4]_i_13_3 ),
        .I5(\rgf_c1bus_wb[4]_i_13_4 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'h00000001FFFF0001)) 
    \sr[4]_i_214 
       (.I0(\sr[4]_i_167 ),
        .I1(\sr[4]_i_167_0 ),
        .I2(\sr[4]_i_167_1 ),
        .I3(\sr[4]_i_167_2 ),
        .I4(\rgf_c1bus_wb[4]_i_13_3 ),
        .I5(\rgf_c1bus_wb[4]_i_13_4 ),
        .O(\sr_reg[6]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [0]),
        .Q(tr[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [10]),
        .Q(tr[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [11]),
        .Q(tr[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [12]),
        .Q(tr[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [13]),
        .Q(tr[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [14]),
        .Q(tr[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [15]),
        .Q(tr[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [1]),
        .Q(tr[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [2]),
        .Q(tr[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [3]),
        .Q(tr[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [4]),
        .Q(tr[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [5]),
        .Q(tr[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [6]),
        .Q(tr[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [7]),
        .Q(tr[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [8]),
        .Q(tr[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\tr_reg[15]_0 [9]),
        .Q(tr[9]),
        .R(SR));
endmodule

(* STRUCTURAL_NETLIST = "yes" *)
module moscoviumss
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdatx,
    fdat,
    bdatr,
    fadr,
    bcmd,
    badrx,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o);
//
//	Moscovium-SS 16 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2024/08/31	ver.1.10
//		instruction: hdown
//
//	2023/10/28	ver.1.08
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.06
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.04
//		instruction: divlqr, divlrr, divur, divsr, mulur, mulsr
//
//	2022/10/22	ver.1.02
//		corresponding to interrupt vector / level
//
//	2022/06/11	ver.1.00
//		Moscovium-SS: Super Scalar Edition
//
// ================================
//
//	2022/06/04	ver.1.12
//		instruction: csft, csfti
//		revised register file block
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core cpu edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [15:0]fdatx;
  input [15:0]fdat;
  input [15:0]bdatr;
  output [15:0]fadr;
  output [2:0]bcmd;
  output [15:0]badrx;
  output [15:0]badr;
  output [15:0]bdatw;
  input crdy;
  input [15:0]cbus_i;
  output [4:0]ccmd;
  output [15:0]abus_o;
  output [15:0]bbus_o;

  wire [15:0]a0bus_0;
  wire [7:0]a0bus_sel_0;
  wire [5:0]a0bus_sel_cr;
  wire [15:0]a1bus_0;
  wire [15:15]a1bus_b02;
  wire [7:4]a1bus_sel_0;
  wire [5:1]a1bus_sel_cr;
  wire [15:0]a1bus_sr;
  wire [15:0]abus_o;
  wire alu0_n_0;
  wire alu0_n_1;
  wire alu0_n_10;
  wire alu0_n_11;
  wire alu0_n_13;
  wire alu0_n_14;
  wire alu0_n_15;
  wire alu0_n_17;
  wire alu0_n_2;
  wire alu0_n_3;
  wire alu0_n_4;
  wire alu0_n_5;
  wire alu0_n_6;
  wire alu0_n_7;
  wire alu0_n_8;
  wire alu0_n_9;
  wire alu1_n_0;
  wire alu1_n_1;
  wire alu1_n_10;
  wire alu1_n_11;
  wire alu1_n_13;
  wire alu1_n_14;
  wire alu1_n_15;
  wire alu1_n_17;
  wire alu1_n_2;
  wire alu1_n_3;
  wire alu1_n_4;
  wire alu1_n_5;
  wire alu1_n_6;
  wire alu1_n_7;
  wire alu1_n_8;
  wire alu1_n_9;
  wire [18:18]\art/add/tout ;
  wire [18:18]\art/add/tout_0 ;
  wire [15:15]\art/p_0_in ;
  wire [15:15]\art/p_0_in_1 ;
  wire [2:1]b0bus_sel_0;
  wire [5:1]b0bus_sel_cr;
  wire [15:0]b0bus_sr;
  wire [4:0]b1bus_b02;
  wire [5:0]b1bus_sel_cr;
  wire [14:0]b1bus_sr;
  wire [15:0]badr;
  wire [15:0]badrx;
  wire [0:0]\bank02/p_0_in ;
  wire [4:0]\bank02/p_0_in2_in ;
  wire [0:0]\bank02/p_1_in ;
  wire [4:0]\bank02/p_1_in3_in ;
  wire [3:3]bank_sel;
  wire [15:0]bbus_o;
  wire [2:0]bcmd;
  wire [5:4]\bctl/ctl/p_0_in ;
  wire [0:0]\bctl/ctl/stat_nx ;
  wire [15:0]bdatr;
  wire [15:0]bdatw;
  wire brdy;
  wire [15:0]c0bus;
  wire [15:0]c1bus;
  wire [15:0]cbus_i;
  wire [4:0]ccmd;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl0_n_0;
  wire ctl0_n_1;
  wire ctl0_n_10;
  wire ctl0_n_11;
  wire ctl0_n_12;
  wire ctl0_n_13;
  wire ctl0_n_14;
  wire ctl0_n_15;
  wire ctl0_n_16;
  wire ctl0_n_17;
  wire ctl0_n_18;
  wire ctl0_n_19;
  wire ctl0_n_20;
  wire ctl0_n_21;
  wire ctl0_n_22;
  wire ctl0_n_23;
  wire ctl0_n_24;
  wire ctl0_n_25;
  wire ctl0_n_26;
  wire ctl0_n_27;
  wire ctl0_n_28;
  wire ctl0_n_5;
  wire ctl0_n_6;
  wire ctl0_n_7;
  wire ctl0_n_8;
  wire ctl0_n_9;
  wire ctl1_n_0;
  wire ctl1_n_1;
  wire ctl1_n_10;
  wire ctl1_n_11;
  wire ctl1_n_12;
  wire ctl1_n_13;
  wire ctl1_n_14;
  wire ctl1_n_15;
  wire ctl1_n_16;
  wire ctl1_n_17;
  wire ctl1_n_18;
  wire ctl1_n_19;
  wire ctl1_n_20;
  wire ctl1_n_21;
  wire ctl1_n_22;
  wire ctl1_n_5;
  wire ctl1_n_6;
  wire ctl1_n_7;
  wire ctl1_n_8;
  wire ctl1_n_9;
  wire ctl_bcc_take0_fl;
  wire ctl_bcc_take1_fl;
  wire [0:0]ctl_sela0;
  wire [2:0]ctl_sela0_rn;
  wire [0:0]ctl_selb0_0;
  wire [1:0]ctl_selb0_rn;
  wire [1:1]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [1:1]ctl_selc0;
  wire [2:0]ctl_selc0_rn;
  wire [1:1]ctl_selc1;
  wire [0:0]ctl_selc1_rn;
  wire [15:0]fadr;
  wire [15:0]fch_ir0;
  wire [15:0]fch_ir1;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire fch_memacc1;
  wire fch_n_1000;
  wire fch_n_1001;
  wire fch_n_1002;
  wire fch_n_1003;
  wire fch_n_1004;
  wire fch_n_1005;
  wire fch_n_1006;
  wire fch_n_1007;
  wire fch_n_1008;
  wire fch_n_1009;
  wire fch_n_1010;
  wire fch_n_1011;
  wire fch_n_1012;
  wire fch_n_1013;
  wire fch_n_1014;
  wire fch_n_1015;
  wire fch_n_1016;
  wire fch_n_1017;
  wire fch_n_1018;
  wire fch_n_1019;
  wire fch_n_1020;
  wire fch_n_1021;
  wire fch_n_1022;
  wire fch_n_1023;
  wire fch_n_1024;
  wire fch_n_1025;
  wire fch_n_1026;
  wire fch_n_1027;
  wire fch_n_1028;
  wire fch_n_1029;
  wire fch_n_1030;
  wire fch_n_1031;
  wire fch_n_1032;
  wire fch_n_1033;
  wire fch_n_1034;
  wire fch_n_1035;
  wire fch_n_1036;
  wire fch_n_1037;
  wire fch_n_1038;
  wire fch_n_1039;
  wire fch_n_1040;
  wire fch_n_1041;
  wire fch_n_1042;
  wire fch_n_1043;
  wire fch_n_1044;
  wire fch_n_1045;
  wire fch_n_1046;
  wire fch_n_1047;
  wire fch_n_1048;
  wire fch_n_1049;
  wire fch_n_105;
  wire fch_n_1050;
  wire fch_n_1051;
  wire fch_n_1052;
  wire fch_n_1053;
  wire fch_n_1054;
  wire fch_n_1055;
  wire fch_n_1056;
  wire fch_n_1057;
  wire fch_n_1058;
  wire fch_n_1059;
  wire fch_n_106;
  wire fch_n_1060;
  wire fch_n_1061;
  wire fch_n_1062;
  wire fch_n_1063;
  wire fch_n_1064;
  wire fch_n_1065;
  wire fch_n_1066;
  wire fch_n_1067;
  wire fch_n_1068;
  wire fch_n_1069;
  wire fch_n_107;
  wire fch_n_1070;
  wire fch_n_1071;
  wire fch_n_1072;
  wire fch_n_1073;
  wire fch_n_1074;
  wire fch_n_1075;
  wire fch_n_1076;
  wire fch_n_1077;
  wire fch_n_1078;
  wire fch_n_1079;
  wire fch_n_108;
  wire fch_n_1080;
  wire fch_n_1081;
  wire fch_n_1082;
  wire fch_n_1083;
  wire fch_n_1084;
  wire fch_n_1085;
  wire fch_n_1086;
  wire fch_n_1087;
  wire fch_n_1088;
  wire fch_n_1089;
  wire fch_n_1090;
  wire fch_n_1091;
  wire fch_n_1092;
  wire fch_n_1093;
  wire fch_n_1094;
  wire fch_n_1095;
  wire fch_n_1096;
  wire fch_n_1097;
  wire fch_n_1098;
  wire fch_n_1099;
  wire fch_n_1100;
  wire fch_n_1101;
  wire fch_n_1102;
  wire fch_n_1103;
  wire fch_n_1104;
  wire fch_n_1105;
  wire fch_n_1106;
  wire fch_n_1107;
  wire fch_n_1108;
  wire fch_n_1109;
  wire fch_n_1110;
  wire fch_n_1111;
  wire fch_n_1112;
  wire fch_n_1113;
  wire fch_n_1114;
  wire fch_n_1115;
  wire fch_n_1116;
  wire fch_n_1117;
  wire fch_n_1118;
  wire fch_n_1119;
  wire fch_n_1120;
  wire fch_n_1121;
  wire fch_n_1122;
  wire fch_n_1123;
  wire fch_n_1124;
  wire fch_n_1125;
  wire fch_n_1126;
  wire fch_n_1127;
  wire fch_n_1128;
  wire fch_n_1129;
  wire fch_n_1130;
  wire fch_n_1131;
  wire fch_n_1132;
  wire fch_n_1133;
  wire fch_n_1134;
  wire fch_n_1135;
  wire fch_n_1136;
  wire fch_n_1137;
  wire fch_n_1138;
  wire fch_n_1139;
  wire fch_n_1140;
  wire fch_n_1141;
  wire fch_n_1142;
  wire fch_n_1143;
  wire fch_n_1144;
  wire fch_n_1145;
  wire fch_n_1146;
  wire fch_n_1147;
  wire fch_n_1148;
  wire fch_n_1149;
  wire fch_n_1150;
  wire fch_n_1151;
  wire fch_n_1152;
  wire fch_n_1153;
  wire fch_n_1154;
  wire fch_n_1155;
  wire fch_n_1156;
  wire fch_n_1157;
  wire fch_n_1158;
  wire fch_n_1159;
  wire fch_n_1160;
  wire fch_n_1161;
  wire fch_n_1162;
  wire fch_n_1163;
  wire fch_n_1164;
  wire fch_n_1165;
  wire fch_n_1166;
  wire fch_n_1167;
  wire fch_n_1168;
  wire fch_n_1169;
  wire fch_n_1170;
  wire fch_n_1171;
  wire fch_n_1172;
  wire fch_n_1173;
  wire fch_n_1174;
  wire fch_n_1175;
  wire fch_n_1176;
  wire fch_n_1177;
  wire fch_n_1178;
  wire fch_n_1179;
  wire fch_n_1180;
  wire fch_n_1181;
  wire fch_n_1182;
  wire fch_n_1183;
  wire fch_n_1184;
  wire fch_n_1185;
  wire fch_n_1186;
  wire fch_n_1187;
  wire fch_n_1188;
  wire fch_n_1189;
  wire fch_n_1190;
  wire fch_n_1191;
  wire fch_n_1192;
  wire fch_n_1193;
  wire fch_n_1194;
  wire fch_n_1195;
  wire fch_n_1196;
  wire fch_n_1197;
  wire fch_n_1198;
  wire fch_n_1199;
  wire fch_n_1200;
  wire fch_n_1201;
  wire fch_n_1202;
  wire fch_n_146;
  wire fch_n_147;
  wire fch_n_148;
  wire fch_n_149;
  wire fch_n_150;
  wire fch_n_151;
  wire fch_n_152;
  wire fch_n_153;
  wire fch_n_154;
  wire fch_n_155;
  wire fch_n_156;
  wire fch_n_157;
  wire fch_n_158;
  wire fch_n_159;
  wire fch_n_160;
  wire fch_n_161;
  wire fch_n_162;
  wire fch_n_163;
  wire fch_n_164;
  wire fch_n_165;
  wire fch_n_166;
  wire fch_n_167;
  wire fch_n_168;
  wire fch_n_169;
  wire fch_n_184;
  wire fch_n_185;
  wire fch_n_186;
  wire fch_n_187;
  wire fch_n_189;
  wire fch_n_190;
  wire fch_n_191;
  wire fch_n_192;
  wire fch_n_193;
  wire fch_n_194;
  wire fch_n_195;
  wire fch_n_196;
  wire fch_n_197;
  wire fch_n_198;
  wire fch_n_199;
  wire fch_n_200;
  wire fch_n_201;
  wire fch_n_202;
  wire fch_n_203;
  wire fch_n_204;
  wire fch_n_205;
  wire fch_n_221;
  wire fch_n_222;
  wire fch_n_223;
  wire fch_n_224;
  wire fch_n_225;
  wire fch_n_226;
  wire fch_n_227;
  wire fch_n_228;
  wire fch_n_229;
  wire fch_n_230;
  wire fch_n_231;
  wire fch_n_232;
  wire fch_n_233;
  wire fch_n_234;
  wire fch_n_235;
  wire fch_n_236;
  wire fch_n_242;
  wire fch_n_248;
  wire fch_n_249;
  wire fch_n_250;
  wire fch_n_251;
  wire fch_n_253;
  wire fch_n_254;
  wire fch_n_255;
  wire fch_n_256;
  wire fch_n_257;
  wire fch_n_258;
  wire fch_n_264;
  wire fch_n_265;
  wire fch_n_267;
  wire fch_n_268;
  wire fch_n_269;
  wire fch_n_270;
  wire fch_n_271;
  wire fch_n_272;
  wire fch_n_273;
  wire fch_n_274;
  wire fch_n_275;
  wire fch_n_276;
  wire fch_n_277;
  wire fch_n_278;
  wire fch_n_279;
  wire fch_n_280;
  wire fch_n_281;
  wire fch_n_282;
  wire fch_n_283;
  wire fch_n_284;
  wire fch_n_289;
  wire fch_n_293;
  wire fch_n_294;
  wire fch_n_295;
  wire fch_n_298;
  wire fch_n_299;
  wire fch_n_300;
  wire fch_n_301;
  wire fch_n_302;
  wire fch_n_303;
  wire fch_n_304;
  wire fch_n_305;
  wire fch_n_322;
  wire fch_n_323;
  wire fch_n_324;
  wire fch_n_325;
  wire fch_n_326;
  wire fch_n_327;
  wire fch_n_328;
  wire fch_n_329;
  wire fch_n_330;
  wire fch_n_331;
  wire fch_n_332;
  wire fch_n_333;
  wire fch_n_334;
  wire fch_n_335;
  wire fch_n_336;
  wire fch_n_337;
  wire fch_n_338;
  wire fch_n_339;
  wire fch_n_340;
  wire fch_n_341;
  wire fch_n_342;
  wire fch_n_343;
  wire fch_n_344;
  wire fch_n_345;
  wire fch_n_346;
  wire fch_n_347;
  wire fch_n_348;
  wire fch_n_349;
  wire fch_n_350;
  wire fch_n_351;
  wire fch_n_352;
  wire fch_n_353;
  wire fch_n_354;
  wire fch_n_355;
  wire fch_n_356;
  wire fch_n_357;
  wire fch_n_358;
  wire fch_n_359;
  wire fch_n_360;
  wire fch_n_361;
  wire fch_n_362;
  wire fch_n_363;
  wire fch_n_364;
  wire fch_n_365;
  wire fch_n_366;
  wire fch_n_367;
  wire fch_n_368;
  wire fch_n_369;
  wire fch_n_37;
  wire fch_n_370;
  wire fch_n_371;
  wire fch_n_372;
  wire fch_n_373;
  wire fch_n_374;
  wire fch_n_375;
  wire fch_n_376;
  wire fch_n_377;
  wire fch_n_378;
  wire fch_n_379;
  wire fch_n_38;
  wire fch_n_380;
  wire fch_n_381;
  wire fch_n_382;
  wire fch_n_383;
  wire fch_n_384;
  wire fch_n_385;
  wire fch_n_386;
  wire fch_n_387;
  wire fch_n_388;
  wire fch_n_389;
  wire fch_n_39;
  wire fch_n_390;
  wire fch_n_391;
  wire fch_n_392;
  wire fch_n_393;
  wire fch_n_394;
  wire fch_n_395;
  wire fch_n_396;
  wire fch_n_397;
  wire fch_n_398;
  wire fch_n_399;
  wire fch_n_400;
  wire fch_n_401;
  wire fch_n_402;
  wire fch_n_403;
  wire fch_n_404;
  wire fch_n_405;
  wire fch_n_406;
  wire fch_n_407;
  wire fch_n_408;
  wire fch_n_409;
  wire fch_n_410;
  wire fch_n_411;
  wire fch_n_412;
  wire fch_n_413;
  wire fch_n_414;
  wire fch_n_415;
  wire fch_n_416;
  wire fch_n_417;
  wire fch_n_418;
  wire fch_n_419;
  wire fch_n_420;
  wire fch_n_421;
  wire fch_n_422;
  wire fch_n_423;
  wire fch_n_424;
  wire fch_n_425;
  wire fch_n_426;
  wire fch_n_427;
  wire fch_n_428;
  wire fch_n_429;
  wire fch_n_430;
  wire fch_n_431;
  wire fch_n_432;
  wire fch_n_433;
  wire fch_n_434;
  wire fch_n_435;
  wire fch_n_436;
  wire fch_n_437;
  wire fch_n_438;
  wire fch_n_439;
  wire fch_n_440;
  wire fch_n_441;
  wire fch_n_442;
  wire fch_n_443;
  wire fch_n_444;
  wire fch_n_445;
  wire fch_n_450;
  wire fch_n_451;
  wire fch_n_452;
  wire fch_n_453;
  wire fch_n_454;
  wire fch_n_455;
  wire fch_n_456;
  wire fch_n_457;
  wire fch_n_458;
  wire fch_n_459;
  wire fch_n_460;
  wire fch_n_461;
  wire fch_n_462;
  wire fch_n_463;
  wire fch_n_464;
  wire fch_n_481;
  wire fch_n_482;
  wire fch_n_483;
  wire fch_n_484;
  wire fch_n_485;
  wire fch_n_486;
  wire fch_n_487;
  wire fch_n_488;
  wire fch_n_489;
  wire fch_n_490;
  wire fch_n_491;
  wire fch_n_492;
  wire fch_n_493;
  wire fch_n_494;
  wire fch_n_495;
  wire fch_n_496;
  wire fch_n_497;
  wire fch_n_498;
  wire fch_n_499;
  wire fch_n_500;
  wire fch_n_501;
  wire fch_n_502;
  wire fch_n_503;
  wire fch_n_504;
  wire fch_n_505;
  wire fch_n_506;
  wire fch_n_507;
  wire fch_n_508;
  wire fch_n_509;
  wire fch_n_510;
  wire fch_n_511;
  wire fch_n_512;
  wire fch_n_513;
  wire fch_n_514;
  wire fch_n_515;
  wire fch_n_516;
  wire fch_n_532;
  wire fch_n_533;
  wire fch_n_534;
  wire fch_n_535;
  wire fch_n_536;
  wire fch_n_537;
  wire fch_n_538;
  wire fch_n_539;
  wire fch_n_540;
  wire fch_n_541;
  wire fch_n_542;
  wire fch_n_543;
  wire fch_n_544;
  wire fch_n_545;
  wire fch_n_546;
  wire fch_n_547;
  wire fch_n_548;
  wire fch_n_549;
  wire fch_n_550;
  wire fch_n_551;
  wire fch_n_552;
  wire fch_n_574;
  wire fch_n_575;
  wire fch_n_576;
  wire fch_n_577;
  wire fch_n_578;
  wire fch_n_579;
  wire fch_n_580;
  wire fch_n_581;
  wire fch_n_582;
  wire fch_n_583;
  wire fch_n_584;
  wire fch_n_585;
  wire fch_n_586;
  wire fch_n_587;
  wire fch_n_588;
  wire fch_n_589;
  wire fch_n_590;
  wire fch_n_591;
  wire fch_n_592;
  wire fch_n_593;
  wire fch_n_594;
  wire fch_n_595;
  wire fch_n_596;
  wire fch_n_597;
  wire fch_n_598;
  wire fch_n_599;
  wire fch_n_600;
  wire fch_n_601;
  wire fch_n_602;
  wire fch_n_603;
  wire fch_n_604;
  wire fch_n_642;
  wire fch_n_645;
  wire fch_n_650;
  wire fch_n_703;
  wire fch_n_704;
  wire fch_n_705;
  wire fch_n_706;
  wire fch_n_707;
  wire fch_n_708;
  wire fch_n_709;
  wire fch_n_710;
  wire fch_n_711;
  wire fch_n_712;
  wire fch_n_713;
  wire fch_n_714;
  wire fch_n_715;
  wire fch_n_716;
  wire fch_n_717;
  wire fch_n_718;
  wire fch_n_719;
  wire fch_n_720;
  wire fch_n_721;
  wire fch_n_722;
  wire fch_n_723;
  wire fch_n_724;
  wire fch_n_725;
  wire fch_n_726;
  wire fch_n_727;
  wire fch_n_728;
  wire fch_n_729;
  wire fch_n_730;
  wire fch_n_731;
  wire fch_n_732;
  wire fch_n_733;
  wire fch_n_734;
  wire fch_n_735;
  wire fch_n_736;
  wire fch_n_737;
  wire fch_n_738;
  wire fch_n_739;
  wire fch_n_740;
  wire fch_n_741;
  wire fch_n_742;
  wire fch_n_743;
  wire fch_n_744;
  wire fch_n_745;
  wire fch_n_746;
  wire fch_n_747;
  wire fch_n_748;
  wire fch_n_749;
  wire fch_n_750;
  wire fch_n_751;
  wire fch_n_752;
  wire fch_n_753;
  wire fch_n_754;
  wire fch_n_755;
  wire fch_n_756;
  wire fch_n_757;
  wire fch_n_758;
  wire fch_n_759;
  wire fch_n_760;
  wire fch_n_761;
  wire fch_n_762;
  wire fch_n_763;
  wire fch_n_764;
  wire fch_n_765;
  wire fch_n_766;
  wire fch_n_767;
  wire fch_n_768;
  wire fch_n_769;
  wire fch_n_770;
  wire fch_n_771;
  wire fch_n_772;
  wire fch_n_773;
  wire fch_n_774;
  wire fch_n_775;
  wire fch_n_776;
  wire fch_n_777;
  wire fch_n_778;
  wire fch_n_779;
  wire fch_n_78;
  wire fch_n_780;
  wire fch_n_781;
  wire fch_n_782;
  wire fch_n_783;
  wire fch_n_784;
  wire fch_n_785;
  wire fch_n_786;
  wire fch_n_787;
  wire fch_n_788;
  wire fch_n_789;
  wire fch_n_790;
  wire fch_n_791;
  wire fch_n_792;
  wire fch_n_793;
  wire fch_n_794;
  wire fch_n_795;
  wire fch_n_796;
  wire fch_n_797;
  wire fch_n_798;
  wire fch_n_799;
  wire fch_n_800;
  wire fch_n_801;
  wire fch_n_802;
  wire fch_n_803;
  wire fch_n_804;
  wire fch_n_805;
  wire fch_n_806;
  wire fch_n_807;
  wire fch_n_808;
  wire fch_n_809;
  wire fch_n_810;
  wire fch_n_811;
  wire fch_n_812;
  wire fch_n_813;
  wire fch_n_814;
  wire fch_n_815;
  wire fch_n_816;
  wire fch_n_817;
  wire fch_n_818;
  wire fch_n_819;
  wire fch_n_820;
  wire fch_n_821;
  wire fch_n_822;
  wire fch_n_823;
  wire fch_n_824;
  wire fch_n_825;
  wire fch_n_826;
  wire fch_n_827;
  wire fch_n_828;
  wire fch_n_829;
  wire fch_n_83;
  wire fch_n_830;
  wire fch_n_831;
  wire fch_n_832;
  wire fch_n_833;
  wire fch_n_834;
  wire fch_n_835;
  wire fch_n_836;
  wire fch_n_837;
  wire fch_n_838;
  wire fch_n_839;
  wire fch_n_84;
  wire fch_n_840;
  wire fch_n_841;
  wire fch_n_842;
  wire fch_n_843;
  wire fch_n_844;
  wire fch_n_845;
  wire fch_n_846;
  wire fch_n_847;
  wire fch_n_848;
  wire fch_n_849;
  wire fch_n_85;
  wire fch_n_850;
  wire fch_n_851;
  wire fch_n_852;
  wire fch_n_853;
  wire fch_n_854;
  wire fch_n_855;
  wire fch_n_856;
  wire fch_n_857;
  wire fch_n_858;
  wire fch_n_859;
  wire fch_n_860;
  wire fch_n_861;
  wire fch_n_862;
  wire fch_n_863;
  wire fch_n_864;
  wire fch_n_865;
  wire fch_n_866;
  wire fch_n_867;
  wire fch_n_868;
  wire fch_n_869;
  wire fch_n_870;
  wire fch_n_871;
  wire fch_n_872;
  wire fch_n_873;
  wire fch_n_874;
  wire fch_n_875;
  wire fch_n_876;
  wire fch_n_877;
  wire fch_n_878;
  wire fch_n_879;
  wire fch_n_88;
  wire fch_n_880;
  wire fch_n_881;
  wire fch_n_882;
  wire fch_n_883;
  wire fch_n_884;
  wire fch_n_885;
  wire fch_n_886;
  wire fch_n_887;
  wire fch_n_888;
  wire fch_n_889;
  wire fch_n_890;
  wire fch_n_891;
  wire fch_n_892;
  wire fch_n_893;
  wire fch_n_894;
  wire fch_n_895;
  wire fch_n_896;
  wire fch_n_897;
  wire fch_n_898;
  wire fch_n_899;
  wire fch_n_900;
  wire fch_n_901;
  wire fch_n_902;
  wire fch_n_903;
  wire fch_n_904;
  wire fch_n_905;
  wire fch_n_906;
  wire fch_n_907;
  wire fch_n_908;
  wire fch_n_909;
  wire fch_n_910;
  wire fch_n_911;
  wire fch_n_912;
  wire fch_n_913;
  wire fch_n_914;
  wire fch_n_915;
  wire fch_n_916;
  wire fch_n_917;
  wire fch_n_918;
  wire fch_n_919;
  wire fch_n_920;
  wire fch_n_921;
  wire fch_n_922;
  wire fch_n_923;
  wire fch_n_924;
  wire fch_n_925;
  wire fch_n_926;
  wire fch_n_927;
  wire fch_n_928;
  wire fch_n_929;
  wire fch_n_930;
  wire fch_n_931;
  wire fch_n_932;
  wire fch_n_933;
  wire fch_n_934;
  wire fch_n_935;
  wire fch_n_936;
  wire fch_n_937;
  wire fch_n_938;
  wire fch_n_939;
  wire fch_n_940;
  wire fch_n_941;
  wire fch_n_942;
  wire fch_n_943;
  wire fch_n_944;
  wire fch_n_945;
  wire fch_n_946;
  wire fch_n_947;
  wire fch_n_948;
  wire fch_n_949;
  wire fch_n_950;
  wire fch_n_951;
  wire fch_n_952;
  wire fch_n_953;
  wire fch_n_954;
  wire fch_n_955;
  wire fch_n_956;
  wire fch_n_957;
  wire fch_n_958;
  wire fch_n_959;
  wire fch_n_960;
  wire fch_n_961;
  wire fch_n_962;
  wire fch_n_963;
  wire fch_n_964;
  wire fch_n_965;
  wire fch_n_966;
  wire fch_n_967;
  wire fch_n_968;
  wire fch_n_969;
  wire fch_n_970;
  wire fch_n_971;
  wire fch_n_972;
  wire fch_n_973;
  wire fch_n_974;
  wire fch_n_975;
  wire fch_n_976;
  wire fch_n_977;
  wire fch_n_978;
  wire fch_n_979;
  wire fch_n_980;
  wire fch_n_981;
  wire fch_n_982;
  wire fch_n_983;
  wire fch_n_984;
  wire fch_n_985;
  wire fch_n_986;
  wire fch_n_987;
  wire fch_n_988;
  wire fch_n_989;
  wire fch_n_990;
  wire fch_n_991;
  wire fch_n_992;
  wire fch_n_993;
  wire fch_n_994;
  wire fch_n_995;
  wire fch_n_996;
  wire fch_n_997;
  wire fch_n_998;
  wire fch_n_999;
  wire [15:13]fch_pc;
  wire [15:0]fch_pc0;
  wire [15:0]fch_pc1;
  (* DONT_TOUCH *) wire fch_term;
  wire [15:0]fdat;
  wire [15:0]fdatx;
  wire [21:21]ir0_id;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [15:1]\ivec/p_0_in ;
  wire [15:0]\ivec/p_1_in ;
  wire [21:21]lir_id_0;
  wire mem_n_0;
  wire mem_n_1;
  wire mem_n_10;
  wire mem_n_11;
  wire mem_n_12;
  wire mem_n_13;
  wire mem_n_14;
  wire mem_n_15;
  wire mem_n_18;
  wire mem_n_19;
  wire mem_n_2;
  wire mem_n_20;
  wire mem_n_22;
  wire mem_n_23;
  wire mem_n_24;
  wire mem_n_25;
  wire mem_n_26;
  wire mem_n_27;
  wire mem_n_28;
  wire mem_n_29;
  wire mem_n_3;
  wire mem_n_30;
  wire mem_n_31;
  wire mem_n_32;
  wire mem_n_33;
  wire mem_n_34;
  wire mem_n_35;
  wire mem_n_36;
  wire mem_n_37;
  wire mem_n_38;
  wire mem_n_4;
  wire mem_n_5;
  wire mem_n_6;
  wire mem_n_7;
  wire mem_n_8;
  wire mem_n_9;
  wire [15:0]p_2_in;
  wire [15:13]p_2_in_4;
  wire [15:0]\pcnt/p_1_in ;
  wire \rctl/p_2_in ;
  wire [15:0]\rctl/rgf_c0bus_wb ;
  wire [15:0]\rctl/rgf_c1bus_wb ;
  wire [2:0]\rctl/rgf_selc0_rn_wb ;
  wire \rctl/rgf_selc0_stat ;
  wire [1:0]\rctl/rgf_selc0_wb ;
  wire [2:0]\rctl/rgf_selc1_rn_wb ;
  wire \rctl/rgf_selc1_stat ;
  wire [1:0]\rctl/rgf_selc1_wb ;
  wire rgf_iv_ve;
  wire rgf_n_10;
  wire rgf_n_11;
  wire rgf_n_12;
  wire rgf_n_13;
  wire rgf_n_14;
  wire rgf_n_15;
  wire rgf_n_159;
  wire rgf_n_16;
  wire rgf_n_160;
  wire rgf_n_161;
  wire rgf_n_165;
  wire rgf_n_166;
  wire rgf_n_169;
  wire rgf_n_17;
  wire rgf_n_170;
  wire rgf_n_171;
  wire rgf_n_172;
  wire rgf_n_173;
  wire rgf_n_174;
  wire rgf_n_175;
  wire rgf_n_176;
  wire rgf_n_177;
  wire rgf_n_178;
  wire rgf_n_179;
  wire rgf_n_18;
  wire rgf_n_180;
  wire rgf_n_181;
  wire rgf_n_182;
  wire rgf_n_183;
  wire rgf_n_186;
  wire rgf_n_187;
  wire rgf_n_188;
  wire rgf_n_189;
  wire rgf_n_19;
  wire rgf_n_190;
  wire rgf_n_191;
  wire rgf_n_192;
  wire rgf_n_193;
  wire rgf_n_194;
  wire rgf_n_195;
  wire rgf_n_196;
  wire rgf_n_197;
  wire rgf_n_198;
  wire rgf_n_199;
  wire rgf_n_2;
  wire rgf_n_20;
  wire rgf_n_200;
  wire rgf_n_201;
  wire rgf_n_21;
  wire rgf_n_218;
  wire rgf_n_219;
  wire rgf_n_22;
  wire rgf_n_220;
  wire rgf_n_221;
  wire rgf_n_222;
  wire rgf_n_223;
  wire rgf_n_224;
  wire rgf_n_225;
  wire rgf_n_226;
  wire rgf_n_227;
  wire rgf_n_228;
  wire rgf_n_229;
  wire rgf_n_23;
  wire rgf_n_230;
  wire rgf_n_231;
  wire rgf_n_232;
  wire rgf_n_233;
  wire rgf_n_234;
  wire rgf_n_235;
  wire rgf_n_236;
  wire rgf_n_237;
  wire rgf_n_238;
  wire rgf_n_239;
  wire rgf_n_24;
  wire rgf_n_240;
  wire rgf_n_241;
  wire rgf_n_242;
  wire rgf_n_243;
  wire rgf_n_244;
  wire rgf_n_245;
  wire rgf_n_246;
  wire rgf_n_247;
  wire rgf_n_248;
  wire rgf_n_249;
  wire rgf_n_25;
  wire rgf_n_250;
  wire rgf_n_251;
  wire rgf_n_252;
  wire rgf_n_253;
  wire rgf_n_254;
  wire rgf_n_255;
  wire rgf_n_256;
  wire rgf_n_257;
  wire rgf_n_258;
  wire rgf_n_259;
  wire rgf_n_26;
  wire rgf_n_260;
  wire rgf_n_261;
  wire rgf_n_262;
  wire rgf_n_263;
  wire rgf_n_264;
  wire rgf_n_265;
  wire rgf_n_266;
  wire rgf_n_267;
  wire rgf_n_268;
  wire rgf_n_269;
  wire rgf_n_27;
  wire rgf_n_270;
  wire rgf_n_271;
  wire rgf_n_272;
  wire rgf_n_273;
  wire rgf_n_274;
  wire rgf_n_275;
  wire rgf_n_276;
  wire rgf_n_277;
  wire rgf_n_278;
  wire rgf_n_279;
  wire rgf_n_28;
  wire rgf_n_280;
  wire rgf_n_281;
  wire rgf_n_282;
  wire rgf_n_283;
  wire rgf_n_284;
  wire rgf_n_285;
  wire rgf_n_286;
  wire rgf_n_287;
  wire rgf_n_288;
  wire rgf_n_289;
  wire rgf_n_29;
  wire rgf_n_290;
  wire rgf_n_291;
  wire rgf_n_292;
  wire rgf_n_293;
  wire rgf_n_294;
  wire rgf_n_295;
  wire rgf_n_296;
  wire rgf_n_297;
  wire rgf_n_298;
  wire rgf_n_299;
  wire rgf_n_3;
  wire rgf_n_30;
  wire rgf_n_300;
  wire rgf_n_301;
  wire rgf_n_302;
  wire rgf_n_303;
  wire rgf_n_304;
  wire rgf_n_305;
  wire rgf_n_306;
  wire rgf_n_307;
  wire rgf_n_308;
  wire rgf_n_309;
  wire rgf_n_31;
  wire rgf_n_310;
  wire rgf_n_311;
  wire rgf_n_312;
  wire rgf_n_313;
  wire rgf_n_314;
  wire rgf_n_316;
  wire rgf_n_317;
  wire rgf_n_318;
  wire rgf_n_319;
  wire rgf_n_32;
  wire rgf_n_320;
  wire rgf_n_321;
  wire rgf_n_322;
  wire rgf_n_323;
  wire rgf_n_33;
  wire rgf_n_334;
  wire rgf_n_335;
  wire rgf_n_336;
  wire rgf_n_337;
  wire rgf_n_338;
  wire rgf_n_339;
  wire rgf_n_34;
  wire rgf_n_340;
  wire rgf_n_35;
  wire rgf_n_357;
  wire rgf_n_358;
  wire rgf_n_359;
  wire rgf_n_36;
  wire rgf_n_360;
  wire rgf_n_361;
  wire rgf_n_362;
  wire rgf_n_363;
  wire rgf_n_364;
  wire rgf_n_365;
  wire rgf_n_366;
  wire rgf_n_367;
  wire rgf_n_368;
  wire rgf_n_369;
  wire rgf_n_37;
  wire rgf_n_370;
  wire rgf_n_371;
  wire rgf_n_372;
  wire rgf_n_373;
  wire rgf_n_374;
  wire rgf_n_375;
  wire rgf_n_376;
  wire rgf_n_377;
  wire rgf_n_378;
  wire rgf_n_379;
  wire rgf_n_38;
  wire rgf_n_380;
  wire rgf_n_381;
  wire rgf_n_382;
  wire rgf_n_383;
  wire rgf_n_384;
  wire rgf_n_385;
  wire rgf_n_386;
  wire rgf_n_387;
  wire rgf_n_388;
  wire rgf_n_389;
  wire rgf_n_39;
  wire rgf_n_390;
  wire rgf_n_391;
  wire rgf_n_392;
  wire rgf_n_393;
  wire rgf_n_394;
  wire rgf_n_395;
  wire rgf_n_396;
  wire rgf_n_397;
  wire rgf_n_398;
  wire rgf_n_399;
  wire rgf_n_4;
  wire rgf_n_40;
  wire rgf_n_400;
  wire rgf_n_401;
  wire rgf_n_402;
  wire rgf_n_403;
  wire rgf_n_404;
  wire rgf_n_405;
  wire rgf_n_406;
  wire rgf_n_407;
  wire rgf_n_408;
  wire rgf_n_409;
  wire rgf_n_41;
  wire rgf_n_410;
  wire rgf_n_411;
  wire rgf_n_412;
  wire rgf_n_413;
  wire rgf_n_414;
  wire rgf_n_415;
  wire rgf_n_416;
  wire rgf_n_417;
  wire rgf_n_418;
  wire rgf_n_419;
  wire rgf_n_42;
  wire rgf_n_420;
  wire rgf_n_421;
  wire rgf_n_422;
  wire rgf_n_423;
  wire rgf_n_424;
  wire rgf_n_425;
  wire rgf_n_426;
  wire rgf_n_427;
  wire rgf_n_428;
  wire rgf_n_429;
  wire rgf_n_43;
  wire rgf_n_430;
  wire rgf_n_431;
  wire rgf_n_432;
  wire rgf_n_433;
  wire rgf_n_434;
  wire rgf_n_435;
  wire rgf_n_436;
  wire rgf_n_437;
  wire rgf_n_438;
  wire rgf_n_439;
  wire rgf_n_44;
  wire rgf_n_440;
  wire rgf_n_441;
  wire rgf_n_442;
  wire rgf_n_443;
  wire rgf_n_444;
  wire rgf_n_445;
  wire rgf_n_446;
  wire rgf_n_447;
  wire rgf_n_448;
  wire rgf_n_449;
  wire rgf_n_45;
  wire rgf_n_450;
  wire rgf_n_46;
  wire rgf_n_47;
  wire rgf_n_471;
  wire rgf_n_472;
  wire rgf_n_473;
  wire rgf_n_474;
  wire rgf_n_475;
  wire rgf_n_476;
  wire rgf_n_477;
  wire rgf_n_478;
  wire rgf_n_479;
  wire rgf_n_48;
  wire rgf_n_480;
  wire rgf_n_481;
  wire rgf_n_482;
  wire rgf_n_483;
  wire rgf_n_484;
  wire rgf_n_485;
  wire rgf_n_486;
  wire rgf_n_487;
  wire rgf_n_488;
  wire rgf_n_489;
  wire rgf_n_49;
  wire rgf_n_490;
  wire rgf_n_491;
  wire rgf_n_492;
  wire rgf_n_493;
  wire rgf_n_495;
  wire rgf_n_496;
  wire rgf_n_497;
  wire rgf_n_498;
  wire rgf_n_499;
  wire rgf_n_5;
  wire rgf_n_50;
  wire rgf_n_500;
  wire rgf_n_501;
  wire rgf_n_502;
  wire rgf_n_503;
  wire rgf_n_504;
  wire rgf_n_505;
  wire rgf_n_506;
  wire rgf_n_507;
  wire rgf_n_508;
  wire rgf_n_509;
  wire rgf_n_51;
  wire rgf_n_510;
  wire rgf_n_511;
  wire rgf_n_512;
  wire rgf_n_513;
  wire rgf_n_514;
  wire rgf_n_515;
  wire rgf_n_516;
  wire rgf_n_517;
  wire rgf_n_518;
  wire rgf_n_519;
  wire rgf_n_52;
  wire rgf_n_520;
  wire rgf_n_521;
  wire rgf_n_522;
  wire rgf_n_523;
  wire rgf_n_53;
  wire rgf_n_54;
  wire rgf_n_55;
  wire rgf_n_56;
  wire rgf_n_569;
  wire rgf_n_57;
  wire rgf_n_570;
  wire rgf_n_571;
  wire rgf_n_572;
  wire rgf_n_573;
  wire rgf_n_574;
  wire rgf_n_575;
  wire rgf_n_576;
  wire rgf_n_577;
  wire rgf_n_578;
  wire rgf_n_579;
  wire rgf_n_58;
  wire rgf_n_580;
  wire rgf_n_581;
  wire rgf_n_582;
  wire rgf_n_583;
  wire rgf_n_584;
  wire rgf_n_585;
  wire rgf_n_586;
  wire rgf_n_587;
  wire rgf_n_588;
  wire rgf_n_589;
  wire rgf_n_59;
  wire rgf_n_590;
  wire rgf_n_591;
  wire rgf_n_592;
  wire rgf_n_593;
  wire rgf_n_594;
  wire rgf_n_595;
  wire rgf_n_6;
  wire rgf_n_60;
  wire rgf_n_61;
  wire rgf_n_62;
  wire rgf_n_63;
  wire rgf_n_64;
  wire rgf_n_65;
  wire rgf_n_66;
  wire rgf_n_67;
  wire rgf_n_68;
  wire rgf_n_69;
  wire rgf_n_7;
  wire rgf_n_70;
  wire rgf_n_71;
  wire rgf_n_72;
  wire rgf_n_73;
  wire rgf_n_74;
  wire rgf_n_75;
  wire rgf_n_76;
  wire rgf_n_77;
  wire rgf_n_78;
  wire rgf_n_79;
  wire rgf_n_8;
  wire rgf_n_80;
  wire rgf_n_81;
  wire rgf_n_82;
  wire rgf_n_83;
  wire rgf_n_84;
  wire rgf_n_85;
  wire rgf_n_86;
  wire rgf_n_87;
  wire rgf_n_88;
  wire rgf_n_89;
  wire rgf_n_9;
  wire rgf_n_90;
  wire rgf_n_91;
  wire rgf_n_92;
  wire rgf_n_93;
  wire [15:0]rgf_pc;
  wire rgf_sr_dr;
  wire [3:0]rgf_sr_flag;
  wire [1:0]rgf_sr_ie;
  wire rgf_sr_ml;
  wire rgf_sr_sd;
  wire [15:0]rgf_tr;
  wire rst_n;
  wire [0:0]\sptr/data3 ;
  wire [0:0]\sptr/p_0_in ;
  wire [1:0]sr_bank;
  wire [15:0]\sreg/p_0_in ;
  wire [7:0]\sreg/p_2_in ;
  wire [2:0]stat;
  wire [2:0]stat_2;
  wire [1:0]stat_nx;
  wire [2:0]stat_nx_3;
  wire \treg/p_0_in ;
  wire [15:0]\treg/p_1_in ;

  mcss_alu alu0
       (.DI({fch_n_578,fch_n_579,fch_n_580}),
        .O({alu0_n_0,alu0_n_1,alu0_n_2,alu0_n_3}),
        .S({fch_n_581,fch_n_582,fch_n_583,fch_n_584}),
        .\rgf_c0bus_wb[4]_i_17 ({fch_n_585,fch_n_586,fch_n_587,fch_n_588}),
        .\rgf_c0bus_wb[4]_i_17_0 ({fch_n_589,fch_n_590,fch_n_591,fch_n_592}),
        .\rgf_c0bus_wb[8]_i_5 ({fch_n_593,fch_n_594,fch_n_595,fch_n_596}),
        .\rgf_c0bus_wb[8]_i_5_0 ({fch_n_597,fch_n_598,fch_n_599,fch_n_600}),
        .\rgf_c0bus_wb_reg[15] ({fch_n_546,fch_n_547,fch_n_548,fch_n_549}),
        .\rgf_c0bus_wb_reg[15]_0 ({rgf_n_511,fch_n_543,fch_n_544,fch_n_545}),
        .\sr[4]_i_206 (alu0_n_17),
        .\sr[6]_i_8 (fch_n_550),
        .\sr[6]_i_8_0 ({fch_n_551,fch_n_552}),
        .tout__1_carry__0_i_8({alu0_n_4,alu0_n_5,alu0_n_6,alu0_n_7}),
        .tout__1_carry__1_i_8({alu0_n_8,alu0_n_9,alu0_n_10,alu0_n_11}),
        .tout__1_carry__2_i_8({\art/p_0_in ,alu0_n_13,alu0_n_14,alu0_n_15}),
        .tout__1_carry__3_i_3__0(\art/add/tout ));
  mcss_alu_0 alu1
       (.DI({fch_n_536,fch_n_537,fch_n_538}),
        .O({alu1_n_0,alu1_n_1,alu1_n_2,alu1_n_3}),
        .S({fch_n_532,fch_n_533,fch_n_534,fch_n_535}),
        .\rgf_c1bus_wb[4]_i_5 ({rgf_n_512,rgf_n_513,fch_n_601,fch_n_602}),
        .\rgf_c1bus_wb[4]_i_5_0 ({rgf_n_514,rgf_n_515,fch_n_603,fch_n_604}),
        .\rgf_c1bus_wb[8]_i_4 ({rgf_n_516,rgf_n_517,rgf_n_518,rgf_n_519}),
        .\rgf_c1bus_wb[8]_i_4_0 ({rgf_n_520,rgf_n_521,rgf_n_522,rgf_n_523}),
        .\rgf_c1bus_wb_reg[15] ({fch_n_542,rgf_n_508,rgf_n_509,rgf_n_510}),
        .\rgf_c1bus_wb_reg[15]_0 ({rgf_n_504,rgf_n_505,rgf_n_506,rgf_n_507}),
        .\sr[4]_i_123 (alu1_n_17),
        .\sr[6]_i_2 (fch_n_541),
        .\sr[6]_i_2_0 ({fch_n_539,fch_n_540}),
        .tout__1_carry__0_i_8__0({alu1_n_4,alu1_n_5,alu1_n_6,alu1_n_7}),
        .tout__1_carry__1_i_8__0({alu1_n_8,alu1_n_9,alu1_n_10,alu1_n_11}),
        .tout__1_carry__2_i_8__0({\art/p_0_in_1 ,alu1_n_13,alu1_n_14,alu1_n_15}),
        .tout__1_carry__3_i_3(\art/add/tout_0 ));
  mcss_fsm ctl0
       (.D(stat_nx_3),
        .Q(stat),
        .SR(\treg/p_0_in ),
        .brdy(brdy),
        .\ccmd[4]_INST_0_i_2 (fch_n_258),
        .clk(clk),
        .crdy(crdy),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .out({fch_ir0[15:9],fch_ir0[7],fch_ir0[2:0]}),
        .rgf_sr_dr(rgf_sr_dr),
        .\stat_reg[0]_0 (ctl0_n_5),
        .\stat_reg[0]_1 (ctl0_n_6),
        .\stat_reg[0]_10 (ctl0_n_22),
        .\stat_reg[0]_11 (ctl0_n_23),
        .\stat_reg[0]_12 (ctl0_n_24),
        .\stat_reg[0]_13 (ctl0_n_28),
        .\stat_reg[0]_14 (fch_n_303),
        .\stat_reg[0]_15 (fch_n_242),
        .\stat_reg[0]_16 (ctl1_n_21),
        .\stat_reg[0]_2 (ctl0_n_7),
        .\stat_reg[0]_3 (ctl0_n_8),
        .\stat_reg[0]_4 (ctl0_n_10),
        .\stat_reg[0]_5 (ctl0_n_15),
        .\stat_reg[0]_6 (ctl0_n_16),
        .\stat_reg[0]_7 (ctl0_n_17),
        .\stat_reg[0]_8 (ctl0_n_18),
        .\stat_reg[0]_9 (ctl0_n_21),
        .\stat_reg[1]_0 (ctl0_n_1),
        .\stat_reg[1]_1 (ctl0_n_9),
        .\stat_reg[1]_2 (ctl0_n_11),
        .\stat_reg[1]_3 (ctl0_n_13),
        .\stat_reg[1]_4 (ctl0_n_14),
        .\stat_reg[1]_5 (ctl0_n_25),
        .\stat_reg[1]_6 (ctl0_n_26),
        .\stat_reg[1]_7 (rgf_n_477),
        .\stat_reg[1]_8 (fch_n_304),
        .\stat_reg[2]_0 (ctl0_n_0),
        .\stat_reg[2]_1 (ctl0_n_12),
        .\stat_reg[2]_2 (ctl0_n_19),
        .\stat_reg[2]_3 (ctl0_n_20),
        .\stat_reg[2]_4 (ctl0_n_27));
  mcss_fsm_1 ctl1
       (.D(stat_nx),
        .Q(stat_2),
        .SR(\treg/p_0_in ),
        .brdy(brdy),
        .brdy_0(ctl1_n_19),
        .clk(clk),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .out({fch_ir1[15:9],fch_ir1[2:0]}),
        .\rgf_selc1_rn_wb_reg[0] (fch_n_284),
        .\sp[15]_i_6 (mem_n_18),
        .\stat_reg[0]_0 (ctl1_n_6),
        .\stat_reg[0]_1 (ctl1_n_7),
        .\stat_reg[0]_2 (ctl1_n_12),
        .\stat_reg[0]_3 (ctl1_n_14),
        .\stat_reg[0]_4 (ctl1_n_15),
        .\stat_reg[0]_5 (ctl1_n_20),
        .\stat_reg[1]_0 (ctl1_n_8),
        .\stat_reg[1]_1 (ctl1_n_9),
        .\stat_reg[1]_2 (ctl1_n_10),
        .\stat_reg[1]_3 (ctl1_n_11),
        .\stat_reg[1]_4 (ctl1_n_13),
        .\stat_reg[1]_5 (ctl1_n_16),
        .\stat_reg[1]_6 (ctl1_n_17),
        .\stat_reg[1]_7 (ctl1_n_18),
        .\stat_reg[1]_8 (ctl1_n_22),
        .\stat_reg[2]_0 (ctl1_n_0),
        .\stat_reg[2]_1 (ctl1_n_1),
        .\stat_reg[2]_2 (ctl1_n_5),
        .\stat_reg[2]_3 (ctl1_n_21),
        .\stat_reg[2]_4 (fch_n_293),
        .\stat_reg[2]_5 (fch_n_294),
        .\stat_reg[2]_6 (fch_n_295),
        .\stat_reg[2]_7 (fch_n_289),
        .\stat_reg[2]_8 (mem_n_15));
  mcss_fch fch
       (.D(fch_pc),
        .DI({fch_n_536,fch_n_537,fch_n_538}),
        .E(fch_n_429),
        .O({fch_n_37,fch_n_38,fch_n_39}),
        .Q(\rctl/rgf_c1bus_wb ),
        .S(rgf_n_483),
        .SR(\treg/p_0_in ),
        .a0bus_0(a0bus_0),
        .a0bus_sel_0({a0bus_sel_0[7],a0bus_sel_0[4:3],a0bus_sel_0[0]}),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:0]}),
        .a1bus_0(a1bus_0),
        .a1bus_b02(a1bus_b02),
        .a1bus_sel_0(a1bus_sel_0),
        .a1bus_sel_cr(a1bus_sel_cr),
        .a1bus_sr(a1bus_sr),
        .abus_o(abus_o),
        .b0bus_sel_0(b0bus_sel_0),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b0bus_sr(b0bus_sr),
        .b1bus_b02(b1bus_b02),
        .b1bus_sel_cr(b1bus_sel_cr),
        .b1bus_sr(b1bus_sr),
        .badr(badr[15:1]),
        .\badr[10]_INST_0_i_2 ({fch_n_593,fch_n_594,fch_n_595,fch_n_596}),
        .\badr[14]_INST_0_i_1 (fch_n_199),
        .\badr[14]_INST_0_i_2 ({fch_n_543,fch_n_544,fch_n_545}),
        .\badr[15]_INST_0_i_1 ({fch_n_539,fch_n_540}),
        .\badr[15]_INST_0_i_114_0 (rgf_n_473),
        .\badr[15]_INST_0_i_1_0 (fch_n_541),
        .\badr[15]_INST_0_i_1_1 (fch_n_542),
        .\badr[15]_INST_0_i_2 (fch_n_230),
        .\badr[15]_INST_0_i_25_0 (rgf_n_472),
        .\badr[15]_INST_0_i_28_0 (ctl1_n_16),
        .\badr[15]_INST_0_i_2_0 ({fch_n_546,fch_n_547,fch_n_548,fch_n_549}),
        .\badr[15]_INST_0_i_2_1 (fch_n_550),
        .\badr[15]_INST_0_i_2_2 ({fch_n_551,fch_n_552}),
        .\badr[1]_INST_0_i_2 (fch_n_231),
        .\badr[2]_INST_0_i_2 ({fch_n_578,fch_n_579,fch_n_580}),
        .\badr[4]_INST_0_i_1 ({fch_n_601,fch_n_602}),
        .\badr[6]_INST_0_i_2 ({fch_n_585,fch_n_586,fch_n_587,fch_n_588}),
        .bank_sel(bank_sel),
        .bbus_o({bbus_o[15:6],bbus_o[4:0]}),
        .\bbus_o[0]_0 (rgf_n_573),
        .\bbus_o[0]_INST_0_i_1_0 (fch_n_232),
        .\bbus_o[1]_0 (rgf_n_572),
        .\bbus_o[1]_INST_0_i_1_0 (fch_n_226),
        .\bbus_o[1]_INST_0_i_1_1 (fch_n_234),
        .\bbus_o[1]_INST_0_i_1_2 (fch_n_235),
        .\bbus_o[2]_0 (rgf_n_571),
        .\bbus_o[2]_INST_0_i_1_0 (fch_n_224),
        .\bbus_o[3]_0 (rgf_n_570),
        .\bbus_o[3]_INST_0_i_1_0 (fch_n_225),
        .\bbus_o[4]_INST_0_i_49_0 (rgf_n_476),
        .bbus_o_0_sp_1(rgf_n_574),
        .bbus_o_13_sp_1(rgf_n_189),
        .bbus_o_14_sp_1(rgf_n_186),
        .bbus_o_1_sp_1(rgf_n_575),
        .bbus_o_2_sp_1(rgf_n_576),
        .bbus_o_3_sp_1(rgf_n_577),
        .bbus_o_6_sp_1(rgf_n_219),
        .bbus_o_7_sp_1(rgf_n_198),
        .\bcmd[1] (ctl0_n_27),
        .\bcmd[1]_0 (ctl1_n_9),
        .\bcmd[1]_INST_0_0 (fch_n_185),
        .\bcmd[2]_INST_0_0 (fch_n_184),
        .bdatr(bdatr[13:9]),
        .\bdatr[15] (c1bus),
        .bdatw({bdatw[15],bdatw[12:0]}),
        .\bdatw[10]_0 (rgf_n_336),
        .\bdatw[11]_0 (rgf_n_193),
        .\bdatw[11]_INST_0_i_16_0 (fch_n_200),
        .\bdatw[12]_0 (rgf_n_192),
        .\bdatw[15] (rgf_n_323),
        .\bdatw[15]_0 (rgf_n_197),
        .\bdatw[15]_1 (rgf_n_579),
        .\bdatw[15]_2 (rgf_n_580),
        .\bdatw[15]_INST_0_i_67_0 (ctl0_n_11),
        .\bdatw[8]_0 (rgf_n_338),
        .\bdatw[8]_INST_0_i_16_0 (fch_n_191),
        .\bdatw[8]_INST_0_i_16_1 (fch_n_194),
        .\bdatw[8]_INST_0_i_16_2 (fch_n_197),
        .\bdatw[9]_0 (rgf_n_195),
        .\bdatw[9]_INST_0_i_16_0 (fch_n_192),
        .bdatw_10_sp_1(rgf_n_194),
        .bdatw_11_sp_1(rgf_n_335),
        .bdatw_12_sp_1(rgf_n_334),
        .bdatw_5_sp_1(rgf_n_191),
        .bdatw_6_sp_1(rgf_n_188),
        .bdatw_8_sp_1(rgf_n_196),
        .bdatw_9_sp_1(rgf_n_337),
        .brdy(brdy),
        .cbus_i({cbus_i[13:12],cbus_i[9],cbus_i[7:1]}),
        .\cbus_i[15] (c0bus),
        .ccmd(ccmd),
        .\ccmd[0]_INST_0_i_1_0 (ctl0_n_24),
        .\ccmd[0]_INST_0_i_1_1 (rgf_n_474),
        .\ccmd[0]_INST_0_i_1_2 (ctl0_n_23),
        .\ccmd[2]_INST_0_i_2_0 (ctl0_n_1),
        .\ccmd[2]_INST_0_i_3_0 (ctl0_n_22),
        .\ccmd[3]_INST_0_i_3_0 (ctl0_n_25),
        .ccmd_4_sp_1(ctl0_n_10),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .ctl_bcc_take0_fl(ctl_bcc_take0_fl),
        .ctl_bcc_take0_fl_reg_0(ctl0_n_28),
        .ctl_bcc_take1_fl(ctl_bcc_take1_fl),
        .ctl_bcc_take1_fl_reg_0(ctl1_n_20),
        .ctl_fetch0_fl_i_16(rgf_n_478),
        .ctl_fetch0_fl_i_16_0(ctl0_n_20),
        .ctl_fetch0_fl_i_8(ctl0_n_15),
        .ctl_fetch0_fl_reg_0(ctl0_n_8),
        .ctl_fetch0_fl_reg_1(rgf_n_501),
        .ctl_fetch0_fl_reg_2(rgf_n_471),
        .ctl_fetch1_fl_i_16(rgf_n_475),
        .ctl_fetch1_fl_reg_i_6(rgf_n_479),
        .ctl_sela0(ctl_sela0),
        .ctl_sela0_rn({ctl_sela0_rn[2],ctl_sela0_rn[0]}),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .fadr(fadr[12:0]),
        .\fadr[3] (rgf_n_484),
        .\fch_irq_lev[1]_i_2_0 (ctl0_n_6),
        .fch_irq_req(fch_irq_req),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_irq_req_fl_reg_0(fch_n_445),
        .fch_issu1_inferred_i_49_0(mem_n_20),
        .fch_leir_nir_reg(fch_n_167),
        .fch_leir_nir_reg_0(fch_n_273),
        .fch_leir_nir_reg_1(fch_n_276),
        .fch_leir_nir_reg_2(fch_n_277),
        .fch_leir_nir_reg_3(fch_n_278),
        .fch_leir_nir_reg_4(fch_n_279),
        .fch_leir_nir_reg_5(fch_n_280),
        .fch_leir_nir_reg_6(fch_n_281),
        .fch_leir_nir_reg_7(fch_n_282),
        .fch_memacc1(fch_memacc1),
        .fch_term(fch_term),
        .fdat(fdat),
        .fdat_0_sp_1(fch_n_300),
        .fdat_12_sp_1(fch_n_301),
        .fdat_5_sp_1(fch_n_302),
        .fdatx(fdatx),
        .fdatx_14_sp_1(fch_n_299),
        .fdatx_5_sp_1(fch_n_298),
        .\grn[15]_i_3__5 (\rctl/rgf_selc0_wb ),
        .\grn_reg[0] (fch_n_333),
        .\grn_reg[0]_0 (fch_n_358),
        .\grn_reg[0]_1 (fch_n_365),
        .\grn_reg[0]_2 (fch_n_371),
        .\grn_reg[0]_3 (fch_n_376),
        .\grn_reg[0]_4 (fch_n_381),
        .\grn_reg[0]_5 (fch_n_386),
        .\grn_reg[0]_6 (fch_n_391),
        .\grn_reg[0]_7 (fch_n_396),
        .\grn_reg[15] (fch_term),
        .\grn_reg[15]_0 (\rctl/rgf_selc0_rn_wb ),
        .\grn_reg[1] (fch_n_332),
        .\grn_reg[1]_0 (fch_n_357),
        .\grn_reg[1]_1 (fch_n_364),
        .\grn_reg[1]_2 (fch_n_370),
        .\grn_reg[1]_3 (fch_n_375),
        .\grn_reg[1]_4 (fch_n_380),
        .\grn_reg[1]_5 (fch_n_385),
        .\grn_reg[1]_6 (fch_n_390),
        .\grn_reg[1]_7 (fch_n_395),
        .\grn_reg[2] (fch_n_331),
        .\grn_reg[2]_0 (fch_n_356),
        .\grn_reg[2]_1 (fch_n_363),
        .\grn_reg[2]_2 (fch_n_369),
        .\grn_reg[2]_3 (fch_n_374),
        .\grn_reg[2]_4 (fch_n_379),
        .\grn_reg[2]_5 (fch_n_384),
        .\grn_reg[2]_6 (fch_n_389),
        .\grn_reg[2]_7 (fch_n_394),
        .\grn_reg[3] (fch_n_330),
        .\grn_reg[3]_0 (fch_n_355),
        .\grn_reg[3]_1 (fch_n_362),
        .\grn_reg[3]_2 (fch_n_368),
        .\grn_reg[3]_3 (fch_n_373),
        .\grn_reg[3]_4 (fch_n_378),
        .\grn_reg[3]_5 (fch_n_383),
        .\grn_reg[3]_6 (fch_n_388),
        .\grn_reg[3]_7 (fch_n_393),
        .\grn_reg[4] (fch_n_328),
        .\grn_reg[4]_0 (fch_n_353),
        .\grn_reg[4]_1 (fch_n_359),
        .\grn_reg[4]_2 (fch_n_366),
        .\grn_reg[4]_3 (fch_n_372),
        .\grn_reg[4]_4 (fch_n_377),
        .\grn_reg[4]_5 (fch_n_382),
        .\grn_reg[4]_6 (fch_n_387),
        .\grn_reg[4]_7 (fch_n_392),
        .\i_/bbus_o[0]_INST_0_i_18 (rgf_n_503),
        .\i_/bbus_o[4]_INST_0_i_20 ({rgf_n_74,rgf_n_75,rgf_n_76,rgf_n_77,rgf_n_78}),
        .\i_/bbus_o[4]_INST_0_i_20_0 ({rgf_n_79,rgf_n_80,rgf_n_81,rgf_n_82,rgf_n_83}),
        .\i_/bbus_o[4]_INST_0_i_21 ({rgf_n_89,rgf_n_90,rgf_n_91,rgf_n_92,rgf_n_93}),
        .\i_/bbus_o[4]_INST_0_i_21_0 ({rgf_n_84,rgf_n_85,rgf_n_86,rgf_n_87,rgf_n_88}),
        .\i_/bbus_o[4]_INST_0_i_22 ({rgf_n_38,rgf_n_39,rgf_n_40,rgf_n_41,rgf_n_42}),
        .\i_/bbus_o[4]_INST_0_i_22_0 ({rgf_n_33,rgf_n_34,rgf_n_35,rgf_n_36,rgf_n_37}),
        .\i_/bbus_o[4]_INST_0_i_23 ({rgf_n_43,rgf_n_44,rgf_n_45,rgf_n_46,rgf_n_47}),
        .\i_/bbus_o[4]_INST_0_i_23_0 ({rgf_n_53,rgf_n_54,rgf_n_55,rgf_n_56,rgf_n_57}),
        .\i_/bdatw[12]_INST_0_i_64 ({rgf_n_48,rgf_n_49,rgf_n_50,rgf_n_51,rgf_n_52}),
        .\i_/rgf_c1bus_wb[4]_i_86 ({rgf_n_58,rgf_n_59,rgf_n_60,rgf_n_61,rgf_n_62,rgf_n_63,rgf_n_64,rgf_n_65,rgf_n_66,rgf_n_67,rgf_n_68,rgf_n_69,rgf_n_70,rgf_n_71,rgf_n_72,rgf_n_73}),
        .\i_/rgf_c1bus_wb[4]_i_87 ({rgf_n_17,rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22,rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32}),
        .\i_/rgf_c1bus_wb[4]_i_96 ({rgf_n_2,rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6,rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16}),
        .ir0_id(ir0_id),
        .\ir1_id_fl_reg[20]_0 (rgf_n_481),
        .\ir1_id_fl_reg[21]_0 (mem_n_19),
        .irq_lev(irq_lev),
        .irq_vec(irq_vec),
        .\iv_reg[15] (\ivec/p_1_in ),
        .\iv_reg[15]_0 ({\ivec/p_0_in ,rgf_iv_ve}),
        .\nir_id_reg[21]_0 ({lir_id_0,rgf_n_502}),
        .\nir_id_reg[24]_0 (rgf_n_482),
        .out({fch_ir0[15:9],fch_ir0[7],fch_ir0[2:0]}),
        .p_0_in(\bank02/p_0_in ),
        .p_0_in2_in(\bank02/p_0_in2_in ),
        .p_1_in(\bank02/p_1_in ),
        .p_1_in3_in(\bank02/p_1_in3_in ),
        .p_2_in(\rctl/p_2_in ),
        .\pc0_reg[15]_0 (fch_pc0),
        .\pc0_reg[15]_1 (rgf_pc),
        .\pc1_reg[15]_0 (fch_pc1),
        .\pc1_reg[15]_1 ({rgf_n_485,rgf_n_486,rgf_n_487}),
        .\pc_reg[13] (rgf_n_166),
        .\pc_reg[14] (rgf_n_165),
        .\pc_reg[15] (p_2_in_4),
        .\pc_reg[15]_0 (\rctl/rgf_c0bus_wb ),
        .\pc_reg[15]_1 (rgf_n_161),
        .\read_cyc_reg[1] (ctl1_n_10),
        .\read_cyc_reg[1]_0 (ctl0_n_12),
        .\rgf_c0bus_wb[0]_i_2_0 (rgf_n_450),
        .\rgf_c0bus_wb[0]_i_2_1 (rgf_n_403),
        .\rgf_c0bus_wb[10]_i_4_0 (rgf_n_419),
        .\rgf_c0bus_wb[10]_i_4_1 (rgf_n_425),
        .\rgf_c0bus_wb[11]_i_11_0 (fch_n_227),
        .\rgf_c0bus_wb[11]_i_3_0 (fch_n_228),
        .\rgf_c0bus_wb[11]_i_4_0 (rgf_n_378),
        .\rgf_c0bus_wb[11]_i_5_0 (rgf_n_413),
        .\rgf_c0bus_wb[12]_i_2_0 (rgf_n_438),
        .\rgf_c0bus_wb[12]_i_3_0 (rgf_n_402),
        .\rgf_c0bus_wb[12]_i_3_1 (rgf_n_442),
        .\rgf_c0bus_wb[13]_i_10_0 (fch_n_229),
        .\rgf_c0bus_wb[13]_i_2_0 (rgf_n_404),
        .\rgf_c0bus_wb[13]_i_2_1 (rgf_n_386),
        .\rgf_c0bus_wb[13]_i_2_2 (rgf_n_433),
        .\rgf_c0bus_wb[13]_i_4_0 (rgf_n_367),
        .\rgf_c0bus_wb[14]_i_5_0 (rgf_n_371),
        .\rgf_c0bus_wb[15]_i_4_0 (rgf_n_384),
        .\rgf_c0bus_wb[15]_i_4_1 (rgf_n_418),
        .\rgf_c0bus_wb[15]_i_4_2 (rgf_n_409),
        .\rgf_c0bus_wb[15]_i_7_0 (fch_n_222),
        .\rgf_c0bus_wb[15]_i_8_0 (fch_n_505),
        .\rgf_c0bus_wb[1]_i_3_0 (rgf_n_436),
        .\rgf_c0bus_wb[2]_i_2_0 (rgf_n_397),
        .\rgf_c0bus_wb[4]_i_2_0 (rgf_n_407),
        .\rgf_c0bus_wb[4]_i_2_1 (rgf_n_427),
        .\rgf_c0bus_wb[4]_i_3_0 (rgf_n_423),
        .\rgf_c0bus_wb[4]_i_3_1 (rgf_n_416),
        .\rgf_c0bus_wb[4]_i_5_0 (mem_n_33),
        .\rgf_c0bus_wb[4]_i_6_0 (rgf_n_447),
        .\rgf_c0bus_wb[4]_i_6_1 (rgf_n_448),
        .\rgf_c0bus_wb[5]_i_2_0 (rgf_n_390),
        .\rgf_c0bus_wb[5]_i_2_1 (rgf_n_430),
        .\rgf_c0bus_wb[5]_i_3_0 (rgf_n_361),
        .\rgf_c0bus_wb[5]_i_3_1 (rgf_n_364),
        .\rgf_c0bus_wb[5]_i_3_2 (rgf_n_400),
        .\rgf_c0bus_wb[9]_i_3_0 (rgf_n_387),
        .\rgf_c0bus_wb[9]_i_3_1 (rgf_n_388),
        .\rgf_c0bus_wb_reg[0] (mem_n_0),
        .\rgf_c0bus_wb_reg[10] (rgf_n_395),
        .\rgf_c0bus_wb_reg[10]_0 (mem_n_4),
        .\rgf_c0bus_wb_reg[10]_1 (rgf_n_398),
        .\rgf_c0bus_wb_reg[10]_2 (rgf_n_369),
        .\rgf_c0bus_wb_reg[10]_3 (rgf_n_372),
        .\rgf_c0bus_wb_reg[10]_i_17_0 (rgf_n_340),
        .\rgf_c0bus_wb_reg[10]_i_17_1 (rgf_n_498),
        .\rgf_c0bus_wb_reg[10]_i_17_2 (rgf_n_449),
        .\rgf_c0bus_wb_reg[11] (mem_n_5),
        .\rgf_c0bus_wb_reg[11]_0 ({alu0_n_8,alu0_n_9,alu0_n_10,alu0_n_11}),
        .\rgf_c0bus_wb_reg[11]_1 (rgf_n_380),
        .\rgf_c0bus_wb_reg[11]_2 (rgf_n_444),
        .\rgf_c0bus_wb_reg[11]_3 (rgf_n_445),
        .\rgf_c0bus_wb_reg[12] (rgf_n_491),
        .\rgf_c0bus_wb_reg[12]_0 (rgf_n_373),
        .\rgf_c0bus_wb_reg[13] (rgf_n_389),
        .\rgf_c0bus_wb_reg[13]_0 (rgf_n_578),
        .\rgf_c0bus_wb_reg[13]_1 (rgf_n_569),
        .\rgf_c0bus_wb_reg[14] (mem_n_6),
        .\rgf_c0bus_wb_reg[14]_0 (rgf_n_495),
        .\rgf_c0bus_wb_reg[15] ({\art/p_0_in ,alu0_n_13,alu0_n_14,alu0_n_15}),
        .\rgf_c0bus_wb_reg[15]_0 (mem_n_7),
        .\rgf_c0bus_wb_reg[1] (rgf_n_385),
        .\rgf_c0bus_wb_reg[1]_0 (mem_n_30),
        .\rgf_c0bus_wb_reg[2] (rgf_n_393),
        .\rgf_c0bus_wb_reg[2]_0 (rgf_n_496),
        .\rgf_c0bus_wb_reg[2]_1 (mem_n_31),
        .\rgf_c0bus_wb_reg[3] ({alu0_n_0,alu0_n_1,alu0_n_2,alu0_n_3}),
        .\rgf_c0bus_wb_reg[3]_0 (mem_n_2),
        .\rgf_c0bus_wb_reg[4] (rgf_n_365),
        .\rgf_c0bus_wb_reg[4]_0 (rgf_n_497),
        .\rgf_c0bus_wb_reg[4]_1 (rgf_n_440),
        .\rgf_c0bus_wb_reg[4]_2 (rgf_n_360),
        .\rgf_c0bus_wb_reg[5] (rgf_n_223),
        .\rgf_c0bus_wb_reg[5]_0 (mem_n_34),
        .\rgf_c0bus_wb_reg[5]_1 (rgf_n_394),
        .\rgf_c0bus_wb_reg[6] (mem_n_35),
        .\rgf_c0bus_wb_reg[6]_0 (rgf_n_431),
        .\rgf_c0bus_wb_reg[6]_1 (rgf_n_405),
        .\rgf_c0bus_wb_reg[7] (mem_n_36),
        .\rgf_c0bus_wb_reg[7]_0 ({alu0_n_4,alu0_n_5,alu0_n_6,alu0_n_7}),
        .\rgf_c0bus_wb_reg[7]_1 (rgf_n_382),
        .\rgf_c0bus_wb_reg[7]_2 (rgf_n_374),
        .\rgf_c0bus_wb_reg[7]_3 (rgf_n_379),
        .\rgf_c0bus_wb_reg[8] (mem_n_3),
        .\rgf_c0bus_wb_reg[8]_0 (rgf_n_432),
        .\rgf_c0bus_wb_reg[8]_1 (rgf_n_391),
        .\rgf_c0bus_wb_reg[8]_2 (rgf_n_441),
        .\rgf_c0bus_wb_reg[8]_3 (rgf_n_376),
        .\rgf_c0bus_wb_reg[8]_4 (rgf_n_375),
        .\rgf_c0bus_wb_reg[9] (rgf_n_492),
        .\rgf_c0bus_wb_reg[9]_0 (rgf_n_429),
        .\rgf_c0bus_wb_reg[9]_1 (rgf_n_434),
        .\rgf_c0bus_wb_reg[9]_2 (mem_n_1),
        .\rgf_c1bus_wb[0]_i_16_0 (ctl1_n_15),
        .\rgf_c1bus_wb[0]_i_4_0 (rgf_n_230),
        .\rgf_c1bus_wb[0]_i_4_1 (rgf_n_265),
        .\rgf_c1bus_wb[11]_i_3_0 (rgf_n_240),
        .\rgf_c1bus_wb[11]_i_6_0 (rgf_n_306),
        .\rgf_c1bus_wb[13]_i_2_0 (rgf_n_275),
        .\rgf_c1bus_wb[13]_i_5_0 (rgf_n_190),
        .\rgf_c1bus_wb[14]_i_28_0 (rgf_n_587),
        .\rgf_c1bus_wb[14]_i_28_1 (rgf_n_584),
        .\rgf_c1bus_wb[14]_i_28_2 (rgf_n_592),
        .\rgf_c1bus_wb[14]_i_3_0 (rgf_n_187),
        .\rgf_c1bus_wb[14]_i_3_1 (rgf_n_201),
        .\rgf_c1bus_wb[14]_i_53_0 (ctl1_n_8),
        .\rgf_c1bus_wb[15]_i_10_0 (rgf_n_199),
        .\rgf_c1bus_wb[15]_i_14_0 (fch_n_187),
        .\rgf_c1bus_wb[15]_i_14_1 (fch_n_198),
        .\rgf_c1bus_wb[15]_i_4_0 (rgf_n_247),
        .\rgf_c1bus_wb[1]_i_2_0 (rgf_n_293),
        .\rgf_c1bus_wb[1]_i_2_1 (rgf_n_282),
        .\rgf_c1bus_wb[4]_i_11_0 (rgf_n_316),
        .\rgf_c1bus_wb[4]_i_11_1 (rgf_n_317),
        .\rgf_c1bus_wb[4]_i_11_2 (rgf_n_318),
        .\rgf_c1bus_wb[4]_i_4_0 (rgf_n_319),
        .\rgf_c1bus_wb[4]_i_4_1 (rgf_n_314),
        .\rgf_c1bus_wb[4]_i_4_2 (rgf_n_320),
        .\rgf_c1bus_wb[4]_i_4_3 (rgf_n_308),
        .\rgf_c1bus_wb[5]_i_9_0 (rgf_n_588),
        .\rgf_c1bus_wb[5]_i_9_1 (rgf_n_583),
        .\rgf_c1bus_wb[5]_i_9_2 (rgf_n_593),
        .\rgf_c1bus_wb[9]_i_3_0 (rgf_n_234),
        .\rgf_c1bus_wb[9]_i_3_1 (rgf_n_272),
        .\rgf_c1bus_wb[9]_i_3_2 (rgf_n_229),
        .\rgf_c1bus_wb_reg[0] (rgf_n_488),
        .\rgf_c1bus_wb_reg[0]_0 (mem_n_29),
        .\rgf_c1bus_wb_reg[10] (rgf_n_288),
        .\rgf_c1bus_wb_reg[10]_0 (rgf_n_284),
        .\rgf_c1bus_wb_reg[11] ({alu1_n_8,alu1_n_9}),
        .\rgf_c1bus_wb_reg[11]_0 (rgf_n_245),
        .\rgf_c1bus_wb_reg[12] (mem_n_9),
        .\rgf_c1bus_wb_reg[12]_0 (rgf_n_253),
        .\rgf_c1bus_wb_reg[12]_1 (rgf_n_268),
        .\rgf_c1bus_wb_reg[13] (mem_n_13),
        .\rgf_c1bus_wb_reg[13]_0 (rgf_n_226),
        .\rgf_c1bus_wb_reg[13]_1 (rgf_n_276),
        .\rgf_c1bus_wb_reg[13]_2 (rgf_n_281),
        .\rgf_c1bus_wb_reg[13]_3 (rgf_n_590),
        .\rgf_c1bus_wb_reg[13]_4 (rgf_n_581),
        .\rgf_c1bus_wb_reg[13]_5 (rgf_n_595),
        .\rgf_c1bus_wb_reg[13]_6 (rgf_n_227),
        .\rgf_c1bus_wb_reg[14] (mem_n_14),
        .\rgf_c1bus_wb_reg[14]_0 (rgf_n_321),
        .\rgf_c1bus_wb_reg[14]_1 (rgf_n_285),
        .\rgf_c1bus_wb_reg[14]_2 (rgf_n_225),
        .\rgf_c1bus_wb_reg[14]_3 (rgf_n_292),
        .\rgf_c1bus_wb_reg[15] ({\art/p_0_in_1 ,alu1_n_15}),
        .\rgf_c1bus_wb_reg[15]_0 (mem_n_23),
        .\rgf_c1bus_wb_reg[15]_1 (rgf_n_313),
        .\rgf_c1bus_wb_reg[1] (rgf_n_302),
        .\rgf_c1bus_wb_reg[1]_0 (mem_n_28),
        .\rgf_c1bus_wb_reg[1]_1 (rgf_n_271),
        .\rgf_c1bus_wb_reg[2] (mem_n_8),
        .\rgf_c1bus_wb_reg[2]_0 (rgf_n_490),
        .\rgf_c1bus_wb_reg[3] (rgf_n_259),
        .\rgf_c1bus_wb_reg[3]_0 (rgf_n_238),
        .\rgf_c1bus_wb_reg[3]_1 (rgf_n_242),
        .\rgf_c1bus_wb_reg[3]_2 ({alu1_n_0,alu1_n_2,alu1_n_3}),
        .\rgf_c1bus_wb_reg[3]_3 (mem_n_27),
        .\rgf_c1bus_wb_reg[4] (rgf_n_264),
        .\rgf_c1bus_wb_reg[4]_0 (rgf_n_270),
        .\rgf_c1bus_wb_reg[4]_1 (rgf_n_269),
        .\rgf_c1bus_wb_reg[4]_2 (mem_n_26),
        .\rgf_c1bus_wb_reg[5] (rgf_n_224),
        .\rgf_c1bus_wb_reg[5]_0 (mem_n_25),
        .\rgf_c1bus_wb_reg[6] (mem_n_10),
        .\rgf_c1bus_wb_reg[6]_0 (rgf_n_218),
        .\rgf_c1bus_wb_reg[6]_1 (rgf_n_200),
        .\rgf_c1bus_wb_reg[6]_2 (rgf_n_312),
        .\rgf_c1bus_wb_reg[6]_3 (rgf_n_295),
        .\rgf_c1bus_wb_reg[7] (rgf_n_236),
        .\rgf_c1bus_wb_reg[7]_0 (mem_n_24),
        .\rgf_c1bus_wb_reg[7]_1 ({alu1_n_4,alu1_n_6,alu1_n_7}),
        .\rgf_c1bus_wb_reg[7]_2 (rgf_n_243),
        .\rgf_c1bus_wb_reg[7]_3 (rgf_n_241),
        .\rgf_c1bus_wb_reg[8] (mem_n_11),
        .\rgf_c1bus_wb_reg[8]_0 (rgf_n_250),
        .\rgf_c1bus_wb_reg[8]_1 (rgf_n_489),
        .\rgf_c1bus_wb_reg[8]_2 (rgf_n_254),
        .\rgf_c1bus_wb_reg[9] (mem_n_12),
        .\rgf_c1bus_wb_reg[9]_0 (rgf_n_274),
        .\rgf_selc0_rn_wb[0]_i_5_0 (rgf_n_477),
        .\rgf_selc0_rn_wb_reg[0] (stat),
        .\rgf_selc0_rn_wb_reg[0]_0 (ctl0_n_9),
        .\rgf_selc0_rn_wb_reg[0]_1 (ctl0_n_26),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .\rgf_selc0_wb[1]_i_4_0 (ctl0_n_5),
        .\rgf_selc0_wb[1]_i_4_1 (rgf_n_500),
        .\rgf_selc1_rn_wb[1]_i_2_0 (ctl1_n_18),
        .\rgf_selc1_rn_wb[1]_i_2_1 (ctl1_n_22),
        .\rgf_selc1_rn_wb_reg[0] (ctl1_n_5),
        .\rgf_selc1_rn_wb_reg[2] (mem_n_37),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg(\pcnt/p_1_in ),
        .rgf_selc1_stat_reg_0(p_2_in),
        .rgf_selc1_stat_reg_1({fch_n_703,fch_n_704,fch_n_705,fch_n_706,fch_n_707,fch_n_708,fch_n_709,fch_n_710,fch_n_711,fch_n_712,fch_n_713,fch_n_714,fch_n_715,fch_n_716,fch_n_717,fch_n_718}),
        .rgf_selc1_stat_reg_10({fch_n_847,fch_n_848,fch_n_849,fch_n_850,fch_n_851,fch_n_852,fch_n_853,fch_n_854,fch_n_855,fch_n_856,fch_n_857,fch_n_858,fch_n_859,fch_n_860,fch_n_861,fch_n_862}),
        .rgf_selc1_stat_reg_11({fch_n_863,fch_n_864,fch_n_865,fch_n_866,fch_n_867,fch_n_868,fch_n_869,fch_n_870,fch_n_871,fch_n_872,fch_n_873,fch_n_874,fch_n_875,fch_n_876,fch_n_877,fch_n_878}),
        .rgf_selc1_stat_reg_12({fch_n_879,fch_n_880,fch_n_881,fch_n_882,fch_n_883,fch_n_884,fch_n_885,fch_n_886,fch_n_887,fch_n_888,fch_n_889,fch_n_890,fch_n_891,fch_n_892,fch_n_893,fch_n_894}),
        .rgf_selc1_stat_reg_13({fch_n_895,fch_n_896,fch_n_897,fch_n_898,fch_n_899,fch_n_900,fch_n_901,fch_n_902,fch_n_903,fch_n_904,fch_n_905,fch_n_906,fch_n_907,fch_n_908,fch_n_909,fch_n_910}),
        .rgf_selc1_stat_reg_14({fch_n_911,fch_n_912,fch_n_913,fch_n_914,fch_n_915,fch_n_916,fch_n_917,fch_n_918,fch_n_919,fch_n_920,fch_n_921,fch_n_922,fch_n_923,fch_n_924,fch_n_925,fch_n_926}),
        .rgf_selc1_stat_reg_15({fch_n_927,fch_n_928,fch_n_929,fch_n_930,fch_n_931,fch_n_932,fch_n_933,fch_n_934,fch_n_935,fch_n_936,fch_n_937,fch_n_938,fch_n_939,fch_n_940,fch_n_941,fch_n_942}),
        .rgf_selc1_stat_reg_16({fch_n_943,fch_n_944,fch_n_945,fch_n_946,fch_n_947,fch_n_948,fch_n_949,fch_n_950,fch_n_951,fch_n_952,fch_n_953,fch_n_954,fch_n_955,fch_n_956,fch_n_957,fch_n_958}),
        .rgf_selc1_stat_reg_17({fch_n_959,fch_n_960,fch_n_961,fch_n_962,fch_n_963,fch_n_964,fch_n_965,fch_n_966,fch_n_967,fch_n_968,fch_n_969,fch_n_970,fch_n_971,fch_n_972,fch_n_973,fch_n_974}),
        .rgf_selc1_stat_reg_18({fch_n_975,fch_n_976,fch_n_977,fch_n_978,fch_n_979,fch_n_980,fch_n_981,fch_n_982,fch_n_983,fch_n_984,fch_n_985,fch_n_986,fch_n_987,fch_n_988,fch_n_989,fch_n_990}),
        .rgf_selc1_stat_reg_19({fch_n_991,fch_n_992,fch_n_993,fch_n_994,fch_n_995,fch_n_996,fch_n_997,fch_n_998,fch_n_999,fch_n_1000,fch_n_1001,fch_n_1002,fch_n_1003,fch_n_1004,fch_n_1005,fch_n_1006}),
        .rgf_selc1_stat_reg_2({fch_n_719,fch_n_720,fch_n_721,fch_n_722,fch_n_723,fch_n_724,fch_n_725,fch_n_726,fch_n_727,fch_n_728,fch_n_729,fch_n_730,fch_n_731,fch_n_732,fch_n_733,fch_n_734}),
        .rgf_selc1_stat_reg_20({fch_n_1007,fch_n_1008,fch_n_1009,fch_n_1010,fch_n_1011,fch_n_1012,fch_n_1013,fch_n_1014,fch_n_1015,fch_n_1016,fch_n_1017,fch_n_1018,fch_n_1019,fch_n_1020,fch_n_1021,fch_n_1022}),
        .rgf_selc1_stat_reg_21({fch_n_1023,fch_n_1024,fch_n_1025,fch_n_1026,fch_n_1027,fch_n_1028,fch_n_1029,fch_n_1030,fch_n_1031,fch_n_1032,fch_n_1033,fch_n_1034,fch_n_1035,fch_n_1036,fch_n_1037,fch_n_1038}),
        .rgf_selc1_stat_reg_22({fch_n_1039,fch_n_1040,fch_n_1041,fch_n_1042,fch_n_1043,fch_n_1044,fch_n_1045,fch_n_1046,fch_n_1047,fch_n_1048,fch_n_1049,fch_n_1050,fch_n_1051,fch_n_1052,fch_n_1053,fch_n_1054}),
        .rgf_selc1_stat_reg_23({fch_n_1055,fch_n_1056,fch_n_1057,fch_n_1058,fch_n_1059,fch_n_1060,fch_n_1061,fch_n_1062,fch_n_1063,fch_n_1064,fch_n_1065,fch_n_1066,fch_n_1067,fch_n_1068,fch_n_1069,fch_n_1070}),
        .rgf_selc1_stat_reg_24({fch_n_1071,fch_n_1072,fch_n_1073,fch_n_1074,fch_n_1075,fch_n_1076,fch_n_1077,fch_n_1078,fch_n_1079,fch_n_1080,fch_n_1081,fch_n_1082,fch_n_1083,fch_n_1084,fch_n_1085,fch_n_1086}),
        .rgf_selc1_stat_reg_25({fch_n_1087,fch_n_1088,fch_n_1089,fch_n_1090,fch_n_1091,fch_n_1092,fch_n_1093,fch_n_1094,fch_n_1095,fch_n_1096,fch_n_1097,fch_n_1098,fch_n_1099,fch_n_1100,fch_n_1101,fch_n_1102}),
        .rgf_selc1_stat_reg_26({fch_n_1103,fch_n_1104,fch_n_1105,fch_n_1106,fch_n_1107,fch_n_1108,fch_n_1109,fch_n_1110,fch_n_1111,fch_n_1112,fch_n_1113,fch_n_1114,fch_n_1115,fch_n_1116,fch_n_1117,fch_n_1118}),
        .rgf_selc1_stat_reg_27({fch_n_1119,fch_n_1120,fch_n_1121,fch_n_1122,fch_n_1123,fch_n_1124,fch_n_1125,fch_n_1126,fch_n_1127,fch_n_1128,fch_n_1129,fch_n_1130,fch_n_1131,fch_n_1132,fch_n_1133,fch_n_1134}),
        .rgf_selc1_stat_reg_28({fch_n_1135,fch_n_1136,fch_n_1137,fch_n_1138,fch_n_1139,fch_n_1140,fch_n_1141,fch_n_1142,fch_n_1143,fch_n_1144,fch_n_1145,fch_n_1146,fch_n_1147,fch_n_1148,fch_n_1149,fch_n_1150}),
        .rgf_selc1_stat_reg_29({fch_n_1151,fch_n_1152,fch_n_1153,fch_n_1154,fch_n_1155,fch_n_1156,fch_n_1157,fch_n_1158,fch_n_1159,fch_n_1160,fch_n_1161,fch_n_1162,fch_n_1163,fch_n_1164,fch_n_1165,fch_n_1166}),
        .rgf_selc1_stat_reg_3({fch_n_735,fch_n_736,fch_n_737,fch_n_738,fch_n_739,fch_n_740,fch_n_741,fch_n_742,fch_n_743,fch_n_744,fch_n_745,fch_n_746,fch_n_747,fch_n_748,fch_n_749,fch_n_750}),
        .rgf_selc1_stat_reg_30({fch_n_1167,fch_n_1168,fch_n_1169,fch_n_1170,fch_n_1171,fch_n_1172,fch_n_1173,fch_n_1174,fch_n_1175,fch_n_1176,fch_n_1177,fch_n_1178,fch_n_1179,fch_n_1180,fch_n_1181,fch_n_1182}),
        .rgf_selc1_stat_reg_31({fch_n_1183,fch_n_1184,fch_n_1185,fch_n_1186,fch_n_1187,fch_n_1188,fch_n_1189,fch_n_1190,fch_n_1191,fch_n_1192,fch_n_1193,fch_n_1194,fch_n_1195,fch_n_1196,fch_n_1197,fch_n_1198}),
        .rgf_selc1_stat_reg_4({fch_n_751,fch_n_752,fch_n_753,fch_n_754,fch_n_755,fch_n_756,fch_n_757,fch_n_758,fch_n_759,fch_n_760,fch_n_761,fch_n_762,fch_n_763,fch_n_764,fch_n_765,fch_n_766}),
        .rgf_selc1_stat_reg_5({fch_n_767,fch_n_768,fch_n_769,fch_n_770,fch_n_771,fch_n_772,fch_n_773,fch_n_774,fch_n_775,fch_n_776,fch_n_777,fch_n_778,fch_n_779,fch_n_780,fch_n_781,fch_n_782}),
        .rgf_selc1_stat_reg_6({fch_n_783,fch_n_784,fch_n_785,fch_n_786,fch_n_787,fch_n_788,fch_n_789,fch_n_790,fch_n_791,fch_n_792,fch_n_793,fch_n_794,fch_n_795,fch_n_796,fch_n_797,fch_n_798}),
        .rgf_selc1_stat_reg_7({fch_n_799,fch_n_800,fch_n_801,fch_n_802,fch_n_803,fch_n_804,fch_n_805,fch_n_806,fch_n_807,fch_n_808,fch_n_809,fch_n_810,fch_n_811,fch_n_812,fch_n_813,fch_n_814}),
        .rgf_selc1_stat_reg_8({fch_n_815,fch_n_816,fch_n_817,fch_n_818,fch_n_819,fch_n_820,fch_n_821,fch_n_822,fch_n_823,fch_n_824,fch_n_825,fch_n_826,fch_n_827,fch_n_828,fch_n_829,fch_n_830}),
        .rgf_selc1_stat_reg_9({fch_n_831,fch_n_832,fch_n_833,fch_n_834,fch_n_835,fch_n_836,fch_n_837,fch_n_838,fch_n_839,fch_n_840,fch_n_841,fch_n_842,fch_n_843,fch_n_844,fch_n_845,fch_n_846}),
        .\rgf_selc1_wb[1]_i_5_0 (rgf_n_499),
        .\rgf_selc1_wb[1]_i_5_1 (ctl1_n_6),
        .\rgf_selc1_wb[1]_i_5_2 (ctl1_n_12),
        .\rgf_selc1_wb_reg[0] (ctl1_n_13),
        .\rgf_selc1_wb_reg[1] (stat_2),
        .\rgf_selc1_wb_reg[1]_0 (ctl1_n_17),
        .rst_n(rst_n),
        .rst_n_0(fch_n_108),
        .rst_n_fl_reg_0({fch_ir1[15:9],fch_ir1[5],fch_ir1[2:0]}),
        .rst_n_fl_reg_1(fch_n_78),
        .rst_n_fl_reg_10(fch_n_439),
        .rst_n_fl_reg_11(fch_n_440),
        .rst_n_fl_reg_12(fch_n_441),
        .rst_n_fl_reg_2(fch_n_258),
        .rst_n_fl_reg_3(fch_n_264),
        .rst_n_fl_reg_4(fch_n_268),
        .rst_n_fl_reg_5(fch_n_269),
        .rst_n_fl_reg_6(fch_n_270),
        .rst_n_fl_reg_7(fch_n_274),
        .rst_n_fl_reg_8(fch_n_275),
        .rst_n_fl_reg_9(fch_n_283),
        .\sp[15]_i_2 (ctl1_n_19),
        .\sp[15]_i_8_0 (ctl0_n_13),
        .\sp_reg[0] (\sptr/data3 ),
        .\sp_reg[0]_0 (\sptr/p_0_in ),
        .\sp_reg[10] (rgf_n_179),
        .\sp_reg[11] (rgf_n_180),
        .\sp_reg[12] (rgf_n_181),
        .\sp_reg[13] (rgf_n_182),
        .\sp_reg[14] (rgf_n_183),
        .\sp_reg[15] ({fch_n_149,fch_n_150,fch_n_151,fch_n_152,fch_n_153,fch_n_154,fch_n_155,fch_n_156,fch_n_157,fch_n_158,fch_n_159,fch_n_160,fch_n_161,fch_n_162,fch_n_163,fch_n_164}),
        .\sp_reg[15]_0 (rgf_n_169),
        .\sp_reg[1] (rgf_n_170),
        .\sp_reg[2] (rgf_n_171),
        .\sp_reg[3] (rgf_n_172),
        .\sp_reg[4] (rgf_n_173),
        .\sp_reg[5] (rgf_n_174),
        .\sp_reg[6] (rgf_n_175),
        .\sp_reg[7] (rgf_n_176),
        .\sp_reg[8] (rgf_n_177),
        .\sp_reg[9] (rgf_n_178),
        .\sr[13]_i_5 (\rctl/rgf_selc1_rn_wb ),
        .\sr[13]_i_5_0 (\rctl/rgf_selc1_wb ),
        .\sr[15]_i_2 (mem_n_38),
        .\sr[3]_i_3 (mem_n_32),
        .\sr[4]_i_100_0 (rgf_n_280),
        .\sr[4]_i_100_1 (rgf_n_278),
        .\sr[4]_i_100_2 (rgf_n_310),
        .\sr[4]_i_102_0 (rgf_n_267),
        .\sr[4]_i_102_1 (rgf_n_589),
        .\sr[4]_i_102_2 (rgf_n_582),
        .\sr[4]_i_102_3 (rgf_n_594),
        .\sr[4]_i_10_0 (rgf_n_228),
        .\sr[4]_i_10_1 (rgf_n_246),
        .\sr[4]_i_10_2 (rgf_n_239),
        .\sr[4]_i_111_0 (rgf_n_262),
        .\sr[4]_i_11_0 (rgf_n_257),
        .\sr[4]_i_127_0 (rgf_n_411),
        .\sr[4]_i_127_1 (rgf_n_412),
        .\sr[4]_i_128 (rgf_n_435),
        .\sr[4]_i_128_0 (rgf_n_428),
        .\sr[4]_i_12_0 (rgf_n_283),
        .\sr[4]_i_15_0 (rgf_n_377),
        .\sr[4]_i_16_0 (rgf_n_368),
        .\sr[4]_i_17_0 (rgf_n_437),
        .\sr[4]_i_17_1 (rgf_n_401),
        .\sr[4]_i_18_0 (rgf_n_399),
        .\sr[4]_i_18_1 (rgf_n_366),
        .\sr[4]_i_18_2 (rgf_n_362),
        .\sr[4]_i_18_3 (rgf_n_363),
        .\sr[4]_i_20_0 (alu0_n_17),
        .\sr[4]_i_25_0 (rgf_n_255),
        .\sr[4]_i_27_0 (rgf_n_266),
        .\sr[4]_i_28_0 (rgf_n_307),
        .\sr[4]_i_28_1 (rgf_n_305),
        .\sr[4]_i_29_0 (rgf_n_273),
        .\sr[4]_i_29_1 (rgf_n_277),
        .\sr[4]_i_29_2 (rgf_n_291),
        .\sr[4]_i_29_3 (rgf_n_303),
        .\sr[4]_i_30_0 (rgf_n_311),
        .\sr[4]_i_30_1 (rgf_n_249),
        .\sr[4]_i_33_0 (rgf_n_248),
        .\sr[4]_i_34_0 (rgf_n_297),
        .\sr[4]_i_35_0 (rgf_n_261),
        .\sr[4]_i_35_1 (rgf_n_244),
        .\sr[4]_i_36_0 (rgf_n_256),
        .\sr[4]_i_36_1 (rgf_n_301),
        .\sr[4]_i_36_2 (rgf_n_263),
        .\sr[4]_i_37_0 (rgf_n_300),
        .\sr[4]_i_39_0 (rgf_n_258),
        .\sr[4]_i_3_0 (alu1_n_17),
        .\sr[4]_i_41_0 (rgf_n_309),
        .\sr[4]_i_43_0 (rgf_n_290),
        .\sr[4]_i_43_1 (rgf_n_289),
        .\sr[4]_i_43_2 (rgf_n_294),
        .\sr[4]_i_44_0 (rgf_n_286),
        .\sr[4]_i_45_0 (rgf_n_298),
        .\sr[4]_i_46_0 (rgf_n_287),
        .\sr[4]_i_46_1 (rgf_n_304),
        .\sr[4]_i_46_2 (rgf_n_296),
        .\sr[4]_i_52_0 (rgf_n_322),
        .\sr[4]_i_53_0 (rgf_n_222),
        .\sr[4]_i_53_1 (rgf_n_220),
        .\sr[4]_i_54_0 (rgf_n_408),
        .\sr[4]_i_54_1 (rgf_n_439),
        .\sr[4]_i_55_0 (rgf_n_446),
        .\sr[4]_i_55_1 (rgf_n_414),
        .\sr[4]_i_55_2 (rgf_n_410),
        .\sr[4]_i_58_0 (rgf_n_424),
        .\sr[4]_i_60_0 (rgf_n_415),
        .\sr[4]_i_60_1 (rgf_n_417),
        .\sr[4]_i_60_2 (rgf_n_421),
        .\sr[4]_i_63_0 (rgf_n_426),
        .\sr[4]_i_63_1 (rgf_n_406),
        .\sr[4]_i_64_0 (rgf_n_370),
        .\sr[4]_i_64_1 (rgf_n_396),
        .\sr[4]_i_65_0 (rgf_n_420),
        .\sr[4]_i_66_0 (rgf_n_392),
        .\sr[4]_i_67_0 (rgf_n_422),
        .\sr[4]_i_68_0 (rgf_n_383),
        .\sr[4]_i_68_1 (rgf_n_443),
        .\sr[4]_i_69_0 (rgf_n_339),
        .\sr[4]_i_6_0 (rgf_n_359),
        .\sr[4]_i_70_0 (rgf_n_358),
        .\sr[4]_i_71_0 (rgf_n_493),
        .\sr[4]_i_72_0 (rgf_n_357),
        .\sr[4]_i_91 (rgf_n_279),
        .\sr[4]_i_98_0 (rgf_n_233),
        .\sr[4]_i_98_1 (rgf_n_232),
        .\sr[4]_i_9_0 (rgf_n_231),
        .\sr[6]_i_16 (rgf_n_586),
        .\sr[6]_i_16_0 (rgf_n_585),
        .\sr[6]_i_16_1 (rgf_n_591),
        .\sr[6]_i_5 (rgf_n_381),
        .\sr[6]_i_5_0 (\art/add/tout ),
        .\sr[6]_i_6_0 (rgf_n_252),
        .\sr[6]_i_6_1 (rgf_n_260),
        .\sr[6]_i_6_2 (rgf_n_251),
        .\sr[6]_i_6_3 (rgf_n_235),
        .\sr[6]_i_9_0 (rgf_n_237),
        .\sr[6]_i_9_1 (rgf_n_299),
        .\sr_reg[0] (fch_n_322),
        .\sr_reg[0]_0 (fch_n_324),
        .\sr_reg[0]_1 (fch_n_325),
        .\sr_reg[0]_10 (fch_n_343),
        .\sr_reg[0]_11 (fch_n_344),
        .\sr_reg[0]_12 (fch_n_345),
        .\sr_reg[0]_13 (fch_n_346),
        .\sr_reg[0]_14 (fch_n_347),
        .\sr_reg[0]_15 (fch_n_348),
        .\sr_reg[0]_16 (fch_n_349),
        .\sr_reg[0]_17 (fch_n_350),
        .\sr_reg[0]_18 (fch_n_351),
        .\sr_reg[0]_19 (fch_n_352),
        .\sr_reg[0]_2 (fch_n_326),
        .\sr_reg[0]_20 (fch_n_397),
        .\sr_reg[0]_21 (fch_n_398),
        .\sr_reg[0]_22 (fch_n_399),
        .\sr_reg[0]_23 (fch_n_400),
        .\sr_reg[0]_24 (fch_n_401),
        .\sr_reg[0]_25 (fch_n_402),
        .\sr_reg[0]_26 (fch_n_403),
        .\sr_reg[0]_27 (fch_n_404),
        .\sr_reg[0]_28 (fch_n_405),
        .\sr_reg[0]_29 (fch_n_406),
        .\sr_reg[0]_3 (fch_n_327),
        .\sr_reg[0]_30 (fch_n_407),
        .\sr_reg[0]_31 (fch_n_408),
        .\sr_reg[0]_32 (fch_n_409),
        .\sr_reg[0]_33 (fch_n_410),
        .\sr_reg[0]_34 (fch_n_411),
        .\sr_reg[0]_35 (fch_n_412),
        .\sr_reg[0]_36 (fch_n_482),
        .\sr_reg[0]_37 (fch_n_483),
        .\sr_reg[0]_38 (fch_n_484),
        .\sr_reg[0]_39 (fch_n_486),
        .\sr_reg[0]_4 (fch_n_334),
        .\sr_reg[0]_40 (fch_n_487),
        .\sr_reg[0]_41 (fch_n_488),
        .\sr_reg[0]_42 (fch_n_490),
        .\sr_reg[0]_43 (fch_n_491),
        .\sr_reg[0]_44 (fch_n_492),
        .\sr_reg[0]_45 (fch_n_494),
        .\sr_reg[0]_46 (fch_n_495),
        .\sr_reg[0]_47 (fch_n_496),
        .\sr_reg[0]_48 (fch_n_498),
        .\sr_reg[0]_49 (fch_n_499),
        .\sr_reg[0]_5 (fch_n_338),
        .\sr_reg[0]_50 (fch_n_500),
        .\sr_reg[0]_51 (fch_n_502),
        .\sr_reg[0]_52 (fch_n_503),
        .\sr_reg[0]_53 (fch_n_504),
        .\sr_reg[0]_54 (fch_n_574),
        .\sr_reg[0]_55 (fch_n_576),
        .\sr_reg[0]_56 (fch_n_577),
        .\sr_reg[0]_57 (fch_n_1199),
        .\sr_reg[0]_58 (fch_n_1200),
        .\sr_reg[0]_59 (fch_n_1201),
        .\sr_reg[0]_6 (fch_n_339),
        .\sr_reg[0]_7 (fch_n_340),
        .\sr_reg[0]_8 (fch_n_341),
        .\sr_reg[0]_9 (fch_n_342),
        .\sr_reg[15] (\sreg/p_0_in ),
        .\sr_reg[15]_0 ({\sreg/p_2_in [7:4],rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,\sreg/p_2_in [0],rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[1] (fch_n_413),
        .\sr_reg[1]_0 (fch_n_414),
        .\sr_reg[1]_1 (fch_n_415),
        .\sr_reg[1]_10 (fch_n_424),
        .\sr_reg[1]_11 (fch_n_425),
        .\sr_reg[1]_12 (fch_n_426),
        .\sr_reg[1]_13 (fch_n_427),
        .\sr_reg[1]_14 (fch_n_481),
        .\sr_reg[1]_15 (fch_n_485),
        .\sr_reg[1]_16 (fch_n_489),
        .\sr_reg[1]_17 (fch_n_493),
        .\sr_reg[1]_18 (fch_n_497),
        .\sr_reg[1]_19 (fch_n_501),
        .\sr_reg[1]_2 (fch_n_416),
        .\sr_reg[1]_20 (fch_n_575),
        .\sr_reg[1]_21 (fch_n_1202),
        .\sr_reg[1]_3 (fch_n_417),
        .\sr_reg[1]_4 (fch_n_418),
        .\sr_reg[1]_5 (fch_n_419),
        .\sr_reg[1]_6 (fch_n_420),
        .\sr_reg[1]_7 (fch_n_421),
        .\sr_reg[1]_8 (fch_n_422),
        .\sr_reg[1]_9 (fch_n_423),
        .\sr_reg[4] (fch_n_289),
        .\sr_reg[4]_0 (fch_n_304),
        .\sr_reg[4]_1 (rgf_n_159),
        .\sr_reg[5] (fch_n_251),
        .\sr_reg[5]_0 (rgf_n_160),
        .\sr_reg[6] (fch_n_195),
        .\sr_reg[6]_0 (fch_n_233),
        .\sr_reg[6]_1 (\art/add/tout_0 ),
        .\stat[0]_i_15_0 (ctl0_n_21),
        .\stat[0]_i_2__1_0 (ctl1_n_7),
        .\stat[0]_i_30_0 (ctl0_n_19),
        .\stat[0]_i_8_0 (ctl0_n_17),
        .\stat[2]_i_2__1 (rgf_n_480),
        .\stat[2]_i_4 (fch_n_146),
        .\stat_reg[0] (fch_n_147),
        .\stat_reg[0]_0 (fch_n_165),
        .\stat_reg[0]_1 (fch_n_166),
        .\stat_reg[0]_10 (fch_n_256),
        .\stat_reg[0]_11 (fch_n_265),
        .\stat_reg[0]_12 (fch_n_267),
        .\stat_reg[0]_13 (fch_n_271),
        .\stat_reg[0]_14 (fch_n_272),
        .\stat_reg[0]_15 (\bctl/ctl/stat_nx ),
        .\stat_reg[0]_16 (fch_n_293),
        .\stat_reg[0]_17 (fch_n_294),
        .\stat_reg[0]_18 (fch_n_295),
        .\stat_reg[0]_19 (fch_n_323),
        .\stat_reg[0]_2 (fch_n_203),
        .\stat_reg[0]_20 (fch_n_329),
        .\stat_reg[0]_21 (fch_n_354),
        .\stat_reg[0]_22 (fch_n_361),
        .\stat_reg[0]_23 (fch_n_367),
        .\stat_reg[0]_24 (fch_n_430),
        .\stat_reg[0]_25 (fch_n_431),
        .\stat_reg[0]_26 (fch_n_432),
        .\stat_reg[0]_27 (fch_n_433),
        .\stat_reg[0]_28 (fch_n_434),
        .\stat_reg[0]_29 (fch_n_435),
        .\stat_reg[0]_3 (fch_n_221),
        .\stat_reg[0]_30 (fch_n_436),
        .\stat_reg[0]_31 (fch_n_437),
        .\stat_reg[0]_32 (fch_n_438),
        .\stat_reg[0]_33 (fch_n_442),
        .\stat_reg[0]_34 (fch_n_506),
        .\stat_reg[0]_35 (fch_n_507),
        .\stat_reg[0]_36 (fch_n_508),
        .\stat_reg[0]_37 (fch_n_509),
        .\stat_reg[0]_38 (fch_n_510),
        .\stat_reg[0]_39 (fch_n_511),
        .\stat_reg[0]_4 (stat_nx_3),
        .\stat_reg[0]_40 (fch_n_512),
        .\stat_reg[0]_41 (fch_n_513),
        .\stat_reg[0]_42 (fch_n_514),
        .\stat_reg[0]_43 (fch_n_515),
        .\stat_reg[0]_44 (fch_n_516),
        .\stat_reg[0]_45 (fch_n_642),
        .\stat_reg[0]_46 (fch_n_645),
        .\stat_reg[0]_47 (fch_n_650),
        .\stat_reg[0]_48 (mem_n_18),
        .\stat_reg[0]_49 (ctl0_n_0),
        .\stat_reg[0]_5 (fch_n_248),
        .\stat_reg[0]_50 (ctl0_n_14),
        .\stat_reg[0]_51 (ctl0_n_16),
        .\stat_reg[0]_52 (mem_n_22),
        .\stat_reg[0]_53 (ctl1_n_0),
        .\stat_reg[0]_54 (ctl1_n_1),
        .\stat_reg[0]_55 (mem_n_15),
        .\stat_reg[0]_56 (\bctl/ctl/p_0_in ),
        .\stat_reg[0]_6 (fch_n_250),
        .\stat_reg[0]_7 (fch_n_253),
        .\stat_reg[0]_8 (fch_n_254),
        .\stat_reg[0]_9 (fch_n_255),
        .\stat_reg[1] (fch_n_148),
        .\stat_reg[1]_0 (fch_n_168),
        .\stat_reg[1]_1 (fch_n_205),
        .\stat_reg[1]_2 (fch_n_223),
        .\stat_reg[1]_3 (fch_n_249),
        .\stat_reg[1]_4 (fch_n_257),
        .\stat_reg[1]_5 ({bcmd[0],bcmd[2],badr[0]}),
        .\stat_reg[1]_6 (fch_n_284),
        .\stat_reg[1]_7 (fch_n_303),
        .\stat_reg[1]_8 (ctl0_n_7),
        .\stat_reg[2] (ctl_selc0_rn),
        .\stat_reg[2]_0 ({ctl_selc0,fch_n_83}),
        .\stat_reg[2]_1 ({fch_n_84,fch_n_85,ctl_selc1_rn}),
        .\stat_reg[2]_10 (fch_n_204),
        .\stat_reg[2]_11 (fch_n_242),
        .\stat_reg[2]_12 (stat_nx),
        .\stat_reg[2]_13 (fch_n_305),
        .\stat_reg[2]_14 (fch_n_335),
        .\stat_reg[2]_15 (fch_n_336),
        .\stat_reg[2]_16 (fch_n_337),
        .\stat_reg[2]_17 (fch_n_360),
        .\stat_reg[2]_18 (fch_n_428),
        .\stat_reg[2]_19 (fch_n_443),
        .\stat_reg[2]_2 ({ctl_selc1,fch_n_88}),
        .\stat_reg[2]_20 (fch_n_444),
        .\stat_reg[2]_21 (ctl0_n_18),
        .\stat_reg[2]_3 (fch_n_105),
        .\stat_reg[2]_4 (fch_n_169),
        .\stat_reg[2]_5 (bcmd[1]),
        .\stat_reg[2]_6 (fch_n_189),
        .\stat_reg[2]_7 (fch_n_190),
        .\stat_reg[2]_8 (fch_n_193),
        .\stat_reg[2]_9 (fch_n_201),
        .tout__1_carry__0(rgf_n_221),
        .tout__1_carry__0_i_1_0({fch_n_589,fch_n_590,fch_n_591,fch_n_592}),
        .tout__1_carry__0_i_3__0_0({fch_n_603,fch_n_604}),
        .tout__1_carry__1_i_1_0({fch_n_597,fch_n_598,fch_n_599,fch_n_600}),
        .tout__1_carry_i_11_0(fch_n_106),
        .tout__1_carry_i_1_0({fch_n_581,fch_n_582,fch_n_583,fch_n_584}),
        .tout__1_carry_i_1__0_0({fch_n_532,fch_n_533,fch_n_534,fch_n_535}),
        .tout__1_carry_i_22_0(ctl1_n_11),
        .tout__1_carry_i_25_0(ctl1_n_14),
        .\tr_reg[0] (fch_n_196),
        .\tr_reg[0]_0 (fch_n_202),
        .\tr_reg[0]_1 (fch_n_236),
        .\tr_reg[10] (fch_n_459),
        .\tr_reg[11] (fch_n_460),
        .\tr_reg[12] (fch_n_461),
        .\tr_reg[13] (fch_n_462),
        .\tr_reg[14] (fch_n_463),
        .\tr_reg[15] (fch_n_464),
        .\tr_reg[15]_0 (\treg/p_1_in ),
        .\tr_reg[15]_1 (rgf_tr),
        .\tr_reg[1] (fch_n_450),
        .\tr_reg[2] (fch_n_451),
        .\tr_reg[3] (fch_n_452),
        .\tr_reg[4] (fch_n_107),
        .\tr_reg[4]_0 (fch_n_186),
        .\tr_reg[4]_1 (fch_n_453),
        .\tr_reg[5] (fch_n_454),
        .\tr_reg[6] (fch_n_455),
        .\tr_reg[7] (fch_n_456),
        .\tr_reg[8] (fch_n_457),
        .\tr_reg[9] (fch_n_458));
  mcss_mem mem
       (.D(\bctl/ctl/stat_nx ),
        .O(alu1_n_1),
        .Q(\bctl/ctl/p_0_in ),
        .SR(\treg/p_0_in ),
        .bdatr(bdatr),
        .bdatr_15_sp_1(mem_n_23),
        .bdatr_2_sp_1(mem_n_8),
        .bdatr_6_sp_1(mem_n_10),
        .brdy(brdy),
        .brdy_0(mem_n_15),
        .brdy_1(mem_n_37),
        .brdy_2(mem_n_38),
        .cbus_i({cbus_i[15:14],cbus_i[11:10],cbus_i[8],cbus_i[3],cbus_i[0]}),
        .\cbus_i[15] (mem_n_7),
        .cbus_i_0_sp_1(mem_n_0),
        .cbus_i_3_sp_1(mem_n_2),
        .clk(clk),
        .fch_irq_req_fl(fch_irq_req_fl),
        .fch_memacc1(fch_memacc1),
        .fdat(fdat[15:2]),
        .\fdat[8] (lir_id_0),
        .fdatx(fdatx),
        .\fdatx[8]_0 (mem_n_20),
        .fdatx_8_sp_1(mem_n_19),
        .ir0_id(ir0_id),
        .\ir0_id_fl[21]_i_5 (fch_n_299),
        .\nir_id[21]_i_2 (fch_n_301),
        .\nir_id_reg[21] (fch_n_300),
        .out(fch_term),
        .\read_cyc_reg[0] (mem_n_24),
        .\read_cyc_reg[0]_0 (mem_n_26),
        .\read_cyc_reg[0]_1 (mem_n_30),
        .\read_cyc_reg[0]_2 (mem_n_32),
        .\read_cyc_reg[0]_3 (mem_n_36),
        .\read_cyc_reg[1] (mem_n_25),
        .\read_cyc_reg[1]_0 (mem_n_27),
        .\read_cyc_reg[1]_1 (mem_n_28),
        .\read_cyc_reg[1]_2 (mem_n_29),
        .\read_cyc_reg[2] (mem_n_9),
        .\read_cyc_reg[2]_0 (mem_n_11),
        .\read_cyc_reg[2]_1 (mem_n_12),
        .\read_cyc_reg[2]_2 (mem_n_13),
        .\read_cyc_reg[2]_3 (mem_n_14),
        .\read_cyc_reg[2]_4 ({bcmd[0],bcmd[2],badr[0]}),
        .\read_cyc_reg[3] (mem_n_1),
        .\read_cyc_reg[3]_0 (mem_n_3),
        .\read_cyc_reg[3]_1 (mem_n_4),
        .\read_cyc_reg[3]_2 (mem_n_5),
        .\read_cyc_reg[3]_3 (mem_n_6),
        .\read_cyc_reg[3]_4 (mem_n_31),
        .\read_cyc_reg[3]_5 (mem_n_33),
        .\read_cyc_reg[3]_6 (mem_n_34),
        .\read_cyc_reg[3]_7 (mem_n_35),
        .\rgf_c0bus_wb_reg[15] (fch_n_221),
        .\rgf_c1bus_wb_reg[14] (fch_n_106),
        .\rgf_c1bus_wb_reg[14]_0 ({alu1_n_13,alu1_n_14}),
        .\rgf_c1bus_wb_reg[6] (alu1_n_5),
        .\rgf_c1bus_wb_reg[9] ({alu1_n_10,alu1_n_11}),
        .\stat[0]_i_24__0 ({fch_ir1[5],fch_ir1[0]}),
        .\stat[0]_i_4 (fch_ir0[14:13]),
        .\stat[2]_i_7__0 (fch_n_445),
        .\stat_reg[1] (mem_n_18),
        .\stat_reg[1]_0 (mem_n_22));
  mcss_rgf rgf
       (.D(fch_pc),
        .E(fch_n_429),
        .O({fch_n_37,fch_n_38,fch_n_39}),
        .Q(stat_2[0]),
        .S(rgf_n_483),
        .SR(\treg/p_0_in ),
        .a0bus_0(a0bus_0),
        .a0bus_sel_0({a0bus_sel_0[7],a0bus_sel_0[4:3],a0bus_sel_0[0]}),
        .a0bus_sel_cr({a0bus_sel_cr[5],a0bus_sel_cr[2:0]}),
        .a1bus_0(a1bus_0),
        .a1bus_sel_0(a1bus_sel_0),
        .a1bus_sel_cr(a1bus_sel_cr),
        .a1bus_sr(a1bus_sr),
        .\abus_o[0] (fch_n_236),
        .\abus_o[10] (fch_n_459),
        .\abus_o[11] (fch_n_460),
        .\abus_o[12] (fch_n_461),
        .\abus_o[13] (fch_n_462),
        .\abus_o[14] (fch_n_463),
        .\abus_o[15] (fch_n_464),
        .\abus_o[1] (fch_n_450),
        .\abus_o[2] (fch_n_451),
        .\abus_o[3] (fch_n_452),
        .\abus_o[4] (fch_n_453),
        .\abus_o[5] (fch_n_454),
        .\abus_o[6] (fch_n_455),
        .\abus_o[7] (fch_n_456),
        .\abus_o[8] (fch_n_457),
        .\abus_o[9] (fch_n_458),
        .b0bus_sel_0(b0bus_sel_0),
        .b0bus_sel_cr(b0bus_sel_cr),
        .b0bus_sr(b0bus_sr),
        .b1bus_b02(b1bus_b02),
        .b1bus_sel_cr(b1bus_sel_cr),
        .b1bus_sr(b1bus_sr),
        .\badr[0]_INST_0_i_1 (rgf_n_268),
        .\badr[10]_INST_0_i_1 (rgf_n_240),
        .\badr[10]_INST_0_i_1_0 (rgf_n_244),
        .\badr[10]_INST_0_i_1_1 (rgf_n_272),
        .\badr[10]_INST_0_i_1_2 ({rgf_n_516,rgf_n_517,rgf_n_518,rgf_n_519}),
        .\badr[10]_INST_0_i_2 (rgf_n_378),
        .\badr[10]_INST_0_i_2_0 (rgf_n_387),
        .\badr[11]_INST_0_i_1 (rgf_n_284),
        .\badr[11]_INST_0_i_2 (rgf_n_419),
        .\badr[12]_INST_0_i_1 (rgf_n_265),
        .\badr[12]_INST_0_i_2 (rgf_n_391),
        .\badr[12]_INST_0_i_2_0 (rgf_n_444),
        .\badr[13]_INST_0_i_1 (rgf_n_293),
        .\badr[13]_INST_0_i_1_0 ({rgf_n_508,rgf_n_509,rgf_n_510}),
        .\badr[13]_INST_0_i_2 (rgf_n_371),
        .\badr[13]_INST_0_i_2_0 (rgf_n_402),
        .\badr[14]_INST_0_i_1 (rgf_n_245),
        .\badr[14]_INST_0_i_1_0 (rgf_n_298),
        .\badr[14]_INST_0_i_1_1 ({rgf_n_504,rgf_n_505,rgf_n_506,rgf_n_507}),
        .\badr[14]_INST_0_i_2 (rgf_n_388),
        .\badr[14]_INST_0_i_2_0 (rgf_n_397),
        .\badr[14]_INST_0_i_2_1 (rgf_n_436),
        .\badr[14]_INST_0_i_2_2 (rgf_n_511),
        .\badr[15]_INST_0_i_1 (rgf_n_227),
        .\badr[15]_INST_0_i_1_0 (rgf_n_234),
        .\badr[15]_INST_0_i_1_1 (rgf_n_249),
        .\badr[15]_INST_0_i_1_2 (rgf_n_255),
        .\badr[15]_INST_0_i_2 (rgf_n_446),
        .\badr[15]_INST_0_i_208 (fch_ir0[15:11]),
        .\badr[1]_INST_0_i_1 (rgf_n_235),
        .\badr[1]_INST_0_i_2 (rgf_n_370),
        .\badr[1]_INST_0_i_2_0 (rgf_n_433),
        .\badr[2]_INST_0_i_1 (rgf_n_242),
        .\badr[2]_INST_0_i_1_0 (rgf_n_287),
        .\badr[2]_INST_0_i_1_1 (rgf_n_294),
        .\badr[2]_INST_0_i_2 (rgf_n_380),
        .\badr[2]_INST_0_i_2_0 (rgf_n_424),
        .\badr[3]_INST_0_i_1 (rgf_n_230),
        .\badr[3]_INST_0_i_1_0 (rgf_n_247),
        .\badr[3]_INST_0_i_2 (rgf_n_376),
        .\badr[3]_INST_0_i_2_0 (rgf_n_415),
        .\badr[4]_INST_0_i_2 (rgf_n_383),
        .\badr[4]_INST_0_i_2_0 (rgf_n_390),
        .\badr[5]_INST_0_i_1 (rgf_n_222),
        .\badr[5]_INST_0_i_1_0 (rgf_n_260),
        .\badr[5]_INST_0_i_2 (rgf_n_369),
        .\badr[5]_INST_0_i_2_0 (rgf_n_403),
        .\badr[6]_INST_0_i_1 (rgf_n_218),
        .\badr[6]_INST_0_i_1_0 (rgf_n_241),
        .\badr[6]_INST_0_i_1_1 (rgf_n_251),
        .\badr[6]_INST_0_i_1_2 (rgf_n_303),
        .\badr[6]_INST_0_i_1_3 ({rgf_n_512,rgf_n_513}),
        .\badr[6]_INST_0_i_2 (rgf_n_358),
        .\badr[6]_INST_0_i_2_0 (rgf_n_379),
        .\badr[6]_INST_0_i_2_1 (rgf_n_400),
        .\badr[7]_INST_0_i_1 (rgf_n_248),
        .\badr[7]_INST_0_i_2 (rgf_n_420),
        .\badr[8]_INST_0_i_2 (rgf_n_375),
        .\badr[8]_INST_0_i_2_0 (rgf_n_392),
        .\badr[8]_INST_0_i_2_1 (rgf_n_443),
        .\badr[9]_INST_0_i_1 (rgf_n_237),
        .\badr[9]_INST_0_i_1_0 (rgf_n_290),
        .\badr[9]_INST_0_i_2 (rgf_n_372),
        .\badr[9]_INST_0_i_2_0 (rgf_n_404),
        .badrx(badrx),
        .badrx_15_sp_1(fch_n_257),
        .bbus_o(bbus_o[5]),
        .\bbus_o[0]_INST_0_i_7 (fch_n_381),
        .\bbus_o[0]_INST_0_i_7_0 (fch_n_396),
        .\bbus_o[0]_INST_0_i_7_1 (fch_n_386),
        .\bbus_o[0]_INST_0_i_7_2 (fch_n_391),
        .\bbus_o[0]_INST_0_i_7_3 (fch_n_376),
        .\bbus_o[0]_INST_0_i_7_4 (fch_n_371),
        .\bbus_o[0]_INST_0_i_7_5 (fch_n_365),
        .\bbus_o[0]_INST_0_i_7_6 (fch_n_358),
        .\bbus_o[1]_INST_0_i_7 (fch_n_380),
        .\bbus_o[1]_INST_0_i_7_0 (fch_n_395),
        .\bbus_o[1]_INST_0_i_7_1 (fch_n_385),
        .\bbus_o[1]_INST_0_i_7_2 (fch_n_390),
        .\bbus_o[1]_INST_0_i_7_3 (fch_n_375),
        .\bbus_o[1]_INST_0_i_7_4 (fch_n_370),
        .\bbus_o[1]_INST_0_i_7_5 (fch_n_364),
        .\bbus_o[1]_INST_0_i_7_6 (fch_n_357),
        .\bbus_o[2]_INST_0_i_7 (fch_n_379),
        .\bbus_o[2]_INST_0_i_7_0 (fch_n_394),
        .\bbus_o[2]_INST_0_i_7_1 (fch_n_384),
        .\bbus_o[2]_INST_0_i_7_2 (fch_n_389),
        .\bbus_o[2]_INST_0_i_7_3 (fch_n_374),
        .\bbus_o[2]_INST_0_i_7_4 (fch_n_369),
        .\bbus_o[2]_INST_0_i_7_5 (fch_n_363),
        .\bbus_o[2]_INST_0_i_7_6 (fch_n_356),
        .\bbus_o[3]_INST_0_i_7 (fch_n_378),
        .\bbus_o[3]_INST_0_i_7_0 (fch_n_393),
        .\bbus_o[3]_INST_0_i_7_1 (fch_n_383),
        .\bbus_o[3]_INST_0_i_7_2 (fch_n_388),
        .\bbus_o[3]_INST_0_i_7_3 (fch_n_373),
        .\bbus_o[3]_INST_0_i_7_4 (fch_n_368),
        .\bbus_o[3]_INST_0_i_7_5 (fch_n_362),
        .\bbus_o[3]_INST_0_i_7_6 (fch_n_355),
        .\bbus_o[4]_INST_0_i_7 (fch_n_377),
        .\bbus_o[4]_INST_0_i_7_0 (fch_n_392),
        .\bbus_o[4]_INST_0_i_7_1 (fch_n_382),
        .\bbus_o[4]_INST_0_i_7_2 (fch_n_387),
        .\bbus_o[4]_INST_0_i_7_3 (fch_n_372),
        .\bbus_o[4]_INST_0_i_7_4 (fch_n_366),
        .\bbus_o[4]_INST_0_i_7_5 (fch_n_359),
        .\bbus_o[4]_INST_0_i_7_6 (fch_n_353),
        .\bbus_o[5] (fch_n_436),
        .\bbus_o[5]_0 (fch_n_506),
        .\bbus_o[5]_1 (fch_n_221),
        .\bbus_o[6] (fch_n_435),
        .\bbus_o[6]_0 (fch_n_507),
        .\bbus_o[7] (fch_n_256),
        .\bbus_o[7]_0 (fch_n_508),
        .bdatw(bdatw[14:13]),
        .\bdatw[10] (fch_n_264),
        .\bdatw[10]_0 (fch_n_277),
        .\bdatw[10]_1 (fch_n_250),
        .\bdatw[10]_2 (fch_n_511),
        .\bdatw[10]_INST_0_i_43 (fch_n_325),
        .\bdatw[10]_INST_0_i_43_0 (fch_n_331),
        .\bdatw[11] (fch_n_268),
        .\bdatw[11]_0 (fch_n_276),
        .\bdatw[11]_1 (fch_n_434),
        .\bdatw[11]_2 (fch_n_512),
        .\bdatw[11]_INST_0_i_44 (fch_n_324),
        .\bdatw[11]_INST_0_i_44_0 (fch_n_330),
        .\bdatw[12] (fch_n_271),
        .\bdatw[12]_0 (fch_n_275),
        .\bdatw[12]_1 (fch_n_433),
        .\bdatw[12]_2 (fch_n_513),
        .\bdatw[12]_INST_0_i_42 (fch_n_322),
        .\bdatw[12]_INST_0_i_42_0 (fch_n_328),
        .\bdatw[13] (mem_n_18),
        .\bdatw[13]_0 (fch_n_184),
        .\bdatw[13]_1 (fch_n_185),
        .\bdatw[13]_2 (fch_n_269),
        .\bdatw[13]_3 (fch_n_274),
        .\bdatw[13]_4 (fch_n_432),
        .\bdatw[13]_5 (fch_n_514),
        .\bdatw[14] (fch_n_270),
        .\bdatw[14]_0 (fch_n_273),
        .\bdatw[14]_1 (fch_n_431),
        .\bdatw[14]_2 (fch_n_515),
        .\bdatw[15] (fch_n_430),
        .\bdatw[15]_0 (fch_n_516),
        .\bdatw[8] (fch_n_442),
        .\bdatw[8]_0 (fch_n_279),
        .\bdatw[8]_1 (fch_n_255),
        .\bdatw[8]_2 (fch_n_509),
        .\bdatw[8]_INST_0_i_43 (fch_n_327),
        .\bdatw[8]_INST_0_i_43_0 (fch_n_333),
        .\bdatw[9] (fch_n_272),
        .\bdatw[9]_0 (fch_n_278),
        .\bdatw[9]_1 (fch_n_254),
        .\bdatw[9]_2 (fch_n_510),
        .\bdatw[9]_INST_0_i_42 (fch_n_326),
        .\bdatw[9]_INST_0_i_42_0 (fch_n_332),
        .clk(clk),
        .ctl_fetch1_fl_i_15(fch_n_283),
        .ctl_sela0(ctl_sela0),
        .ctl_sela0_rn({ctl_sela0_rn[2],ctl_sela0_rn[0]}),
        .ctl_selb0_0(ctl_selb0_0),
        .ctl_selb0_rn(ctl_selb0_rn),
        .ctl_selb1_0(ctl_selb1_0),
        .ctl_selb1_rn(ctl_selb1_rn),
        .fadr(fadr[15:13]),
        .\fadr[15] (fch_n_248),
        .\fadr[15]_0 (fch_n_249),
        .fch_irq_req(fch_irq_req),
        .fdat({fdat[15:6],fdat[3:0]}),
        .\fdat[15] (rgf_n_502),
        .fdat_12_sp_1(rgf_n_482),
        .fdatx({fdatx[15:6],fdatx[3:0]}),
        .\fdatx[15] (rgf_n_481),
        .\grn_reg[0] (\bank02/p_1_in ),
        .\grn_reg[0]_0 (\bank02/p_0_in ),
        .\grn_reg[15] ({rgf_n_17,rgf_n_18,rgf_n_19,rgf_n_20,rgf_n_21,rgf_n_22,rgf_n_23,rgf_n_24,rgf_n_25,rgf_n_26,rgf_n_27,rgf_n_28,rgf_n_29,rgf_n_30,rgf_n_31,rgf_n_32}),
        .\grn_reg[15]_0 ({rgf_n_58,rgf_n_59,rgf_n_60,rgf_n_61,rgf_n_62,rgf_n_63,rgf_n_64,rgf_n_65,rgf_n_66,rgf_n_67,rgf_n_68,rgf_n_69,rgf_n_70,rgf_n_71,rgf_n_72,rgf_n_73}),
        .\grn_reg[15]_1 (a1bus_b02),
        .\grn_reg[15]_10 (fch_n_504),
        .\grn_reg[15]_11 ({fch_n_751,fch_n_752,fch_n_753,fch_n_754,fch_n_755,fch_n_756,fch_n_757,fch_n_758,fch_n_759,fch_n_760,fch_n_761,fch_n_762,fch_n_763,fch_n_764,fch_n_765,fch_n_766}),
        .\grn_reg[15]_12 (fch_n_1199),
        .\grn_reg[15]_13 ({fch_n_767,fch_n_768,fch_n_769,fch_n_770,fch_n_771,fch_n_772,fch_n_773,fch_n_774,fch_n_775,fch_n_776,fch_n_777,fch_n_778,fch_n_779,fch_n_780,fch_n_781,fch_n_782}),
        .\grn_reg[15]_14 (fch_n_500),
        .\grn_reg[15]_15 ({fch_n_783,fch_n_784,fch_n_785,fch_n_786,fch_n_787,fch_n_788,fch_n_789,fch_n_790,fch_n_791,fch_n_792,fch_n_793,fch_n_794,fch_n_795,fch_n_796,fch_n_797,fch_n_798}),
        .\grn_reg[15]_16 (fch_n_484),
        .\grn_reg[15]_17 ({fch_n_799,fch_n_800,fch_n_801,fch_n_802,fch_n_803,fch_n_804,fch_n_805,fch_n_806,fch_n_807,fch_n_808,fch_n_809,fch_n_810,fch_n_811,fch_n_812,fch_n_813,fch_n_814}),
        .\grn_reg[15]_18 (fch_n_575),
        .\grn_reg[15]_19 ({fch_n_815,fch_n_816,fch_n_817,fch_n_818,fch_n_819,fch_n_820,fch_n_821,fch_n_822,fch_n_823,fch_n_824,fch_n_825,fch_n_826,fch_n_827,fch_n_828,fch_n_829,fch_n_830}),
        .\grn_reg[15]_2 (fch_n_577),
        .\grn_reg[15]_20 (fch_n_493),
        .\grn_reg[15]_21 ({fch_n_831,fch_n_832,fch_n_833,fch_n_834,fch_n_835,fch_n_836,fch_n_837,fch_n_838,fch_n_839,fch_n_840,fch_n_841,fch_n_842,fch_n_843,fch_n_844,fch_n_845,fch_n_846}),
        .\grn_reg[15]_22 (fch_n_489),
        .\grn_reg[15]_23 ({fch_n_847,fch_n_848,fch_n_849,fch_n_850,fch_n_851,fch_n_852,fch_n_853,fch_n_854,fch_n_855,fch_n_856,fch_n_857,fch_n_858,fch_n_859,fch_n_860,fch_n_861,fch_n_862}),
        .\grn_reg[15]_24 (fch_n_485),
        .\grn_reg[15]_25 ({fch_n_863,fch_n_864,fch_n_865,fch_n_866,fch_n_867,fch_n_868,fch_n_869,fch_n_870,fch_n_871,fch_n_872,fch_n_873,fch_n_874,fch_n_875,fch_n_876,fch_n_877,fch_n_878}),
        .\grn_reg[15]_26 (fch_n_501),
        .\grn_reg[15]_27 ({fch_n_879,fch_n_880,fch_n_881,fch_n_882,fch_n_883,fch_n_884,fch_n_885,fch_n_886,fch_n_887,fch_n_888,fch_n_889,fch_n_890,fch_n_891,fch_n_892,fch_n_893,fch_n_894}),
        .\grn_reg[15]_28 (fch_n_1202),
        .\grn_reg[15]_29 ({fch_n_895,fch_n_896,fch_n_897,fch_n_898,fch_n_899,fch_n_900,fch_n_901,fch_n_902,fch_n_903,fch_n_904,fch_n_905,fch_n_906,fch_n_907,fch_n_908,fch_n_909,fch_n_910}),
        .\grn_reg[15]_3 (p_2_in),
        .\grn_reg[15]_30 (fch_n_497),
        .\grn_reg[15]_31 ({fch_n_911,fch_n_912,fch_n_913,fch_n_914,fch_n_915,fch_n_916,fch_n_917,fch_n_918,fch_n_919,fch_n_920,fch_n_921,fch_n_922,fch_n_923,fch_n_924,fch_n_925,fch_n_926}),
        .\grn_reg[15]_32 (fch_n_481),
        .\grn_reg[15]_33 ({fch_n_927,fch_n_928,fch_n_929,fch_n_930,fch_n_931,fch_n_932,fch_n_933,fch_n_934,fch_n_935,fch_n_936,fch_n_937,fch_n_938,fch_n_939,fch_n_940,fch_n_941,fch_n_942}),
        .\grn_reg[15]_34 (fch_n_574),
        .\grn_reg[15]_35 ({fch_n_943,fch_n_944,fch_n_945,fch_n_946,fch_n_947,fch_n_948,fch_n_949,fch_n_950,fch_n_951,fch_n_952,fch_n_953,fch_n_954,fch_n_955,fch_n_956,fch_n_957,fch_n_958}),
        .\grn_reg[15]_36 (fch_n_494),
        .\grn_reg[15]_37 ({fch_n_959,fch_n_960,fch_n_961,fch_n_962,fch_n_963,fch_n_964,fch_n_965,fch_n_966,fch_n_967,fch_n_968,fch_n_969,fch_n_970,fch_n_971,fch_n_972,fch_n_973,fch_n_974}),
        .\grn_reg[15]_38 (fch_n_490),
        .\grn_reg[15]_39 ({fch_n_975,fch_n_976,fch_n_977,fch_n_978,fch_n_979,fch_n_980,fch_n_981,fch_n_982,fch_n_983,fch_n_984,fch_n_985,fch_n_986,fch_n_987,fch_n_988,fch_n_989,fch_n_990}),
        .\grn_reg[15]_4 (fch_n_496),
        .\grn_reg[15]_40 (fch_n_486),
        .\grn_reg[15]_41 ({fch_n_991,fch_n_992,fch_n_993,fch_n_994,fch_n_995,fch_n_996,fch_n_997,fch_n_998,fch_n_999,fch_n_1000,fch_n_1001,fch_n_1002,fch_n_1003,fch_n_1004,fch_n_1005,fch_n_1006}),
        .\grn_reg[15]_42 (fch_n_502),
        .\grn_reg[15]_43 ({fch_n_1007,fch_n_1008,fch_n_1009,fch_n_1010,fch_n_1011,fch_n_1012,fch_n_1013,fch_n_1014,fch_n_1015,fch_n_1016,fch_n_1017,fch_n_1018,fch_n_1019,fch_n_1020,fch_n_1021,fch_n_1022}),
        .\grn_reg[15]_44 (fch_n_1201),
        .\grn_reg[15]_45 ({fch_n_1023,fch_n_1024,fch_n_1025,fch_n_1026,fch_n_1027,fch_n_1028,fch_n_1029,fch_n_1030,fch_n_1031,fch_n_1032,fch_n_1033,fch_n_1034,fch_n_1035,fch_n_1036,fch_n_1037,fch_n_1038}),
        .\grn_reg[15]_46 (fch_n_498),
        .\grn_reg[15]_47 ({fch_n_1039,fch_n_1040,fch_n_1041,fch_n_1042,fch_n_1043,fch_n_1044,fch_n_1045,fch_n_1046,fch_n_1047,fch_n_1048,fch_n_1049,fch_n_1050,fch_n_1051,fch_n_1052,fch_n_1053,fch_n_1054}),
        .\grn_reg[15]_48 (fch_n_482),
        .\grn_reg[15]_49 ({fch_n_1055,fch_n_1056,fch_n_1057,fch_n_1058,fch_n_1059,fch_n_1060,fch_n_1061,fch_n_1062,fch_n_1063,fch_n_1064,fch_n_1065,fch_n_1066,fch_n_1067,fch_n_1068,fch_n_1069,fch_n_1070}),
        .\grn_reg[15]_5 ({fch_n_703,fch_n_704,fch_n_705,fch_n_706,fch_n_707,fch_n_708,fch_n_709,fch_n_710,fch_n_711,fch_n_712,fch_n_713,fch_n_714,fch_n_715,fch_n_716,fch_n_717,fch_n_718}),
        .\grn_reg[15]_50 (fch_n_576),
        .\grn_reg[15]_51 ({fch_n_1071,fch_n_1072,fch_n_1073,fch_n_1074,fch_n_1075,fch_n_1076,fch_n_1077,fch_n_1078,fch_n_1079,fch_n_1080,fch_n_1081,fch_n_1082,fch_n_1083,fch_n_1084,fch_n_1085,fch_n_1086}),
        .\grn_reg[15]_52 (fch_n_495),
        .\grn_reg[15]_53 ({fch_n_1087,fch_n_1088,fch_n_1089,fch_n_1090,fch_n_1091,fch_n_1092,fch_n_1093,fch_n_1094,fch_n_1095,fch_n_1096,fch_n_1097,fch_n_1098,fch_n_1099,fch_n_1100,fch_n_1101,fch_n_1102}),
        .\grn_reg[15]_54 (fch_n_491),
        .\grn_reg[15]_55 ({fch_n_1103,fch_n_1104,fch_n_1105,fch_n_1106,fch_n_1107,fch_n_1108,fch_n_1109,fch_n_1110,fch_n_1111,fch_n_1112,fch_n_1113,fch_n_1114,fch_n_1115,fch_n_1116,fch_n_1117,fch_n_1118}),
        .\grn_reg[15]_56 (fch_n_487),
        .\grn_reg[15]_57 ({fch_n_1119,fch_n_1120,fch_n_1121,fch_n_1122,fch_n_1123,fch_n_1124,fch_n_1125,fch_n_1126,fch_n_1127,fch_n_1128,fch_n_1129,fch_n_1130,fch_n_1131,fch_n_1132,fch_n_1133,fch_n_1134}),
        .\grn_reg[15]_58 (fch_n_503),
        .\grn_reg[15]_59 ({fch_n_1135,fch_n_1136,fch_n_1137,fch_n_1138,fch_n_1139,fch_n_1140,fch_n_1141,fch_n_1142,fch_n_1143,fch_n_1144,fch_n_1145,fch_n_1146,fch_n_1147,fch_n_1148,fch_n_1149,fch_n_1150}),
        .\grn_reg[15]_6 (fch_n_492),
        .\grn_reg[15]_60 (fch_n_1200),
        .\grn_reg[15]_61 ({fch_n_1151,fch_n_1152,fch_n_1153,fch_n_1154,fch_n_1155,fch_n_1156,fch_n_1157,fch_n_1158,fch_n_1159,fch_n_1160,fch_n_1161,fch_n_1162,fch_n_1163,fch_n_1164,fch_n_1165,fch_n_1166}),
        .\grn_reg[15]_62 (fch_n_499),
        .\grn_reg[15]_63 ({fch_n_1167,fch_n_1168,fch_n_1169,fch_n_1170,fch_n_1171,fch_n_1172,fch_n_1173,fch_n_1174,fch_n_1175,fch_n_1176,fch_n_1177,fch_n_1178,fch_n_1179,fch_n_1180,fch_n_1181,fch_n_1182}),
        .\grn_reg[15]_64 (fch_n_483),
        .\grn_reg[15]_65 ({fch_n_1183,fch_n_1184,fch_n_1185,fch_n_1186,fch_n_1187,fch_n_1188,fch_n_1189,fch_n_1190,fch_n_1191,fch_n_1192,fch_n_1193,fch_n_1194,fch_n_1195,fch_n_1196,fch_n_1197,fch_n_1198}),
        .\grn_reg[15]_7 ({fch_n_719,fch_n_720,fch_n_721,fch_n_722,fch_n_723,fch_n_724,fch_n_725,fch_n_726,fch_n_727,fch_n_728,fch_n_729,fch_n_730,fch_n_731,fch_n_732,fch_n_733,fch_n_734}),
        .\grn_reg[15]_8 (fch_n_488),
        .\grn_reg[15]_9 ({fch_n_735,fch_n_736,fch_n_737,fch_n_738,fch_n_739,fch_n_740,fch_n_741,fch_n_742,fch_n_743,fch_n_744,fch_n_745,fch_n_746,fch_n_747,fch_n_748,fch_n_749,fch_n_750}),
        .\grn_reg[4] ({rgf_n_33,rgf_n_34,rgf_n_35,rgf_n_36,rgf_n_37}),
        .\grn_reg[4]_0 ({rgf_n_38,rgf_n_39,rgf_n_40,rgf_n_41,rgf_n_42}),
        .\grn_reg[4]_1 ({rgf_n_43,rgf_n_44,rgf_n_45,rgf_n_46,rgf_n_47}),
        .\grn_reg[4]_2 ({rgf_n_48,rgf_n_49,rgf_n_50,rgf_n_51,rgf_n_52}),
        .\grn_reg[4]_3 ({rgf_n_53,rgf_n_54,rgf_n_55,rgf_n_56,rgf_n_57}),
        .\grn_reg[4]_4 ({rgf_n_74,rgf_n_75,rgf_n_76,rgf_n_77,rgf_n_78}),
        .\grn_reg[4]_5 ({rgf_n_79,rgf_n_80,rgf_n_81,rgf_n_82,rgf_n_83}),
        .\grn_reg[4]_6 ({rgf_n_84,rgf_n_85,rgf_n_86,rgf_n_87,rgf_n_88}),
        .\grn_reg[4]_7 ({rgf_n_89,rgf_n_90,rgf_n_91,rgf_n_92,rgf_n_93}),
        .\grn_reg[4]_8 (\bank02/p_1_in3_in ),
        .\grn_reg[4]_9 (\bank02/p_0_in2_in ),
        .\i_/badr[15]_INST_0_i_19 (fch_n_337),
        .\i_/badr[15]_INST_0_i_19_0 (fch_n_336),
        .\i_/badr[15]_INST_0_i_19_1 (fch_n_335),
        .\i_/badr[15]_INST_0_i_43 (fch_n_428),
        .\i_/badr[15]_INST_0_i_43_0 (fch_n_444),
        .\i_/bbus_o[4]_INST_0_i_20 (fch_n_438),
        .\i_/bbus_o[4]_INST_0_i_20_0 (fch_n_437),
        .\i_/bdatw[15]_INST_0_i_112 (fch_n_650),
        .\i_/bdatw[15]_INST_0_i_112_0 (fch_n_267),
        .\i_/bdatw[15]_INST_0_i_112_1 (fch_n_265),
        .\i_/bdatw[15]_INST_0_i_113 (fch_n_323),
        .\i_/bdatw[15]_INST_0_i_24 (fch_n_645),
        .\i_/bdatw[15]_INST_0_i_24_0 (fch_n_367),
        .\i_/bdatw[15]_INST_0_i_44 (fch_n_329),
        .\i_/bdatw[15]_INST_0_i_77 (fch_n_354),
        .\i_/bdatw[15]_INST_0_i_9 (fch_n_642),
        .\i_/bdatw[15]_INST_0_i_9_0 (fch_n_360),
        .\i_/bdatw[15]_INST_0_i_9_1 (fch_n_251),
        .\i_/bdatw[15]_INST_0_i_9_2 (fch_n_253),
        .\i_/bdatw[15]_INST_0_i_9_3 (fch_n_361),
        .\ir0_id_fl[20]_i_4 (fch_n_298),
        .irq(irq),
        .irq_0(rgf_n_478),
        .irq_lev(irq_lev),
        .\iv_reg[15] ({\ivec/p_0_in ,rgf_iv_ve}),
        .\iv_reg[15]_0 (rgf_n_579),
        .\iv_reg[15]_1 (\ivec/p_1_in ),
        .\nir_id_reg[20] (fch_n_302),
        .out({rgf_n_2,rgf_n_3,rgf_n_4,rgf_n_5,rgf_n_6,rgf_n_7,rgf_n_8,rgf_n_9,rgf_n_10,rgf_n_11,rgf_n_12,rgf_n_13,rgf_n_14,rgf_n_15,rgf_n_16}),
        .p_2_in(\rctl/p_2_in ),
        .\pc0_reg[15] (p_2_in_4),
        .\pc0_reg[15]_0 (fch_n_147),
        .\pc0_reg[15]_1 (fch_n_148),
        .\pc_reg[13] (rgf_n_166),
        .\pc_reg[13]_0 (fch_n_146),
        .\pc_reg[14] (rgf_n_165),
        .\pc_reg[15] (rgf_pc),
        .\pc_reg[15]_0 (rgf_n_161),
        .\pc_reg[15]_1 ({rgf_n_485,rgf_n_486,rgf_n_487}),
        .\pc_reg[15]_2 (\pcnt/p_1_in ),
        .\pc_reg[1] (rgf_n_484),
        .\rgf_c0bus_wb[0]_i_14 (rgf_n_384),
        .\rgf_c0bus_wb[10]_i_4 (fch_n_227),
        .\rgf_c0bus_wb[10]_i_8 (rgf_n_431),
        .\rgf_c0bus_wb[11]_i_11 (rgf_n_368),
        .\rgf_c0bus_wb[11]_i_11_0 (rgf_n_373),
        .\rgf_c0bus_wb[11]_i_11_1 (rgf_n_399),
        .\rgf_c0bus_wb[11]_i_11_2 (rgf_n_401),
        .\rgf_c0bus_wb[11]_i_22 (rgf_n_374),
        .\rgf_c0bus_wb[11]_i_22_0 (rgf_n_421),
        .\rgf_c0bus_wb[11]_i_3 (rgf_n_340),
        .\rgf_c0bus_wb[11]_i_3_0 (rgf_n_357),
        .\rgf_c0bus_wb[11]_i_3_1 (rgf_n_449),
        .\rgf_c0bus_wb[11]_i_3_2 (rgf_n_495),
        .\rgf_c0bus_wb[11]_i_3_3 (rgf_n_498),
        .\rgf_c0bus_wb[11]_i_8 (rgf_n_382),
        .\rgf_c0bus_wb[11]_i_9 (rgf_n_361),
        .\rgf_c0bus_wb[11]_i_9_0 (rgf_n_364),
        .\rgf_c0bus_wb[11]_i_9_1 (rgf_n_377),
        .\rgf_c0bus_wb[11]_i_9_2 (rgf_n_432),
        .\rgf_c0bus_wb[11]_i_9_3 (rgf_n_496),
        .\rgf_c0bus_wb[11]_i_9_4 (rgf_n_497),
        .\rgf_c0bus_wb[12]_i_2 (fch_n_234),
        .\rgf_c0bus_wb[12]_i_24 (rgf_n_426),
        .\rgf_c0bus_wb[12]_i_25 (rgf_n_438),
        .\rgf_c0bus_wb[13]_i_27 (rgf_n_366),
        .\rgf_c0bus_wb[13]_i_28 (rgf_n_434),
        .\rgf_c0bus_wb[13]_i_29 (rgf_n_389),
        .\rgf_c0bus_wb[13]_i_30 (rgf_n_408),
        .\rgf_c0bus_wb[13]_i_4 (fch_n_231),
        .\rgf_c0bus_wb[14]_i_2 (fch_n_204),
        .\rgf_c0bus_wb[15]_i_14 (fch_n_225),
        .\rgf_c0bus_wb[15]_i_18 (rgf_n_339),
        .\rgf_c0bus_wb[15]_i_25 (rgf_n_381),
        .\rgf_c0bus_wb[15]_i_26 (rgf_n_405),
        .\rgf_c0bus_wb[15]_i_6 (rgf_n_491),
        .\rgf_c0bus_wb[15]_i_6_0 (rgf_n_492),
        .\rgf_c0bus_wb[15]_i_6_1 (rgf_n_493),
        .\rgf_c0bus_wb[3]_i_7 (fch_n_232),
        .\rgf_c0bus_wb[3]_i_7_0 (fch_n_202),
        .\rgf_c0bus_wb[4]_i_21 (fch_pc0),
        .\rgf_c0bus_wb[4]_i_26 (rgf_n_360),
        .\rgf_c0bus_wb[4]_i_29 (rgf_n_414),
        .\rgf_c0bus_wb[4]_i_31 (rgf_n_418),
        .\rgf_c0bus_wb[4]_i_32 (rgf_n_365),
        .\rgf_c0bus_wb[4]_i_33 (rgf_n_417),
        .\rgf_c0bus_wb[6]_i_11 (fch_n_223),
        .\rgf_c0bus_wb[7]_i_7 (rgf_n_393),
        .\rgf_c0bus_wb[7]_i_7_0 (rgf_n_394),
        .\rgf_c0bus_wb[8]_i_6 (rgf_n_437),
        .\rgf_c0bus_wb_reg[10] (fch_n_224),
        .\rgf_c0bus_wb_reg[10]_0 (fch_n_228),
        .\rgf_c0bus_wb_reg[10]_1 (fch_n_226),
        .\rgf_c0bus_wb_reg[15] (\rctl/rgf_c0bus_wb ),
        .\rgf_c0bus_wb_reg[15]_0 (c0bus),
        .\rgf_c0bus_wb_reg[7]_i_11 (fch_n_203),
        .\rgf_c1bus_wb[11]_i_10 (rgf_n_254),
        .\rgf_c1bus_wb[11]_i_10_0 (rgf_n_263),
        .\rgf_c1bus_wb[11]_i_10_1 (rgf_n_301),
        .\rgf_c1bus_wb[11]_i_10_2 (rgf_n_304),
        .\rgf_c1bus_wb[11]_i_10_3 (rgf_n_311),
        .\rgf_c1bus_wb[11]_i_10_4 (rgf_n_312),
        .\rgf_c1bus_wb[11]_i_10_5 (rgf_n_490),
        .\rgf_c1bus_wb[11]_i_13 (rgf_n_243),
        .\rgf_c1bus_wb[12]_i_2 (fch_n_197),
        .\rgf_c1bus_wb[12]_i_20 (rgf_n_253),
        .\rgf_c1bus_wb[13]_i_16 (rgf_n_274),
        .\rgf_c1bus_wb[13]_i_9 (rgf_n_224),
        .\rgf_c1bus_wb[14]_i_11 (fch_n_440),
        .\rgf_c1bus_wb[14]_i_11_0 (fch_n_281),
        .\rgf_c1bus_wb[14]_i_28 (rgf_n_256),
        .\rgf_c1bus_wb[14]_i_28_0 (rgf_n_258),
        .\rgf_c1bus_wb[14]_i_28_1 (rgf_n_266),
        .\rgf_c1bus_wb[14]_i_28_2 (rgf_n_269),
        .\rgf_c1bus_wb[14]_i_28_3 (rgf_n_270),
        .\rgf_c1bus_wb[14]_i_28_4 (rgf_n_273),
        .\rgf_c1bus_wb[14]_i_28_5 (rgf_n_275),
        .\rgf_c1bus_wb[14]_i_28_6 (rgf_n_289),
        .\rgf_c1bus_wb[14]_i_28_7 (rgf_n_291),
        .\rgf_c1bus_wb[14]_i_30 (rgf_n_225),
        .\rgf_c1bus_wb[14]_i_32 (rgf_n_292),
        .\rgf_c1bus_wb[14]_i_32_0 (rgf_n_295),
        .\rgf_c1bus_wb[15]_i_14 (rgf_n_239),
        .\rgf_c1bus_wb[15]_i_14_0 (rgf_n_246),
        .\rgf_c1bus_wb[15]_i_14_1 (rgf_n_257),
        .\rgf_c1bus_wb[15]_i_14_2 (rgf_n_283),
        .\rgf_c1bus_wb[15]_i_14_3 (rgf_n_288),
        .\rgf_c1bus_wb[15]_i_19 (fch_n_441),
        .\rgf_c1bus_wb[15]_i_19_0 (fch_n_280),
        .\rgf_c1bus_wb[15]_i_27 (rgf_n_313),
        .\rgf_c1bus_wb[1]_i_14 (rgf_n_302),
        .\rgf_c1bus_wb[4]_i_22 (fch_pc1),
        .\rgf_c1bus_wb[4]_i_28 (rgf_n_307),
        .\rgf_c1bus_wb[4]_i_32 (fch_n_408),
        .\rgf_c1bus_wb[4]_i_32_0 (fch_n_348),
        .\rgf_c1bus_wb[4]_i_33 (fch_n_424),
        .\rgf_c1bus_wb[4]_i_34 (fch_n_409),
        .\rgf_c1bus_wb[4]_i_34_0 (fch_n_349),
        .\rgf_c1bus_wb[4]_i_36 (fch_n_410),
        .\rgf_c1bus_wb[4]_i_36_0 (fch_n_350),
        .\rgf_c1bus_wb[4]_i_37 (fch_n_426),
        .\rgf_c1bus_wb[4]_i_38 (fch_n_411),
        .\rgf_c1bus_wb[4]_i_38_0 (fch_n_351),
        .\rgf_c1bus_wb[4]_i_40 (fch_n_397),
        .\rgf_c1bus_wb[4]_i_41 (fch_n_414),
        .\rgf_c1bus_wb[4]_i_42 (fch_n_398),
        .\rgf_c1bus_wb[4]_i_42_0 (fch_n_338),
        .\rgf_c1bus_wb[4]_i_44 (fch_n_352),
        .\rgf_c1bus_wb[4]_i_45 (fch_n_334),
        .\rgf_c1bus_wb[4]_i_47 (fch_n_413),
        .\rgf_c1bus_wb[4]_i_48 (fch_n_400),
        .\rgf_c1bus_wb[4]_i_48_0 (fch_n_340),
        .\rgf_c1bus_wb[4]_i_50 (fch_n_399),
        .\rgf_c1bus_wb[4]_i_50_0 (fch_n_339),
        .\rgf_c1bus_wb[4]_i_51 (fch_n_415),
        .\rgf_c1bus_wb[4]_i_52 (fch_n_407),
        .\rgf_c1bus_wb[4]_i_52_0 (fch_n_347),
        .\rgf_c1bus_wb[4]_i_53 (fch_n_422),
        .\rgf_c1bus_wb[4]_i_54 (fch_n_406),
        .\rgf_c1bus_wb[4]_i_54_0 (fch_n_346),
        .\rgf_c1bus_wb[4]_i_56 (fch_n_405),
        .\rgf_c1bus_wb[4]_i_56_0 (fch_n_345),
        .\rgf_c1bus_wb[4]_i_57 (fch_n_420),
        .\rgf_c1bus_wb[4]_i_58 (fch_n_404),
        .\rgf_c1bus_wb[4]_i_58_0 (fch_n_344),
        .\rgf_c1bus_wb[4]_i_60 (fch_n_403),
        .\rgf_c1bus_wb[4]_i_60_0 (fch_n_343),
        .\rgf_c1bus_wb[4]_i_61 (fch_n_419),
        .\rgf_c1bus_wb[4]_i_62 (fch_n_402),
        .\rgf_c1bus_wb[4]_i_62_0 (fch_n_342),
        .\rgf_c1bus_wb[4]_i_64 (fch_n_401),
        .\rgf_c1bus_wb[4]_i_64_0 (fch_n_341),
        .\rgf_c1bus_wb[4]_i_65 (fch_n_417),
        .\rgf_c1bus_wb[4]_i_67 (fch_n_425),
        .\rgf_c1bus_wb[4]_i_9 (rgf_n_264),
        .\rgf_c1bus_wb[4]_i_9_0 (rgf_n_276),
        .\rgf_c1bus_wb[5]_i_10 (fch_n_189),
        .\rgf_c1bus_wb[7]_i_4 (rgf_n_259),
        .\rgf_c1bus_wb[7]_i_4_0 (rgf_n_488),
        .\rgf_c1bus_wb[9]_i_17 (rgf_n_271),
        .\rgf_c1bus_wb_reg[0] (fch_term),
        .\rgf_c1bus_wb_reg[10] (fch_n_186),
        .\rgf_c1bus_wb_reg[15] (\rctl/rgf_c1bus_wb ),
        .\rgf_c1bus_wb_reg[15]_0 (c1bus),
        .\rgf_c1bus_wb_reg[3] (fch_n_187),
        .\rgf_c1bus_wb_reg[4] (fch_n_193),
        .\rgf_c1bus_wb_reg[5] (fch_n_168),
        .\rgf_c1bus_wb_reg[5]_0 (fch_n_190),
        .\rgf_c1bus_wb_reg[5]_1 (fch_n_192),
        .\rgf_c1bus_wb_reg[7] (fch_n_191),
        .\rgf_selc0_rn_wb_reg[2] (\rctl/rgf_selc0_rn_wb ),
        .\rgf_selc0_rn_wb_reg[2]_0 (ctl_selc0_rn),
        .rgf_selc0_stat(\rctl/rgf_selc0_stat ),
        .\rgf_selc0_wb_reg[1] (\rctl/rgf_selc0_wb ),
        .\rgf_selc0_wb_reg[1]_0 ({ctl_selc0,fch_n_83}),
        .\rgf_selc1_rn_wb_reg[2] (\rctl/rgf_selc1_rn_wb ),
        .\rgf_selc1_rn_wb_reg[2]_0 ({fch_n_84,fch_n_85,ctl_selc1_rn}),
        .rgf_selc1_stat(\rctl/rgf_selc1_stat ),
        .rgf_selc1_stat_reg(fch_n_78),
        .\rgf_selc1_wb[1]_i_16 (fch_ir1[14:11]),
        .\rgf_selc1_wb_reg[0] (fch_n_443),
        .\rgf_selc1_wb_reg[1] (\rctl/rgf_selc1_wb ),
        .\rgf_selc1_wb_reg[1]_0 ({ctl_selc1,fch_n_88}),
        .rst_n(rst_n),
        .\sp_reg[0] (\sptr/p_0_in ),
        .\sp_reg[0]_0 (rgf_n_447),
        .\sp_reg[0]_1 (rgf_n_573),
        .\sp_reg[0]_2 (rgf_n_591),
        .\sp_reg[10] (rgf_n_179),
        .\sp_reg[11] (rgf_n_180),
        .\sp_reg[11]_0 (rgf_n_412),
        .\sp_reg[12] (rgf_n_181),
        .\sp_reg[13] (rgf_n_182),
        .\sp_reg[13]_0 (rgf_n_411),
        .\sp_reg[14] (rgf_n_183),
        .\sp_reg[14]_0 (fch_n_165),
        .\sp_reg[14]_1 (fch_n_166),
        .\sp_reg[15] (rgf_n_169),
        .\sp_reg[15]_0 (rgf_n_318),
        .\sp_reg[15]_1 ({fch_n_149,fch_n_150,fch_n_151,fch_n_152,fch_n_153,fch_n_154,fch_n_155,fch_n_156,fch_n_157,fch_n_158,fch_n_159,fch_n_160,fch_n_161,fch_n_162,fch_n_163,fch_n_164}),
        .\sp_reg[1] (\sptr/data3 ),
        .\sp_reg[1]_0 (rgf_n_170),
        .\sp_reg[1]_1 (rgf_n_423),
        .\sp_reg[1]_2 (rgf_n_572),
        .\sp_reg[1]_3 (rgf_n_592),
        .\sp_reg[2] (rgf_n_171),
        .\sp_reg[2]_0 (rgf_n_407),
        .\sp_reg[2]_1 (rgf_n_571),
        .\sp_reg[2]_2 (rgf_n_593),
        .\sp_reg[3] (rgf_n_172),
        .\sp_reg[3]_0 (rgf_n_570),
        .\sp_reg[3]_1 (rgf_n_594),
        .\sp_reg[4] (rgf_n_173),
        .\sp_reg[4]_0 (rgf_n_427),
        .\sp_reg[4]_1 (rgf_n_569),
        .\sp_reg[4]_2 (rgf_n_595),
        .\sp_reg[5] (rgf_n_174),
        .\sp_reg[6] (rgf_n_175),
        .\sp_reg[7] (rgf_n_176),
        .\sp_reg[8] (rgf_n_177),
        .\sp_reg[9] (rgf_n_178),
        .\sr[4]_i_129 (fch_n_235),
        .\sr[4]_i_133 (rgf_n_359),
        .\sr[4]_i_15 (fch_n_222),
        .\sr[4]_i_156 (rgf_n_231),
        .\sr[4]_i_15_0 (fch_n_107),
        .\sr[4]_i_15_1 (fch_n_229),
        .\sr[4]_i_195 (rgf_n_363),
        .\sr[4]_i_200 (rgf_n_362),
        .\sr[4]_i_219 (rgf_n_261),
        .\sr[4]_i_220 (rgf_n_309),
        .\sr[4]_i_232 (rgf_n_422),
        .\sr[4]_i_235 (fch_n_416),
        .\sr[4]_i_237 (fch_n_418),
        .\sr[4]_i_239 (fch_n_412),
        .\sr[4]_i_240 (fch_n_427),
        .\sr[4]_i_243 (fch_n_423),
        .\sr[4]_i_245 (fch_n_421),
        .\sr[4]_i_27 (fch_n_198),
        .\sr[4]_i_30 (fch_n_195),
        .\sr[4]_i_38 (fch_n_201),
        .\sr[4]_i_44 (fch_n_199),
        .\sr[4]_i_55 (fch_n_233),
        .\sr[4]_i_66 (fch_n_230),
        .\sr[4]_i_67 (fch_n_205),
        .\sr[4]_i_84 (fch_n_200),
        .\sr[6]_i_11 (fch_n_196),
        .\sr[6]_i_11_0 (fch_n_194),
        .\sr[6]_i_11_1 (fch_n_305),
        .\sr[6]_i_15 (fch_n_169),
        .\sr_reg[0] (rgf_n_448),
        .\sr_reg[0]_0 (rgf_n_503),
        .\sr_reg[0]_1 (bank_sel),
        .\sr_reg[0]_2 (rgf_n_585),
        .\sr_reg[10] (rgf_n_479),
        .\sr_reg[14] (rgf_n_428),
        .\sr_reg[15] ({\sreg/p_2_in [7:4],rgf_sr_ml,rgf_sr_dr,rgf_sr_sd,\sreg/p_2_in [0],rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[15]_0 (rgf_n_317),
        .\sr_reg[15]_1 (rgf_n_580),
        .\sr_reg[15]_2 (\sreg/p_0_in ),
        .\sr_reg[1] (rgf_n_584),
        .\sr_reg[2] (rgf_n_583),
        .\sr_reg[3] (rgf_n_582),
        .\sr_reg[4] (rgf_n_159),
        .\sr_reg[4]_0 (rgf_n_471),
        .\sr_reg[4]_1 (rgf_n_480),
        .\sr_reg[4]_2 (rgf_n_581),
        .\sr_reg[5] (rgf_n_160),
        .\sr_reg[5]_0 (rgf_n_472),
        .\sr_reg[5]_1 (rgf_n_474),
        .\sr_reg[5]_2 (rgf_n_476),
        .\sr_reg[5]_3 (rgf_n_499),
        .\sr_reg[5]_4 (rgf_n_500),
        .\sr_reg[5]_5 (rgf_n_501),
        .\sr_reg[5]_6 (fch_n_108),
        .\sr_reg[6] (rgf_n_226),
        .\sr_reg[6]_0 (rgf_n_228),
        .\sr_reg[6]_1 (rgf_n_229),
        .\sr_reg[6]_10 (rgf_n_282),
        .\sr_reg[6]_11 (rgf_n_285),
        .\sr_reg[6]_12 (rgf_n_286),
        .\sr_reg[6]_13 (rgf_n_296),
        .\sr_reg[6]_14 (rgf_n_297),
        .\sr_reg[6]_15 (rgf_n_300),
        .\sr_reg[6]_16 (rgf_n_305),
        .\sr_reg[6]_17 (rgf_n_306),
        .\sr_reg[6]_18 (rgf_n_314),
        .\sr_reg[6]_19 (rgf_n_367),
        .\sr_reg[6]_2 (rgf_n_236),
        .\sr_reg[6]_20 (rgf_n_385),
        .\sr_reg[6]_21 (rgf_n_386),
        .\sr_reg[6]_22 (rgf_n_395),
        .\sr_reg[6]_23 (rgf_n_396),
        .\sr_reg[6]_24 (rgf_n_398),
        .\sr_reg[6]_25 (rgf_n_406),
        .\sr_reg[6]_26 (rgf_n_409),
        .\sr_reg[6]_27 (rgf_n_410),
        .\sr_reg[6]_28 (rgf_n_413),
        .\sr_reg[6]_29 (rgf_n_416),
        .\sr_reg[6]_3 (rgf_n_238),
        .\sr_reg[6]_30 (rgf_n_425),
        .\sr_reg[6]_31 (rgf_n_429),
        .\sr_reg[6]_32 (rgf_n_430),
        .\sr_reg[6]_33 (rgf_n_435),
        .\sr_reg[6]_34 (rgf_n_439),
        .\sr_reg[6]_35 (rgf_n_440),
        .\sr_reg[6]_36 (rgf_n_441),
        .\sr_reg[6]_37 (rgf_n_442),
        .\sr_reg[6]_38 (rgf_n_445),
        .\sr_reg[6]_39 (rgf_n_450),
        .\sr_reg[6]_4 (rgf_n_250),
        .\sr_reg[6]_40 (rgf_n_475),
        .\sr_reg[6]_41 (rgf_n_477),
        .\sr_reg[6]_42 (rgf_n_489),
        .\sr_reg[6]_5 (rgf_n_252),
        .\sr_reg[6]_6 (rgf_n_267),
        .\sr_reg[6]_7 (rgf_n_277),
        .\sr_reg[6]_8 (rgf_n_279),
        .\sr_reg[6]_9 (rgf_n_281),
        .\sr_reg[7] (rgf_n_473),
        .\stat_reg[1] (rgf_n_188),
        .\stat_reg[1]_0 (rgf_n_191),
        .\stat_reg[1]_1 (rgf_n_197),
        .\stat_reg[2] (rgf_n_200),
        .\stat_reg[2]_0 (rgf_n_220),
        .\stat_reg[2]_1 (rgf_n_299),
        .\stat_reg[2]_2 (rgf_n_321),
        .\stat_reg[2]_3 (rgf_n_322),
        .tout__1_carry__0_i_1__0({rgf_n_514,rgf_n_515}),
        .tout__1_carry__0_i_7__0(fch_n_439),
        .tout__1_carry__0_i_7__0_0(fch_n_282),
        .tout__1_carry__1_i_1__0({rgf_n_520,rgf_n_521,rgf_n_522,rgf_n_523}),
        .tout__1_carry__2(fch_n_105),
        .tout__1_carry__2_0(fch_n_167),
        .tout__1_carry__2_1(fch_n_505),
        .\tr_reg[0] (rgf_n_574),
        .\tr_reg[0]_0 (rgf_n_586),
        .\tr_reg[10] (rgf_n_194),
        .\tr_reg[10]_0 (rgf_n_336),
        .\tr_reg[11] (rgf_n_193),
        .\tr_reg[11]_0 (rgf_n_232),
        .\tr_reg[11]_1 (rgf_n_335),
        .\tr_reg[12] (rgf_n_192),
        .\tr_reg[12]_0 (rgf_n_262),
        .\tr_reg[12]_1 (rgf_n_308),
        .\tr_reg[12]_2 (rgf_n_334),
        .\tr_reg[13] (rgf_n_189),
        .\tr_reg[13]_0 (rgf_n_190),
        .\tr_reg[13]_1 (rgf_n_233),
        .\tr_reg[14] (rgf_n_186),
        .\tr_reg[14]_0 (rgf_n_187),
        .\tr_reg[14]_1 (rgf_n_280),
        .\tr_reg[14]_2 (rgf_n_320),
        .\tr_reg[15] (rgf_tr),
        .\tr_reg[15]_0 (rgf_n_316),
        .\tr_reg[15]_1 (rgf_n_323),
        .\tr_reg[15]_2 (\treg/p_1_in ),
        .\tr_reg[1] (rgf_n_278),
        .\tr_reg[1]_0 (rgf_n_319),
        .\tr_reg[1]_1 (rgf_n_575),
        .\tr_reg[1]_2 (rgf_n_587),
        .\tr_reg[2] (rgf_n_576),
        .\tr_reg[2]_0 (rgf_n_588),
        .\tr_reg[3] (rgf_n_310),
        .\tr_reg[3]_0 (rgf_n_577),
        .\tr_reg[3]_1 (rgf_n_589),
        .\tr_reg[4] (rgf_n_578),
        .\tr_reg[4]_0 (rgf_n_590),
        .\tr_reg[5] (rgf_n_221),
        .\tr_reg[5]_0 (rgf_n_223),
        .\tr_reg[6] (rgf_n_201),
        .\tr_reg[6]_0 (rgf_n_219),
        .\tr_reg[7] (rgf_n_198),
        .\tr_reg[7]_0 (rgf_n_199),
        .\tr_reg[8] (rgf_n_196),
        .\tr_reg[8]_0 (rgf_n_338),
        .\tr_reg[9] (rgf_n_195),
        .\tr_reg[9]_0 (rgf_n_337));
endmodule
