
(* STRUCTURAL_NETLIST = "yes" *)
module moscoviumss
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdatx,
    fdat,
    bdatr,
    fadr,
    bcmd,
    badrx,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o);
//
//	Moscovium-SS 16 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2023/10/28	ver.1.08
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.06
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.04
//		instruction: divlqr, divlrr, divur, divsr, mulur, mulsr
//
//	2022/10/22	ver.1.02
//		corresponding to interrupt vector / level
//
//	2022/06/11	ver.1.00
//		Moscovium-SS: Super Scalar Edition
//
// ================================
//
//	2022/06/04	ver.1.12
//		instruction: csft, csfti
//		revised register file block
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [15:0]fdatx;
  input [15:0]fdat;
  input [15:0]bdatr;
  output [15:0]fadr;
  output [2:0]bcmd;
  output [15:0]badrx;
  output [15:0]badr;
  output [15:0]bdatw;
  input crdy;
  input [15:0]cbus_i;
  output [4:0]ccmd;
  output [15:0]abus_o;
  output [15:0]bbus_o;

  wire \<const0> ;
  wire \<const1> ;
  wire [15:0]a0bus_0;
  wire [15:0]a1bus_0;
  wire [15:0]abus_o;
  wire [18:18]\alu0/art/add/tout ;
  wire \alu0/art/add/tout__1_carry__0_n_0 ;
  wire \alu0/art/add/tout__1_carry__0_n_1 ;
  wire \alu0/art/add/tout__1_carry__0_n_2 ;
  wire \alu0/art/add/tout__1_carry__0_n_3 ;
  wire \alu0/art/add/tout__1_carry__0_n_4 ;
  wire \alu0/art/add/tout__1_carry__0_n_5 ;
  wire \alu0/art/add/tout__1_carry__0_n_6 ;
  wire \alu0/art/add/tout__1_carry__0_n_7 ;
  wire \alu0/art/add/tout__1_carry__1_n_0 ;
  wire \alu0/art/add/tout__1_carry__1_n_1 ;
  wire \alu0/art/add/tout__1_carry__1_n_2 ;
  wire \alu0/art/add/tout__1_carry__1_n_3 ;
  wire \alu0/art/add/tout__1_carry__1_n_4 ;
  wire \alu0/art/add/tout__1_carry__1_n_5 ;
  wire \alu0/art/add/tout__1_carry__1_n_6 ;
  wire \alu0/art/add/tout__1_carry__1_n_7 ;
  wire \alu0/art/add/tout__1_carry__2_n_0 ;
  wire \alu0/art/add/tout__1_carry__2_n_1 ;
  wire \alu0/art/add/tout__1_carry__2_n_2 ;
  wire \alu0/art/add/tout__1_carry__2_n_3 ;
  wire \alu0/art/add/tout__1_carry__2_n_5 ;
  wire \alu0/art/add/tout__1_carry__2_n_6 ;
  wire \alu0/art/add/tout__1_carry__2_n_7 ;
  wire \alu0/art/add/tout__1_carry__3_n_3 ;
  wire \alu0/art/add/tout__1_carry_n_0 ;
  wire \alu0/art/add/tout__1_carry_n_1 ;
  wire \alu0/art/add/tout__1_carry_n_2 ;
  wire \alu0/art/add/tout__1_carry_n_3 ;
  wire \alu0/art/add/tout__1_carry_n_4 ;
  wire \alu0/art/add/tout__1_carry_n_5 ;
  wire \alu0/art/add/tout__1_carry_n_6 ;
  wire \alu0/art/add/tout__1_carry_n_7 ;
  wire [15:15]\alu0/art/p_0_in ;
  wire [18:18]\alu1/art/add/tout ;
  wire \alu1/art/add/tout__1_carry__0_n_0 ;
  wire \alu1/art/add/tout__1_carry__0_n_1 ;
  wire \alu1/art/add/tout__1_carry__0_n_2 ;
  wire \alu1/art/add/tout__1_carry__0_n_3 ;
  wire \alu1/art/add/tout__1_carry__0_n_4 ;
  wire \alu1/art/add/tout__1_carry__0_n_5 ;
  wire \alu1/art/add/tout__1_carry__0_n_6 ;
  wire \alu1/art/add/tout__1_carry__0_n_7 ;
  wire \alu1/art/add/tout__1_carry__1_n_0 ;
  wire \alu1/art/add/tout__1_carry__1_n_1 ;
  wire \alu1/art/add/tout__1_carry__1_n_2 ;
  wire \alu1/art/add/tout__1_carry__1_n_3 ;
  wire \alu1/art/add/tout__1_carry__1_n_4 ;
  wire \alu1/art/add/tout__1_carry__1_n_5 ;
  wire \alu1/art/add/tout__1_carry__1_n_6 ;
  wire \alu1/art/add/tout__1_carry__1_n_7 ;
  wire \alu1/art/add/tout__1_carry__2_n_0 ;
  wire \alu1/art/add/tout__1_carry__2_n_1 ;
  wire \alu1/art/add/tout__1_carry__2_n_2 ;
  wire \alu1/art/add/tout__1_carry__2_n_3 ;
  wire \alu1/art/add/tout__1_carry__2_n_5 ;
  wire \alu1/art/add/tout__1_carry__2_n_6 ;
  wire \alu1/art/add/tout__1_carry__2_n_7 ;
  wire \alu1/art/add/tout__1_carry__3_n_3 ;
  wire \alu1/art/add/tout__1_carry_n_0 ;
  wire \alu1/art/add/tout__1_carry_n_1 ;
  wire \alu1/art/add/tout__1_carry_n_2 ;
  wire \alu1/art/add/tout__1_carry_n_3 ;
  wire \alu1/art/add/tout__1_carry_n_4 ;
  wire \alu1/art/add/tout__1_carry_n_5 ;
  wire \alu1/art/add/tout__1_carry_n_6 ;
  wire \alu1/art/add/tout__1_carry_n_7 ;
  wire [15:15]\alu1/art/p_0_in ;
  wire [0:0]alu_sr_flag1;
  wire [15:0]badr;
  wire \badr[0]_INST_0_i_12_n_0 ;
  wire \badr[0]_INST_0_i_29_n_0 ;
  wire \badr[0]_INST_0_i_29_n_1 ;
  wire \badr[0]_INST_0_i_29_n_2 ;
  wire \badr[0]_INST_0_i_29_n_3 ;
  wire \badr[0]_INST_0_i_3_n_0 ;
  wire \badr[0]_INST_0_i_44_n_0 ;
  wire \badr[0]_INST_0_i_45_n_0 ;
  wire \badr[0]_INST_0_i_46_n_0 ;
  wire \badr[0]_INST_0_i_47_n_0 ;
  wire \badr[0]_INST_0_i_48_n_0 ;
  wire \badr[0]_INST_0_i_49_n_0 ;
  wire \badr[0]_INST_0_i_50_n_0 ;
  wire \badr[0]_INST_0_i_51_n_0 ;
  wire \badr[0]_INST_0_i_52_n_0 ;
  wire \badr[0]_INST_0_i_6_n_0 ;
  wire \badr[0]_INST_0_i_9_n_0 ;
  wire \badr[10]_INST_0_i_12_n_0 ;
  wire \badr[10]_INST_0_i_3_n_0 ;
  wire \badr[10]_INST_0_i_43_n_0 ;
  wire \badr[10]_INST_0_i_44_n_0 ;
  wire \badr[10]_INST_0_i_45_n_0 ;
  wire \badr[10]_INST_0_i_46_n_0 ;
  wire \badr[10]_INST_0_i_47_n_0 ;
  wire \badr[10]_INST_0_i_48_n_0 ;
  wire \badr[10]_INST_0_i_49_n_0 ;
  wire \badr[10]_INST_0_i_50_n_0 ;
  wire \badr[10]_INST_0_i_6_n_0 ;
  wire \badr[10]_INST_0_i_9_n_0 ;
  wire \badr[11]_INST_0_i_12_n_0 ;
  wire \badr[11]_INST_0_i_29_n_0 ;
  wire \badr[11]_INST_0_i_29_n_1 ;
  wire \badr[11]_INST_0_i_29_n_2 ;
  wire \badr[11]_INST_0_i_29_n_3 ;
  wire \badr[11]_INST_0_i_3_n_0 ;
  wire \badr[11]_INST_0_i_44_n_0 ;
  wire \badr[11]_INST_0_i_45_n_0 ;
  wire \badr[11]_INST_0_i_46_n_0 ;
  wire \badr[11]_INST_0_i_47_n_0 ;
  wire \badr[11]_INST_0_i_48_n_0 ;
  wire \badr[11]_INST_0_i_49_n_0 ;
  wire \badr[11]_INST_0_i_50_n_0 ;
  wire \badr[11]_INST_0_i_51_n_0 ;
  wire \badr[11]_INST_0_i_52_n_0 ;
  wire \badr[11]_INST_0_i_53_n_0 ;
  wire \badr[11]_INST_0_i_54_n_0 ;
  wire \badr[11]_INST_0_i_55_n_0 ;
  wire \badr[11]_INST_0_i_6_n_0 ;
  wire \badr[11]_INST_0_i_9_n_0 ;
  wire \badr[12]_INST_0_i_12_n_0 ;
  wire \badr[12]_INST_0_i_3_n_0 ;
  wire \badr[12]_INST_0_i_43_n_0 ;
  wire \badr[12]_INST_0_i_44_n_0 ;
  wire \badr[12]_INST_0_i_45_n_0 ;
  wire \badr[12]_INST_0_i_46_n_0 ;
  wire \badr[12]_INST_0_i_47_n_0 ;
  wire \badr[12]_INST_0_i_48_n_0 ;
  wire \badr[12]_INST_0_i_49_n_0 ;
  wire \badr[12]_INST_0_i_50_n_0 ;
  wire \badr[12]_INST_0_i_6_n_0 ;
  wire \badr[12]_INST_0_i_9_n_0 ;
  wire \badr[13]_INST_0_i_12_n_0 ;
  wire \badr[13]_INST_0_i_3_n_0 ;
  wire \badr[13]_INST_0_i_43_n_0 ;
  wire \badr[13]_INST_0_i_44_n_0 ;
  wire \badr[13]_INST_0_i_45_n_0 ;
  wire \badr[13]_INST_0_i_46_n_0 ;
  wire \badr[13]_INST_0_i_47_n_0 ;
  wire \badr[13]_INST_0_i_48_n_0 ;
  wire \badr[13]_INST_0_i_49_n_0 ;
  wire \badr[13]_INST_0_i_50_n_0 ;
  wire \badr[13]_INST_0_i_6_n_0 ;
  wire \badr[13]_INST_0_i_9_n_0 ;
  wire \badr[14]_INST_0_i_12_n_0 ;
  wire \badr[14]_INST_0_i_3_n_0 ;
  wire \badr[14]_INST_0_i_43_n_0 ;
  wire \badr[14]_INST_0_i_44_n_0 ;
  wire \badr[14]_INST_0_i_45_n_0 ;
  wire \badr[14]_INST_0_i_46_n_0 ;
  wire \badr[14]_INST_0_i_47_n_0 ;
  wire \badr[14]_INST_0_i_48_n_0 ;
  wire \badr[14]_INST_0_i_49_n_0 ;
  wire \badr[14]_INST_0_i_50_n_0 ;
  wire \badr[14]_INST_0_i_6_n_0 ;
  wire \badr[14]_INST_0_i_9_n_0 ;
  wire \badr[15]_INST_0_i_104_n_0 ;
  wire \badr[15]_INST_0_i_105_n_0 ;
  wire \badr[15]_INST_0_i_108_n_0 ;
  wire \badr[15]_INST_0_i_109_n_0 ;
  wire \badr[15]_INST_0_i_110_n_0 ;
  wire \badr[15]_INST_0_i_111_n_0 ;
  wire \badr[15]_INST_0_i_112_n_0 ;
  wire \badr[15]_INST_0_i_113_n_0 ;
  wire \badr[15]_INST_0_i_114_n_0 ;
  wire \badr[15]_INST_0_i_115_n_0 ;
  wire \badr[15]_INST_0_i_116_n_0 ;
  wire \badr[15]_INST_0_i_117_n_0 ;
  wire \badr[15]_INST_0_i_118_n_0 ;
  wire \badr[15]_INST_0_i_120_n_0 ;
  wire \badr[15]_INST_0_i_121_n_0 ;
  wire \badr[15]_INST_0_i_122_n_0 ;
  wire \badr[15]_INST_0_i_123_n_0 ;
  wire \badr[15]_INST_0_i_12_n_0 ;
  wire \badr[15]_INST_0_i_140_n_0 ;
  wire \badr[15]_INST_0_i_141_n_0 ;
  wire \badr[15]_INST_0_i_142_n_0 ;
  wire \badr[15]_INST_0_i_143_n_0 ;
  wire \badr[15]_INST_0_i_144_n_0 ;
  wire \badr[15]_INST_0_i_145_n_0 ;
  wire \badr[15]_INST_0_i_146_n_0 ;
  wire \badr[15]_INST_0_i_147_n_0 ;
  wire \badr[15]_INST_0_i_148_n_0 ;
  wire \badr[15]_INST_0_i_159_n_0 ;
  wire \badr[15]_INST_0_i_15_n_0 ;
  wire \badr[15]_INST_0_i_160_n_0 ;
  wire \badr[15]_INST_0_i_163_n_0 ;
  wire \badr[15]_INST_0_i_164_n_0 ;
  wire \badr[15]_INST_0_i_165_n_0 ;
  wire \badr[15]_INST_0_i_166_n_0 ;
  wire \badr[15]_INST_0_i_167_n_0 ;
  wire \badr[15]_INST_0_i_168_n_0 ;
  wire \badr[15]_INST_0_i_169_n_0 ;
  wire \badr[15]_INST_0_i_170_n_0 ;
  wire \badr[15]_INST_0_i_171_n_0 ;
  wire \badr[15]_INST_0_i_172_n_0 ;
  wire \badr[15]_INST_0_i_173_n_0 ;
  wire \badr[15]_INST_0_i_174_n_0 ;
  wire \badr[15]_INST_0_i_175_n_0 ;
  wire \badr[15]_INST_0_i_176_n_0 ;
  wire \badr[15]_INST_0_i_177_n_0 ;
  wire \badr[15]_INST_0_i_178_n_0 ;
  wire \badr[15]_INST_0_i_179_n_0 ;
  wire \badr[15]_INST_0_i_17_n_0 ;
  wire \badr[15]_INST_0_i_180_n_0 ;
  wire \badr[15]_INST_0_i_181_n_0 ;
  wire \badr[15]_INST_0_i_182_n_0 ;
  wire \badr[15]_INST_0_i_183_n_0 ;
  wire \badr[15]_INST_0_i_184_n_0 ;
  wire \badr[15]_INST_0_i_185_n_0 ;
  wire \badr[15]_INST_0_i_186_n_0 ;
  wire \badr[15]_INST_0_i_187_n_0 ;
  wire \badr[15]_INST_0_i_188_n_0 ;
  wire \badr[15]_INST_0_i_189_n_0 ;
  wire \badr[15]_INST_0_i_18_n_0 ;
  wire \badr[15]_INST_0_i_190_n_0 ;
  wire \badr[15]_INST_0_i_191_n_0 ;
  wire \badr[15]_INST_0_i_192_n_0 ;
  wire \badr[15]_INST_0_i_193_n_0 ;
  wire \badr[15]_INST_0_i_194_n_0 ;
  wire \badr[15]_INST_0_i_195_n_0 ;
  wire \badr[15]_INST_0_i_196_n_0 ;
  wire \badr[15]_INST_0_i_197_n_0 ;
  wire \badr[15]_INST_0_i_198_n_0 ;
  wire \badr[15]_INST_0_i_199_n_0 ;
  wire \badr[15]_INST_0_i_200_n_0 ;
  wire \badr[15]_INST_0_i_201_n_0 ;
  wire \badr[15]_INST_0_i_202_n_0 ;
  wire \badr[15]_INST_0_i_203_n_0 ;
  wire \badr[15]_INST_0_i_204_n_0 ;
  wire \badr[15]_INST_0_i_205_n_0 ;
  wire \badr[15]_INST_0_i_206_n_0 ;
  wire \badr[15]_INST_0_i_207_n_0 ;
  wire \badr[15]_INST_0_i_208_n_0 ;
  wire \badr[15]_INST_0_i_210_n_0 ;
  wire \badr[15]_INST_0_i_211_n_0 ;
  wire \badr[15]_INST_0_i_212_n_0 ;
  wire \badr[15]_INST_0_i_213_n_0 ;
  wire \badr[15]_INST_0_i_214_n_0 ;
  wire \badr[15]_INST_0_i_215_n_0 ;
  wire \badr[15]_INST_0_i_216_n_0 ;
  wire \badr[15]_INST_0_i_217_n_0 ;
  wire \badr[15]_INST_0_i_218_n_0 ;
  wire \badr[15]_INST_0_i_219_n_0 ;
  wire \badr[15]_INST_0_i_220_n_0 ;
  wire \badr[15]_INST_0_i_221_n_0 ;
  wire \badr[15]_INST_0_i_222_n_0 ;
  wire \badr[15]_INST_0_i_223_n_0 ;
  wire \badr[15]_INST_0_i_224_n_0 ;
  wire \badr[15]_INST_0_i_225_n_0 ;
  wire \badr[15]_INST_0_i_226_n_0 ;
  wire \badr[15]_INST_0_i_227_n_0 ;
  wire \badr[15]_INST_0_i_228_n_0 ;
  wire \badr[15]_INST_0_i_229_n_0 ;
  wire \badr[15]_INST_0_i_230_n_0 ;
  wire \badr[15]_INST_0_i_231_n_0 ;
  wire \badr[15]_INST_0_i_232_n_0 ;
  wire \badr[15]_INST_0_i_233_n_0 ;
  wire \badr[15]_INST_0_i_234_n_0 ;
  wire \badr[15]_INST_0_i_235_n_0 ;
  wire \badr[15]_INST_0_i_236_n_0 ;
  wire \badr[15]_INST_0_i_237_n_0 ;
  wire \badr[15]_INST_0_i_238_n_0 ;
  wire \badr[15]_INST_0_i_239_n_0 ;
  wire \badr[15]_INST_0_i_240_n_0 ;
  wire \badr[15]_INST_0_i_241_n_0 ;
  wire \badr[15]_INST_0_i_242_n_0 ;
  wire \badr[15]_INST_0_i_243_n_0 ;
  wire \badr[15]_INST_0_i_244_n_0 ;
  wire \badr[15]_INST_0_i_245_n_0 ;
  wire \badr[15]_INST_0_i_246_n_0 ;
  wire \badr[15]_INST_0_i_247_n_0 ;
  wire \badr[15]_INST_0_i_248_n_0 ;
  wire \badr[15]_INST_0_i_249_n_0 ;
  wire \badr[15]_INST_0_i_250_n_0 ;
  wire \badr[15]_INST_0_i_251_n_0 ;
  wire \badr[15]_INST_0_i_252_n_0 ;
  wire \badr[15]_INST_0_i_253_n_0 ;
  wire \badr[15]_INST_0_i_254_n_0 ;
  wire \badr[15]_INST_0_i_255_n_0 ;
  wire \badr[15]_INST_0_i_256_n_0 ;
  wire \badr[15]_INST_0_i_257_n_0 ;
  wire \badr[15]_INST_0_i_258_n_0 ;
  wire \badr[15]_INST_0_i_259_n_0 ;
  wire \badr[15]_INST_0_i_260_n_0 ;
  wire \badr[15]_INST_0_i_261_n_0 ;
  wire \badr[15]_INST_0_i_262_n_0 ;
  wire \badr[15]_INST_0_i_263_n_0 ;
  wire \badr[15]_INST_0_i_264_n_0 ;
  wire \badr[15]_INST_0_i_265_n_0 ;
  wire \badr[15]_INST_0_i_266_n_0 ;
  wire \badr[15]_INST_0_i_267_n_0 ;
  wire \badr[15]_INST_0_i_268_n_0 ;
  wire \badr[15]_INST_0_i_269_n_0 ;
  wire \badr[15]_INST_0_i_270_n_0 ;
  wire \badr[15]_INST_0_i_271_n_0 ;
  wire \badr[15]_INST_0_i_272_n_0 ;
  wire \badr[15]_INST_0_i_273_n_0 ;
  wire \badr[15]_INST_0_i_274_n_0 ;
  wire \badr[15]_INST_0_i_275_n_0 ;
  wire \badr[15]_INST_0_i_276_n_0 ;
  wire \badr[15]_INST_0_i_277_n_0 ;
  wire \badr[15]_INST_0_i_278_n_0 ;
  wire \badr[15]_INST_0_i_279_n_0 ;
  wire \badr[15]_INST_0_i_280_n_0 ;
  wire \badr[15]_INST_0_i_281_n_0 ;
  wire \badr[15]_INST_0_i_282_n_0 ;
  wire \badr[15]_INST_0_i_283_n_0 ;
  wire \badr[15]_INST_0_i_284_n_0 ;
  wire \badr[15]_INST_0_i_285_n_0 ;
  wire \badr[15]_INST_0_i_286_n_0 ;
  wire \badr[15]_INST_0_i_287_n_0 ;
  wire \badr[15]_INST_0_i_288_n_0 ;
  wire \badr[15]_INST_0_i_289_n_0 ;
  wire \badr[15]_INST_0_i_28_n_0 ;
  wire \badr[15]_INST_0_i_290_n_0 ;
  wire \badr[15]_INST_0_i_291_n_0 ;
  wire \badr[15]_INST_0_i_292_n_0 ;
  wire \badr[15]_INST_0_i_293_n_0 ;
  wire \badr[15]_INST_0_i_294_n_0 ;
  wire \badr[15]_INST_0_i_295_n_0 ;
  wire \badr[15]_INST_0_i_296_n_0 ;
  wire \badr[15]_INST_0_i_297_n_0 ;
  wire \badr[15]_INST_0_i_298_n_0 ;
  wire \badr[15]_INST_0_i_299_n_0 ;
  wire \badr[15]_INST_0_i_300_n_0 ;
  wire \badr[15]_INST_0_i_301_n_0 ;
  wire \badr[15]_INST_0_i_302_n_0 ;
  wire \badr[15]_INST_0_i_303_n_0 ;
  wire \badr[15]_INST_0_i_304_n_0 ;
  wire \badr[15]_INST_0_i_305_n_0 ;
  wire \badr[15]_INST_0_i_306_n_0 ;
  wire \badr[15]_INST_0_i_307_n_0 ;
  wire \badr[15]_INST_0_i_308_n_0 ;
  wire \badr[15]_INST_0_i_309_n_0 ;
  wire \badr[15]_INST_0_i_310_n_0 ;
  wire \badr[15]_INST_0_i_311_n_0 ;
  wire \badr[15]_INST_0_i_312_n_0 ;
  wire \badr[15]_INST_0_i_313_n_0 ;
  wire \badr[15]_INST_0_i_314_n_0 ;
  wire \badr[15]_INST_0_i_315_n_0 ;
  wire \badr[15]_INST_0_i_316_n_0 ;
  wire \badr[15]_INST_0_i_317_n_0 ;
  wire \badr[15]_INST_0_i_318_n_0 ;
  wire \badr[15]_INST_0_i_319_n_0 ;
  wire \badr[15]_INST_0_i_320_n_0 ;
  wire \badr[15]_INST_0_i_321_n_0 ;
  wire \badr[15]_INST_0_i_322_n_0 ;
  wire \badr[15]_INST_0_i_323_n_0 ;
  wire \badr[15]_INST_0_i_324_n_0 ;
  wire \badr[15]_INST_0_i_325_n_0 ;
  wire \badr[15]_INST_0_i_326_n_0 ;
  wire \badr[15]_INST_0_i_327_n_0 ;
  wire \badr[15]_INST_0_i_328_n_0 ;
  wire \badr[15]_INST_0_i_329_n_0 ;
  wire \badr[15]_INST_0_i_36_n_1 ;
  wire \badr[15]_INST_0_i_36_n_2 ;
  wire \badr[15]_INST_0_i_36_n_3 ;
  wire \badr[15]_INST_0_i_39_n_0 ;
  wire \badr[15]_INST_0_i_3_n_0 ;
  wire \badr[15]_INST_0_i_40_n_0 ;
  wire \badr[15]_INST_0_i_41_n_0 ;
  wire \badr[15]_INST_0_i_42_n_0 ;
  wire \badr[15]_INST_0_i_52_n_0 ;
  wire \badr[15]_INST_0_i_62_n_0 ;
  wire \badr[15]_INST_0_i_63_n_0 ;
  wire \badr[15]_INST_0_i_64_n_0 ;
  wire \badr[15]_INST_0_i_65_n_0 ;
  wire \badr[15]_INST_0_i_67_n_0 ;
  wire \badr[15]_INST_0_i_68_n_0 ;
  wire \badr[15]_INST_0_i_69_n_0 ;
  wire \badr[15]_INST_0_i_6_n_0 ;
  wire \badr[15]_INST_0_i_70_n_0 ;
  wire \badr[15]_INST_0_i_87_n_0 ;
  wire \badr[15]_INST_0_i_88_n_0 ;
  wire \badr[15]_INST_0_i_89_n_0 ;
  wire \badr[15]_INST_0_i_90_n_0 ;
  wire \badr[15]_INST_0_i_91_n_0 ;
  wire \badr[15]_INST_0_i_92_n_0 ;
  wire \badr[15]_INST_0_i_93_n_0 ;
  wire \badr[15]_INST_0_i_9_n_0 ;
  wire \badr[1]_INST_0_i_12_n_0 ;
  wire \badr[1]_INST_0_i_3_n_0 ;
  wire \badr[1]_INST_0_i_43_n_0 ;
  wire \badr[1]_INST_0_i_44_n_0 ;
  wire \badr[1]_INST_0_i_45_n_0 ;
  wire \badr[1]_INST_0_i_46_n_0 ;
  wire \badr[1]_INST_0_i_47_n_0 ;
  wire \badr[1]_INST_0_i_48_n_0 ;
  wire \badr[1]_INST_0_i_49_n_0 ;
  wire \badr[1]_INST_0_i_50_n_0 ;
  wire \badr[1]_INST_0_i_6_n_0 ;
  wire \badr[1]_INST_0_i_9_n_0 ;
  wire \badr[2]_INST_0_i_12_n_0 ;
  wire \badr[2]_INST_0_i_3_n_0 ;
  wire \badr[2]_INST_0_i_43_n_0 ;
  wire \badr[2]_INST_0_i_44_n_0 ;
  wire \badr[2]_INST_0_i_45_n_0 ;
  wire \badr[2]_INST_0_i_46_n_0 ;
  wire \badr[2]_INST_0_i_47_n_0 ;
  wire \badr[2]_INST_0_i_48_n_0 ;
  wire \badr[2]_INST_0_i_49_n_0 ;
  wire \badr[2]_INST_0_i_50_n_0 ;
  wire \badr[2]_INST_0_i_6_n_0 ;
  wire \badr[2]_INST_0_i_9_n_0 ;
  wire \badr[3]_INST_0_i_12_n_0 ;
  wire \badr[3]_INST_0_i_29_n_0 ;
  wire \badr[3]_INST_0_i_29_n_1 ;
  wire \badr[3]_INST_0_i_29_n_2 ;
  wire \badr[3]_INST_0_i_29_n_3 ;
  wire \badr[3]_INST_0_i_3_n_0 ;
  wire \badr[3]_INST_0_i_44_n_0 ;
  wire \badr[3]_INST_0_i_45_n_0 ;
  wire \badr[3]_INST_0_i_46_n_0 ;
  wire \badr[3]_INST_0_i_47_n_0 ;
  wire \badr[3]_INST_0_i_48_n_0 ;
  wire \badr[3]_INST_0_i_49_n_0 ;
  wire \badr[3]_INST_0_i_50_n_0 ;
  wire \badr[3]_INST_0_i_51_n_0 ;
  wire \badr[3]_INST_0_i_52_n_0 ;
  wire \badr[3]_INST_0_i_53_n_0 ;
  wire \badr[3]_INST_0_i_54_n_0 ;
  wire \badr[3]_INST_0_i_6_n_0 ;
  wire \badr[3]_INST_0_i_9_n_0 ;
  wire \badr[4]_INST_0_i_12_n_0 ;
  wire \badr[4]_INST_0_i_3_n_0 ;
  wire \badr[4]_INST_0_i_43_n_0 ;
  wire \badr[4]_INST_0_i_44_n_0 ;
  wire \badr[4]_INST_0_i_45_n_0 ;
  wire \badr[4]_INST_0_i_46_n_0 ;
  wire \badr[4]_INST_0_i_47_n_0 ;
  wire \badr[4]_INST_0_i_48_n_0 ;
  wire \badr[4]_INST_0_i_49_n_0 ;
  wire \badr[4]_INST_0_i_50_n_0 ;
  wire \badr[4]_INST_0_i_6_n_0 ;
  wire \badr[4]_INST_0_i_9_n_0 ;
  wire \badr[5]_INST_0_i_12_n_0 ;
  wire \badr[5]_INST_0_i_3_n_0 ;
  wire \badr[5]_INST_0_i_43_n_0 ;
  wire \badr[5]_INST_0_i_44_n_0 ;
  wire \badr[5]_INST_0_i_45_n_0 ;
  wire \badr[5]_INST_0_i_46_n_0 ;
  wire \badr[5]_INST_0_i_47_n_0 ;
  wire \badr[5]_INST_0_i_48_n_0 ;
  wire \badr[5]_INST_0_i_49_n_0 ;
  wire \badr[5]_INST_0_i_50_n_0 ;
  wire \badr[5]_INST_0_i_6_n_0 ;
  wire \badr[5]_INST_0_i_9_n_0 ;
  wire \badr[6]_INST_0_i_12_n_0 ;
  wire \badr[6]_INST_0_i_3_n_0 ;
  wire \badr[6]_INST_0_i_43_n_0 ;
  wire \badr[6]_INST_0_i_44_n_0 ;
  wire \badr[6]_INST_0_i_45_n_0 ;
  wire \badr[6]_INST_0_i_46_n_0 ;
  wire \badr[6]_INST_0_i_47_n_0 ;
  wire \badr[6]_INST_0_i_48_n_0 ;
  wire \badr[6]_INST_0_i_49_n_0 ;
  wire \badr[6]_INST_0_i_50_n_0 ;
  wire \badr[6]_INST_0_i_6_n_0 ;
  wire \badr[6]_INST_0_i_9_n_0 ;
  wire \badr[7]_INST_0_i_12_n_0 ;
  wire \badr[7]_INST_0_i_29_n_0 ;
  wire \badr[7]_INST_0_i_29_n_1 ;
  wire \badr[7]_INST_0_i_29_n_2 ;
  wire \badr[7]_INST_0_i_29_n_3 ;
  wire \badr[7]_INST_0_i_3_n_0 ;
  wire \badr[7]_INST_0_i_44_n_0 ;
  wire \badr[7]_INST_0_i_45_n_0 ;
  wire \badr[7]_INST_0_i_46_n_0 ;
  wire \badr[7]_INST_0_i_47_n_0 ;
  wire \badr[7]_INST_0_i_48_n_0 ;
  wire \badr[7]_INST_0_i_49_n_0 ;
  wire \badr[7]_INST_0_i_50_n_0 ;
  wire \badr[7]_INST_0_i_51_n_0 ;
  wire \badr[7]_INST_0_i_52_n_0 ;
  wire \badr[7]_INST_0_i_53_n_0 ;
  wire \badr[7]_INST_0_i_54_n_0 ;
  wire \badr[7]_INST_0_i_55_n_0 ;
  wire \badr[7]_INST_0_i_6_n_0 ;
  wire \badr[7]_INST_0_i_9_n_0 ;
  wire \badr[8]_INST_0_i_12_n_0 ;
  wire \badr[8]_INST_0_i_3_n_0 ;
  wire \badr[8]_INST_0_i_43_n_0 ;
  wire \badr[8]_INST_0_i_44_n_0 ;
  wire \badr[8]_INST_0_i_45_n_0 ;
  wire \badr[8]_INST_0_i_46_n_0 ;
  wire \badr[8]_INST_0_i_47_n_0 ;
  wire \badr[8]_INST_0_i_48_n_0 ;
  wire \badr[8]_INST_0_i_49_n_0 ;
  wire \badr[8]_INST_0_i_50_n_0 ;
  wire \badr[8]_INST_0_i_6_n_0 ;
  wire \badr[8]_INST_0_i_9_n_0 ;
  wire \badr[9]_INST_0_i_12_n_0 ;
  wire \badr[9]_INST_0_i_3_n_0 ;
  wire \badr[9]_INST_0_i_43_n_0 ;
  wire \badr[9]_INST_0_i_44_n_0 ;
  wire \badr[9]_INST_0_i_45_n_0 ;
  wire \badr[9]_INST_0_i_46_n_0 ;
  wire \badr[9]_INST_0_i_47_n_0 ;
  wire \badr[9]_INST_0_i_48_n_0 ;
  wire \badr[9]_INST_0_i_49_n_0 ;
  wire \badr[9]_INST_0_i_50_n_0 ;
  wire \badr[9]_INST_0_i_6_n_0 ;
  wire \badr[9]_INST_0_i_9_n_0 ;
  wire [15:0]badrx;
  wire \badrx[15]_INST_0_i_1_n_0 ;
  wire \badrx[15]_INST_0_i_2_n_0 ;
  wire \badrx[15]_INST_0_i_3_n_0 ;
  wire \badrx[15]_INST_0_i_4_n_0 ;
  wire \badrx[15]_INST_0_i_5_n_0 ;
  wire \bank02/a0buso/gr0_bus1 ;
  wire \bank02/a0buso/gr1_bus1 ;
  wire \bank02/a0buso/gr2_bus1 ;
  wire \bank02/a0buso/gr3_bus1 ;
  wire \bank02/a0buso/gr4_bus1 ;
  wire \bank02/a0buso/gr5_bus1 ;
  wire \bank02/a0buso/gr6_bus1 ;
  wire \bank02/a0buso/gr7_bus1 ;
  wire \bank02/a0buso2l/gr0_bus1 ;
  wire \bank02/a0buso2l/gr1_bus1 ;
  wire \bank02/a0buso2l/gr2_bus1 ;
  wire \bank02/a0buso2l/gr3_bus1 ;
  wire \bank02/a0buso2l/gr4_bus1 ;
  wire \bank02/a0buso2l/gr5_bus1 ;
  wire \bank02/a0buso2l/gr6_bus1 ;
  wire \bank02/a0buso2l/gr7_bus1 ;
  wire \bank02/a1buso/gr0_bus1 ;
  wire \bank02/a1buso/gr1_bus1 ;
  wire \bank02/a1buso/gr2_bus1 ;
  wire \bank02/a1buso/gr3_bus1 ;
  wire \bank02/a1buso/gr4_bus1 ;
  wire \bank02/a1buso/gr5_bus1 ;
  wire \bank02/a1buso/gr6_bus1 ;
  wire \bank02/a1buso/gr7_bus1 ;
  wire \bank02/a1buso2l/gr0_bus1 ;
  wire \bank02/a1buso2l/gr1_bus1 ;
  wire \bank02/a1buso2l/gr2_bus1 ;
  wire \bank02/a1buso2l/gr3_bus1 ;
  wire \bank02/a1buso2l/gr4_bus1 ;
  wire \bank02/a1buso2l/gr5_bus1 ;
  wire \bank02/a1buso2l/gr6_bus1 ;
  wire \bank02/a1buso2l/gr7_bus1 ;
  wire \bank02/b0buso/gr0_bus1 ;
  wire \bank02/b0buso/gr1_bus1 ;
  wire \bank02/b0buso/gr2_bus1 ;
  wire \bank02/b0buso/gr3_bus1 ;
  wire \bank02/b0buso/gr4_bus1 ;
  wire \bank02/b0buso/gr5_bus1 ;
  wire \bank02/b0buso/gr6_bus1 ;
  wire \bank02/b0buso/gr7_bus1 ;
  wire \bank02/b0buso2l/gr0_bus1 ;
  wire \bank02/b0buso2l/gr1_bus1 ;
  wire \bank02/b0buso2l/gr2_bus1 ;
  wire \bank02/b0buso2l/gr3_bus1 ;
  wire \bank02/b0buso2l/gr4_bus1 ;
  wire \bank02/b0buso2l/gr5_bus1 ;
  wire \bank02/b0buso2l/gr6_bus1 ;
  wire \bank02/b0buso2l/gr7_bus1 ;
  wire \bank02/b1buso/gr0_bus1 ;
  wire \bank02/b1buso/gr1_bus1 ;
  wire \bank02/b1buso/gr2_bus1 ;
  wire \bank02/b1buso/gr3_bus1 ;
  wire \bank02/b1buso/gr4_bus1 ;
  wire \bank02/b1buso/gr5_bus1 ;
  wire \bank02/b1buso/gr6_bus1 ;
  wire \bank02/b1buso/gr7_bus1 ;
  wire \bank02/b1buso2l/gr0_bus1 ;
  wire \bank02/b1buso2l/gr1_bus1 ;
  wire \bank02/b1buso2l/gr2_bus1 ;
  wire \bank02/b1buso2l/gr3_bus1 ;
  wire \bank02/b1buso2l/gr4_bus1 ;
  wire \bank02/b1buso2l/gr5_bus1 ;
  wire \bank02/b1buso2l/gr6_bus1 ;
  wire \bank02/b1buso2l/gr7_bus1 ;
  wire \bank02/grn01/grn[0]_i_1_n_0 ;
  wire \bank02/grn01/grn[10]_i_1_n_0 ;
  wire \bank02/grn01/grn[11]_i_1_n_0 ;
  wire \bank02/grn01/grn[12]_i_1_n_0 ;
  wire \bank02/grn01/grn[13]_i_1_n_0 ;
  wire \bank02/grn01/grn[14]_i_1_n_0 ;
  wire \bank02/grn01/grn[15]_i_2_n_0 ;
  wire \bank02/grn01/grn[1]_i_1_n_0 ;
  wire \bank02/grn01/grn[2]_i_1_n_0 ;
  wire \bank02/grn01/grn[3]_i_1_n_0 ;
  wire \bank02/grn01/grn[4]_i_1_n_0 ;
  wire \bank02/grn01/grn[5]_i_1_n_0 ;
  wire \bank02/grn01/grn[6]_i_1_n_0 ;
  wire \bank02/grn01/grn[7]_i_1_n_0 ;
  wire \bank02/grn01/grn[8]_i_1_n_0 ;
  wire \bank02/grn01/grn[9]_i_1_n_0 ;
  wire \bank02/grn02/grn[0]_i_1_n_0 ;
  wire \bank02/grn02/grn[10]_i_1_n_0 ;
  wire \bank02/grn02/grn[11]_i_1_n_0 ;
  wire \bank02/grn02/grn[12]_i_1_n_0 ;
  wire \bank02/grn02/grn[13]_i_1_n_0 ;
  wire \bank02/grn02/grn[14]_i_1_n_0 ;
  wire \bank02/grn02/grn[15]_i_2_n_0 ;
  wire \bank02/grn02/grn[1]_i_1_n_0 ;
  wire \bank02/grn02/grn[2]_i_1_n_0 ;
  wire \bank02/grn02/grn[3]_i_1_n_0 ;
  wire \bank02/grn02/grn[4]_i_1_n_0 ;
  wire \bank02/grn02/grn[5]_i_1_n_0 ;
  wire \bank02/grn02/grn[6]_i_1_n_0 ;
  wire \bank02/grn02/grn[7]_i_1_n_0 ;
  wire \bank02/grn02/grn[8]_i_1_n_0 ;
  wire \bank02/grn02/grn[9]_i_1_n_0 ;
  wire \bank02/grn03/grn[0]_i_1_n_0 ;
  wire \bank02/grn03/grn[10]_i_1_n_0 ;
  wire \bank02/grn03/grn[11]_i_1_n_0 ;
  wire \bank02/grn03/grn[12]_i_1_n_0 ;
  wire \bank02/grn03/grn[13]_i_1_n_0 ;
  wire \bank02/grn03/grn[14]_i_1_n_0 ;
  wire \bank02/grn03/grn[15]_i_2_n_0 ;
  wire \bank02/grn03/grn[1]_i_1_n_0 ;
  wire \bank02/grn03/grn[2]_i_1_n_0 ;
  wire \bank02/grn03/grn[3]_i_1_n_0 ;
  wire \bank02/grn03/grn[4]_i_1_n_0 ;
  wire \bank02/grn03/grn[5]_i_1_n_0 ;
  wire \bank02/grn03/grn[6]_i_1_n_0 ;
  wire \bank02/grn03/grn[7]_i_1_n_0 ;
  wire \bank02/grn03/grn[8]_i_1_n_0 ;
  wire \bank02/grn03/grn[9]_i_1_n_0 ;
  wire \bank02/grn04/grn[0]_i_1_n_0 ;
  wire \bank02/grn04/grn[10]_i_1_n_0 ;
  wire \bank02/grn04/grn[11]_i_1_n_0 ;
  wire \bank02/grn04/grn[12]_i_1_n_0 ;
  wire \bank02/grn04/grn[13]_i_1_n_0 ;
  wire \bank02/grn04/grn[14]_i_1_n_0 ;
  wire \bank02/grn04/grn[15]_i_2_n_0 ;
  wire \bank02/grn04/grn[1]_i_1_n_0 ;
  wire \bank02/grn04/grn[2]_i_1_n_0 ;
  wire \bank02/grn04/grn[3]_i_1_n_0 ;
  wire \bank02/grn04/grn[4]_i_1_n_0 ;
  wire \bank02/grn04/grn[5]_i_1_n_0 ;
  wire \bank02/grn04/grn[6]_i_1_n_0 ;
  wire \bank02/grn04/grn[7]_i_1_n_0 ;
  wire \bank02/grn04/grn[8]_i_1_n_0 ;
  wire \bank02/grn04/grn[9]_i_1_n_0 ;
  wire \bank02/grn05/grn[0]_i_1_n_0 ;
  wire \bank02/grn05/grn[10]_i_1_n_0 ;
  wire \bank02/grn05/grn[11]_i_1_n_0 ;
  wire \bank02/grn05/grn[12]_i_1_n_0 ;
  wire \bank02/grn05/grn[13]_i_1_n_0 ;
  wire \bank02/grn05/grn[14]_i_1_n_0 ;
  wire \bank02/grn05/grn[15]_i_2_n_0 ;
  wire \bank02/grn05/grn[1]_i_1_n_0 ;
  wire \bank02/grn05/grn[2]_i_1_n_0 ;
  wire \bank02/grn05/grn[3]_i_1_n_0 ;
  wire \bank02/grn05/grn[4]_i_1_n_0 ;
  wire \bank02/grn05/grn[5]_i_1_n_0 ;
  wire \bank02/grn05/grn[6]_i_1_n_0 ;
  wire \bank02/grn05/grn[7]_i_1_n_0 ;
  wire \bank02/grn05/grn[8]_i_1_n_0 ;
  wire \bank02/grn05/grn[9]_i_1_n_0 ;
  wire \bank02/grn06/grn[0]_i_1_n_0 ;
  wire \bank02/grn06/grn[10]_i_1_n_0 ;
  wire \bank02/grn06/grn[11]_i_1_n_0 ;
  wire \bank02/grn06/grn[12]_i_1_n_0 ;
  wire \bank02/grn06/grn[13]_i_1_n_0 ;
  wire \bank02/grn06/grn[14]_i_1_n_0 ;
  wire \bank02/grn06/grn[15]_i_2_n_0 ;
  wire \bank02/grn06/grn[1]_i_1_n_0 ;
  wire \bank02/grn06/grn[2]_i_1_n_0 ;
  wire \bank02/grn06/grn[3]_i_1_n_0 ;
  wire \bank02/grn06/grn[4]_i_1_n_0 ;
  wire \bank02/grn06/grn[5]_i_1_n_0 ;
  wire \bank02/grn06/grn[6]_i_1_n_0 ;
  wire \bank02/grn06/grn[7]_i_1_n_0 ;
  wire \bank02/grn06/grn[8]_i_1_n_0 ;
  wire \bank02/grn06/grn[9]_i_1_n_0 ;
  wire \bank02/grn07/grn[0]_i_1_n_0 ;
  wire \bank02/grn07/grn[10]_i_1_n_0 ;
  wire \bank02/grn07/grn[11]_i_1_n_0 ;
  wire \bank02/grn07/grn[12]_i_1_n_0 ;
  wire \bank02/grn07/grn[13]_i_1_n_0 ;
  wire \bank02/grn07/grn[14]_i_1_n_0 ;
  wire \bank02/grn07/grn[15]_i_2_n_0 ;
  wire \bank02/grn07/grn[1]_i_1_n_0 ;
  wire \bank02/grn07/grn[2]_i_1_n_0 ;
  wire \bank02/grn07/grn[3]_i_1_n_0 ;
  wire \bank02/grn07/grn[4]_i_1_n_0 ;
  wire \bank02/grn07/grn[5]_i_1_n_0 ;
  wire \bank02/grn07/grn[6]_i_1_n_0 ;
  wire \bank02/grn07/grn[7]_i_1_n_0 ;
  wire \bank02/grn07/grn[8]_i_1_n_0 ;
  wire \bank02/grn07/grn[9]_i_1_n_0 ;
  wire \bank02/grn20/grn[0]_i_1_n_0 ;
  wire \bank02/grn20/grn[10]_i_1_n_0 ;
  wire \bank02/grn20/grn[11]_i_1_n_0 ;
  wire \bank02/grn20/grn[12]_i_1_n_0 ;
  wire \bank02/grn20/grn[13]_i_1_n_0 ;
  wire \bank02/grn20/grn[14]_i_1_n_0 ;
  wire \bank02/grn20/grn[15]_i_2_n_0 ;
  wire \bank02/grn20/grn[1]_i_1_n_0 ;
  wire \bank02/grn20/grn[2]_i_1_n_0 ;
  wire \bank02/grn20/grn[3]_i_1_n_0 ;
  wire \bank02/grn20/grn[4]_i_1_n_0 ;
  wire \bank02/grn20/grn[5]_i_1_n_0 ;
  wire \bank02/grn20/grn[6]_i_1_n_0 ;
  wire \bank02/grn20/grn[7]_i_1_n_0 ;
  wire \bank02/grn20/grn[8]_i_1_n_0 ;
  wire \bank02/grn20/grn[9]_i_1_n_0 ;
  wire \bank02/grn21/grn[0]_i_1_n_0 ;
  wire \bank02/grn21/grn[10]_i_1_n_0 ;
  wire \bank02/grn21/grn[11]_i_1_n_0 ;
  wire \bank02/grn21/grn[12]_i_1_n_0 ;
  wire \bank02/grn21/grn[13]_i_1_n_0 ;
  wire \bank02/grn21/grn[14]_i_1_n_0 ;
  wire \bank02/grn21/grn[15]_i_2_n_0 ;
  wire \bank02/grn21/grn[1]_i_1_n_0 ;
  wire \bank02/grn21/grn[2]_i_1_n_0 ;
  wire \bank02/grn21/grn[3]_i_1_n_0 ;
  wire \bank02/grn21/grn[4]_i_1_n_0 ;
  wire \bank02/grn21/grn[5]_i_1_n_0 ;
  wire \bank02/grn21/grn[6]_i_1_n_0 ;
  wire \bank02/grn21/grn[7]_i_1_n_0 ;
  wire \bank02/grn21/grn[8]_i_1_n_0 ;
  wire \bank02/grn21/grn[9]_i_1_n_0 ;
  wire \bank02/grn22/grn[0]_i_1_n_0 ;
  wire \bank02/grn22/grn[10]_i_1_n_0 ;
  wire \bank02/grn22/grn[11]_i_1_n_0 ;
  wire \bank02/grn22/grn[12]_i_1_n_0 ;
  wire \bank02/grn22/grn[13]_i_1_n_0 ;
  wire \bank02/grn22/grn[14]_i_1_n_0 ;
  wire \bank02/grn22/grn[15]_i_2_n_0 ;
  wire \bank02/grn22/grn[1]_i_1_n_0 ;
  wire \bank02/grn22/grn[2]_i_1_n_0 ;
  wire \bank02/grn22/grn[3]_i_1_n_0 ;
  wire \bank02/grn22/grn[4]_i_1_n_0 ;
  wire \bank02/grn22/grn[5]_i_1_n_0 ;
  wire \bank02/grn22/grn[6]_i_1_n_0 ;
  wire \bank02/grn22/grn[7]_i_1_n_0 ;
  wire \bank02/grn22/grn[8]_i_1_n_0 ;
  wire \bank02/grn22/grn[9]_i_1_n_0 ;
  wire \bank02/grn23/grn[0]_i_1_n_0 ;
  wire \bank02/grn23/grn[10]_i_1_n_0 ;
  wire \bank02/grn23/grn[11]_i_1_n_0 ;
  wire \bank02/grn23/grn[12]_i_1_n_0 ;
  wire \bank02/grn23/grn[13]_i_1_n_0 ;
  wire \bank02/grn23/grn[14]_i_1_n_0 ;
  wire \bank02/grn23/grn[15]_i_2_n_0 ;
  wire \bank02/grn23/grn[1]_i_1_n_0 ;
  wire \bank02/grn23/grn[2]_i_1_n_0 ;
  wire \bank02/grn23/grn[3]_i_1_n_0 ;
  wire \bank02/grn23/grn[4]_i_1_n_0 ;
  wire \bank02/grn23/grn[5]_i_1_n_0 ;
  wire \bank02/grn23/grn[6]_i_1_n_0 ;
  wire \bank02/grn23/grn[7]_i_1_n_0 ;
  wire \bank02/grn23/grn[8]_i_1_n_0 ;
  wire \bank02/grn23/grn[9]_i_1_n_0 ;
  wire \bank02/grn24/grn[0]_i_1_n_0 ;
  wire \bank02/grn24/grn[10]_i_1_n_0 ;
  wire \bank02/grn24/grn[11]_i_1_n_0 ;
  wire \bank02/grn24/grn[12]_i_1_n_0 ;
  wire \bank02/grn24/grn[13]_i_1_n_0 ;
  wire \bank02/grn24/grn[14]_i_1_n_0 ;
  wire \bank02/grn24/grn[15]_i_2_n_0 ;
  wire \bank02/grn24/grn[1]_i_1_n_0 ;
  wire \bank02/grn24/grn[2]_i_1_n_0 ;
  wire \bank02/grn24/grn[3]_i_1_n_0 ;
  wire \bank02/grn24/grn[4]_i_1_n_0 ;
  wire \bank02/grn24/grn[5]_i_1_n_0 ;
  wire \bank02/grn24/grn[6]_i_1_n_0 ;
  wire \bank02/grn24/grn[7]_i_1_n_0 ;
  wire \bank02/grn24/grn[8]_i_1_n_0 ;
  wire \bank02/grn24/grn[9]_i_1_n_0 ;
  wire \bank02/grn25/grn[0]_i_1_n_0 ;
  wire \bank02/grn25/grn[10]_i_1_n_0 ;
  wire \bank02/grn25/grn[11]_i_1_n_0 ;
  wire \bank02/grn25/grn[12]_i_1_n_0 ;
  wire \bank02/grn25/grn[13]_i_1_n_0 ;
  wire \bank02/grn25/grn[14]_i_1_n_0 ;
  wire \bank02/grn25/grn[15]_i_2_n_0 ;
  wire \bank02/grn25/grn[1]_i_1_n_0 ;
  wire \bank02/grn25/grn[2]_i_1_n_0 ;
  wire \bank02/grn25/grn[3]_i_1_n_0 ;
  wire \bank02/grn25/grn[4]_i_1_n_0 ;
  wire \bank02/grn25/grn[5]_i_1_n_0 ;
  wire \bank02/grn25/grn[6]_i_1_n_0 ;
  wire \bank02/grn25/grn[7]_i_1_n_0 ;
  wire \bank02/grn25/grn[8]_i_1_n_0 ;
  wire \bank02/grn25/grn[9]_i_1_n_0 ;
  wire \bank02/grn26/grn[0]_i_1_n_0 ;
  wire \bank02/grn26/grn[10]_i_1_n_0 ;
  wire \bank02/grn26/grn[11]_i_1_n_0 ;
  wire \bank02/grn26/grn[12]_i_1_n_0 ;
  wire \bank02/grn26/grn[13]_i_1_n_0 ;
  wire \bank02/grn26/grn[14]_i_1_n_0 ;
  wire \bank02/grn26/grn[15]_i_2_n_0 ;
  wire \bank02/grn26/grn[1]_i_1_n_0 ;
  wire \bank02/grn26/grn[2]_i_1_n_0 ;
  wire \bank02/grn26/grn[3]_i_1_n_0 ;
  wire \bank02/grn26/grn[4]_i_1_n_0 ;
  wire \bank02/grn26/grn[5]_i_1_n_0 ;
  wire \bank02/grn26/grn[6]_i_1_n_0 ;
  wire \bank02/grn26/grn[7]_i_1_n_0 ;
  wire \bank02/grn26/grn[8]_i_1_n_0 ;
  wire \bank02/grn26/grn[9]_i_1_n_0 ;
  wire \bank02/grn27/grn[0]_i_1_n_0 ;
  wire \bank02/grn27/grn[10]_i_1_n_0 ;
  wire \bank02/grn27/grn[11]_i_1_n_0 ;
  wire \bank02/grn27/grn[12]_i_1_n_0 ;
  wire \bank02/grn27/grn[13]_i_1_n_0 ;
  wire \bank02/grn27/grn[14]_i_1_n_0 ;
  wire \bank02/grn27/grn[15]_i_2_n_0 ;
  wire \bank02/grn27/grn[1]_i_1_n_0 ;
  wire \bank02/grn27/grn[2]_i_1_n_0 ;
  wire \bank02/grn27/grn[3]_i_1_n_0 ;
  wire \bank02/grn27/grn[4]_i_1_n_0 ;
  wire \bank02/grn27/grn[5]_i_1_n_0 ;
  wire \bank02/grn27/grn[6]_i_1_n_0 ;
  wire \bank02/grn27/grn[7]_i_1_n_0 ;
  wire \bank02/grn27/grn[8]_i_1_n_0 ;
  wire \bank02/grn27/grn[9]_i_1_n_0 ;
  wire \bank13/a0buso/gr0_bus1 ;
  wire \bank13/a0buso/gr1_bus1 ;
  wire \bank13/a0buso/gr2_bus1 ;
  wire \bank13/a0buso/gr3_bus1 ;
  wire \bank13/a0buso/gr4_bus1 ;
  wire \bank13/a0buso/gr5_bus1 ;
  wire \bank13/a0buso/gr6_bus1 ;
  wire \bank13/a0buso/gr7_bus1 ;
  wire \bank13/a0buso2l/gr0_bus1 ;
  wire \bank13/a0buso2l/gr3_bus1 ;
  wire \bank13/a0buso2l/gr4_bus1 ;
  wire \bank13/a0buso2l/gr7_bus1 ;
  wire \bank13/a1buso/gr0_bus1 ;
  wire \bank13/a1buso/gr1_bus1 ;
  wire \bank13/a1buso/gr2_bus1 ;
  wire \bank13/a1buso/gr3_bus1 ;
  wire \bank13/a1buso/gr4_bus1 ;
  wire \bank13/a1buso/gr5_bus1 ;
  wire \bank13/a1buso/gr6_bus1 ;
  wire \bank13/a1buso/gr7_bus1 ;
  wire \bank13/a1buso2l/gr0_bus1 ;
  wire \bank13/a1buso2l/gr3_bus1 ;
  wire \bank13/a1buso2l/gr4_bus1 ;
  wire \bank13/a1buso2l/gr7_bus1 ;
  wire \bank13/b0buso/gr0_bus1 ;
  wire \bank13/b0buso/gr1_bus1 ;
  wire \bank13/b0buso/gr2_bus1 ;
  wire \bank13/b0buso/gr3_bus1 ;
  wire \bank13/b0buso/gr4_bus1 ;
  wire \bank13/b0buso/gr5_bus1 ;
  wire \bank13/b0buso/gr6_bus1 ;
  wire \bank13/b0buso/gr7_bus1 ;
  wire \bank13/b0buso2l/gr0_bus1 ;
  wire \bank13/b0buso2l/gr1_bus1 ;
  wire \bank13/b0buso2l/gr2_bus1 ;
  wire \bank13/b0buso2l/gr3_bus1 ;
  wire \bank13/b0buso2l/gr4_bus1 ;
  wire \bank13/b0buso2l/gr5_bus1 ;
  wire \bank13/b0buso2l/gr6_bus1 ;
  wire \bank13/b0buso2l/gr7_bus1 ;
  wire \bank13/b1buso/gr0_bus1 ;
  wire \bank13/b1buso/gr1_bus1 ;
  wire \bank13/b1buso/gr2_bus1 ;
  wire \bank13/b1buso/gr3_bus1 ;
  wire \bank13/b1buso/gr4_bus1 ;
  wire \bank13/b1buso/gr5_bus1 ;
  wire \bank13/b1buso/gr6_bus1 ;
  wire \bank13/b1buso/gr7_bus1 ;
  wire \bank13/b1buso2l/gr0_bus1 ;
  wire \bank13/b1buso2l/gr1_bus1 ;
  wire \bank13/b1buso2l/gr2_bus1 ;
  wire \bank13/b1buso2l/gr3_bus1 ;
  wire \bank13/b1buso2l/gr4_bus1 ;
  wire \bank13/b1buso2l/gr5_bus1 ;
  wire \bank13/b1buso2l/gr6_bus1 ;
  wire \bank13/b1buso2l/gr7_bus1 ;
  wire \bank13/grn00/grn[0]_i_1_n_0 ;
  wire \bank13/grn00/grn[10]_i_1_n_0 ;
  wire \bank13/grn00/grn[11]_i_1_n_0 ;
  wire \bank13/grn00/grn[12]_i_1_n_0 ;
  wire \bank13/grn00/grn[13]_i_1_n_0 ;
  wire \bank13/grn00/grn[14]_i_1_n_0 ;
  wire \bank13/grn00/grn[15]_i_2_n_0 ;
  wire \bank13/grn00/grn[1]_i_1_n_0 ;
  wire \bank13/grn00/grn[2]_i_1_n_0 ;
  wire \bank13/grn00/grn[3]_i_1_n_0 ;
  wire \bank13/grn00/grn[4]_i_1_n_0 ;
  wire \bank13/grn00/grn[5]_i_1_n_0 ;
  wire \bank13/grn00/grn[6]_i_1_n_0 ;
  wire \bank13/grn00/grn[7]_i_1_n_0 ;
  wire \bank13/grn00/grn[8]_i_1_n_0 ;
  wire \bank13/grn00/grn[9]_i_1_n_0 ;
  wire \bank13/grn01/grn[0]_i_1_n_0 ;
  wire \bank13/grn01/grn[10]_i_1_n_0 ;
  wire \bank13/grn01/grn[11]_i_1_n_0 ;
  wire \bank13/grn01/grn[12]_i_1_n_0 ;
  wire \bank13/grn01/grn[13]_i_1_n_0 ;
  wire \bank13/grn01/grn[14]_i_1_n_0 ;
  wire \bank13/grn01/grn[15]_i_2_n_0 ;
  wire \bank13/grn01/grn[1]_i_1_n_0 ;
  wire \bank13/grn01/grn[2]_i_1_n_0 ;
  wire \bank13/grn01/grn[3]_i_1_n_0 ;
  wire \bank13/grn01/grn[4]_i_1_n_0 ;
  wire \bank13/grn01/grn[5]_i_1_n_0 ;
  wire \bank13/grn01/grn[6]_i_1_n_0 ;
  wire \bank13/grn01/grn[7]_i_1_n_0 ;
  wire \bank13/grn01/grn[8]_i_1_n_0 ;
  wire \bank13/grn01/grn[9]_i_1_n_0 ;
  wire \bank13/grn02/grn[0]_i_1_n_0 ;
  wire \bank13/grn02/grn[10]_i_1_n_0 ;
  wire \bank13/grn02/grn[11]_i_1_n_0 ;
  wire \bank13/grn02/grn[12]_i_1_n_0 ;
  wire \bank13/grn02/grn[13]_i_1_n_0 ;
  wire \bank13/grn02/grn[14]_i_1_n_0 ;
  wire \bank13/grn02/grn[15]_i_2_n_0 ;
  wire \bank13/grn02/grn[1]_i_1_n_0 ;
  wire \bank13/grn02/grn[2]_i_1_n_0 ;
  wire \bank13/grn02/grn[3]_i_1_n_0 ;
  wire \bank13/grn02/grn[4]_i_1_n_0 ;
  wire \bank13/grn02/grn[5]_i_1_n_0 ;
  wire \bank13/grn02/grn[6]_i_1_n_0 ;
  wire \bank13/grn02/grn[7]_i_1_n_0 ;
  wire \bank13/grn02/grn[8]_i_1_n_0 ;
  wire \bank13/grn02/grn[9]_i_1_n_0 ;
  wire \bank13/grn03/grn[0]_i_1_n_0 ;
  wire \bank13/grn03/grn[10]_i_1_n_0 ;
  wire \bank13/grn03/grn[11]_i_1_n_0 ;
  wire \bank13/grn03/grn[12]_i_1_n_0 ;
  wire \bank13/grn03/grn[13]_i_1_n_0 ;
  wire \bank13/grn03/grn[14]_i_1_n_0 ;
  wire \bank13/grn03/grn[15]_i_2_n_0 ;
  wire \bank13/grn03/grn[1]_i_1_n_0 ;
  wire \bank13/grn03/grn[2]_i_1_n_0 ;
  wire \bank13/grn03/grn[3]_i_1_n_0 ;
  wire \bank13/grn03/grn[4]_i_1_n_0 ;
  wire \bank13/grn03/grn[5]_i_1_n_0 ;
  wire \bank13/grn03/grn[6]_i_1_n_0 ;
  wire \bank13/grn03/grn[7]_i_1_n_0 ;
  wire \bank13/grn03/grn[8]_i_1_n_0 ;
  wire \bank13/grn03/grn[9]_i_1_n_0 ;
  wire \bank13/grn04/grn[0]_i_1_n_0 ;
  wire \bank13/grn04/grn[10]_i_1_n_0 ;
  wire \bank13/grn04/grn[11]_i_1_n_0 ;
  wire \bank13/grn04/grn[12]_i_1_n_0 ;
  wire \bank13/grn04/grn[13]_i_1_n_0 ;
  wire \bank13/grn04/grn[14]_i_1_n_0 ;
  wire \bank13/grn04/grn[15]_i_2_n_0 ;
  wire \bank13/grn04/grn[1]_i_1_n_0 ;
  wire \bank13/grn04/grn[2]_i_1_n_0 ;
  wire \bank13/grn04/grn[3]_i_1_n_0 ;
  wire \bank13/grn04/grn[4]_i_1_n_0 ;
  wire \bank13/grn04/grn[5]_i_1_n_0 ;
  wire \bank13/grn04/grn[6]_i_1_n_0 ;
  wire \bank13/grn04/grn[7]_i_1_n_0 ;
  wire \bank13/grn04/grn[8]_i_1_n_0 ;
  wire \bank13/grn04/grn[9]_i_1_n_0 ;
  wire \bank13/grn05/grn[0]_i_1_n_0 ;
  wire \bank13/grn05/grn[10]_i_1_n_0 ;
  wire \bank13/grn05/grn[11]_i_1_n_0 ;
  wire \bank13/grn05/grn[12]_i_1_n_0 ;
  wire \bank13/grn05/grn[13]_i_1_n_0 ;
  wire \bank13/grn05/grn[14]_i_1_n_0 ;
  wire \bank13/grn05/grn[15]_i_2_n_0 ;
  wire \bank13/grn05/grn[1]_i_1_n_0 ;
  wire \bank13/grn05/grn[2]_i_1_n_0 ;
  wire \bank13/grn05/grn[3]_i_1_n_0 ;
  wire \bank13/grn05/grn[4]_i_1_n_0 ;
  wire \bank13/grn05/grn[5]_i_1_n_0 ;
  wire \bank13/grn05/grn[6]_i_1_n_0 ;
  wire \bank13/grn05/grn[7]_i_1_n_0 ;
  wire \bank13/grn05/grn[8]_i_1_n_0 ;
  wire \bank13/grn05/grn[9]_i_1_n_0 ;
  wire \bank13/grn06/grn[0]_i_1_n_0 ;
  wire \bank13/grn06/grn[10]_i_1_n_0 ;
  wire \bank13/grn06/grn[11]_i_1_n_0 ;
  wire \bank13/grn06/grn[12]_i_1_n_0 ;
  wire \bank13/grn06/grn[13]_i_1_n_0 ;
  wire \bank13/grn06/grn[14]_i_1_n_0 ;
  wire \bank13/grn06/grn[15]_i_2_n_0 ;
  wire \bank13/grn06/grn[1]_i_1_n_0 ;
  wire \bank13/grn06/grn[2]_i_1_n_0 ;
  wire \bank13/grn06/grn[3]_i_1_n_0 ;
  wire \bank13/grn06/grn[4]_i_1_n_0 ;
  wire \bank13/grn06/grn[5]_i_1_n_0 ;
  wire \bank13/grn06/grn[6]_i_1_n_0 ;
  wire \bank13/grn06/grn[7]_i_1_n_0 ;
  wire \bank13/grn06/grn[8]_i_1_n_0 ;
  wire \bank13/grn06/grn[9]_i_1_n_0 ;
  wire \bank13/grn07/grn[0]_i_1_n_0 ;
  wire \bank13/grn07/grn[10]_i_1_n_0 ;
  wire \bank13/grn07/grn[11]_i_1_n_0 ;
  wire \bank13/grn07/grn[12]_i_1_n_0 ;
  wire \bank13/grn07/grn[13]_i_1_n_0 ;
  wire \bank13/grn07/grn[14]_i_1_n_0 ;
  wire \bank13/grn07/grn[15]_i_2_n_0 ;
  wire \bank13/grn07/grn[1]_i_1_n_0 ;
  wire \bank13/grn07/grn[2]_i_1_n_0 ;
  wire \bank13/grn07/grn[3]_i_1_n_0 ;
  wire \bank13/grn07/grn[4]_i_1_n_0 ;
  wire \bank13/grn07/grn[5]_i_1_n_0 ;
  wire \bank13/grn07/grn[6]_i_1_n_0 ;
  wire \bank13/grn07/grn[7]_i_1_n_0 ;
  wire \bank13/grn07/grn[8]_i_1_n_0 ;
  wire \bank13/grn07/grn[9]_i_1_n_0 ;
  wire \bank13/grn20/grn[0]_i_1_n_0 ;
  wire \bank13/grn20/grn[10]_i_1_n_0 ;
  wire \bank13/grn20/grn[11]_i_1_n_0 ;
  wire \bank13/grn20/grn[12]_i_1_n_0 ;
  wire \bank13/grn20/grn[13]_i_1_n_0 ;
  wire \bank13/grn20/grn[14]_i_1_n_0 ;
  wire \bank13/grn20/grn[15]_i_2_n_0 ;
  wire \bank13/grn20/grn[1]_i_1_n_0 ;
  wire \bank13/grn20/grn[2]_i_1_n_0 ;
  wire \bank13/grn20/grn[3]_i_1_n_0 ;
  wire \bank13/grn20/grn[4]_i_1_n_0 ;
  wire \bank13/grn20/grn[5]_i_1_n_0 ;
  wire \bank13/grn20/grn[6]_i_1_n_0 ;
  wire \bank13/grn20/grn[7]_i_1_n_0 ;
  wire \bank13/grn20/grn[8]_i_1_n_0 ;
  wire \bank13/grn20/grn[9]_i_1_n_0 ;
  wire \bank13/grn21/grn[0]_i_1_n_0 ;
  wire \bank13/grn21/grn[10]_i_1_n_0 ;
  wire \bank13/grn21/grn[11]_i_1_n_0 ;
  wire \bank13/grn21/grn[12]_i_1_n_0 ;
  wire \bank13/grn21/grn[13]_i_1_n_0 ;
  wire \bank13/grn21/grn[14]_i_1_n_0 ;
  wire \bank13/grn21/grn[15]_i_2_n_0 ;
  wire \bank13/grn21/grn[1]_i_1_n_0 ;
  wire \bank13/grn21/grn[2]_i_1_n_0 ;
  wire \bank13/grn21/grn[3]_i_1_n_0 ;
  wire \bank13/grn21/grn[4]_i_1_n_0 ;
  wire \bank13/grn21/grn[5]_i_1_n_0 ;
  wire \bank13/grn21/grn[6]_i_1_n_0 ;
  wire \bank13/grn21/grn[7]_i_1_n_0 ;
  wire \bank13/grn21/grn[8]_i_1_n_0 ;
  wire \bank13/grn21/grn[9]_i_1_n_0 ;
  wire \bank13/grn22/grn[0]_i_1_n_0 ;
  wire \bank13/grn22/grn[10]_i_1_n_0 ;
  wire \bank13/grn22/grn[11]_i_1_n_0 ;
  wire \bank13/grn22/grn[12]_i_1_n_0 ;
  wire \bank13/grn22/grn[13]_i_1_n_0 ;
  wire \bank13/grn22/grn[14]_i_1_n_0 ;
  wire \bank13/grn22/grn[15]_i_2_n_0 ;
  wire \bank13/grn22/grn[1]_i_1_n_0 ;
  wire \bank13/grn22/grn[2]_i_1_n_0 ;
  wire \bank13/grn22/grn[3]_i_1_n_0 ;
  wire \bank13/grn22/grn[4]_i_1_n_0 ;
  wire \bank13/grn22/grn[5]_i_1_n_0 ;
  wire \bank13/grn22/grn[6]_i_1_n_0 ;
  wire \bank13/grn22/grn[7]_i_1_n_0 ;
  wire \bank13/grn22/grn[8]_i_1_n_0 ;
  wire \bank13/grn22/grn[9]_i_1_n_0 ;
  wire \bank13/grn23/grn[0]_i_1_n_0 ;
  wire \bank13/grn23/grn[10]_i_1_n_0 ;
  wire \bank13/grn23/grn[11]_i_1_n_0 ;
  wire \bank13/grn23/grn[12]_i_1_n_0 ;
  wire \bank13/grn23/grn[13]_i_1_n_0 ;
  wire \bank13/grn23/grn[14]_i_1_n_0 ;
  wire \bank13/grn23/grn[15]_i_2_n_0 ;
  wire \bank13/grn23/grn[1]_i_1_n_0 ;
  wire \bank13/grn23/grn[2]_i_1_n_0 ;
  wire \bank13/grn23/grn[3]_i_1_n_0 ;
  wire \bank13/grn23/grn[4]_i_1_n_0 ;
  wire \bank13/grn23/grn[5]_i_1_n_0 ;
  wire \bank13/grn23/grn[6]_i_1_n_0 ;
  wire \bank13/grn23/grn[7]_i_1_n_0 ;
  wire \bank13/grn23/grn[8]_i_1_n_0 ;
  wire \bank13/grn23/grn[9]_i_1_n_0 ;
  wire \bank13/grn24/grn[0]_i_1_n_0 ;
  wire \bank13/grn24/grn[10]_i_1_n_0 ;
  wire \bank13/grn24/grn[11]_i_1_n_0 ;
  wire \bank13/grn24/grn[12]_i_1_n_0 ;
  wire \bank13/grn24/grn[13]_i_1_n_0 ;
  wire \bank13/grn24/grn[14]_i_1_n_0 ;
  wire \bank13/grn24/grn[15]_i_2_n_0 ;
  wire \bank13/grn24/grn[1]_i_1_n_0 ;
  wire \bank13/grn24/grn[2]_i_1_n_0 ;
  wire \bank13/grn24/grn[3]_i_1_n_0 ;
  wire \bank13/grn24/grn[4]_i_1_n_0 ;
  wire \bank13/grn24/grn[5]_i_1_n_0 ;
  wire \bank13/grn24/grn[6]_i_1_n_0 ;
  wire \bank13/grn24/grn[7]_i_1_n_0 ;
  wire \bank13/grn24/grn[8]_i_1_n_0 ;
  wire \bank13/grn24/grn[9]_i_1_n_0 ;
  wire \bank13/grn25/grn[0]_i_1_n_0 ;
  wire \bank13/grn25/grn[10]_i_1_n_0 ;
  wire \bank13/grn25/grn[11]_i_1_n_0 ;
  wire \bank13/grn25/grn[12]_i_1_n_0 ;
  wire \bank13/grn25/grn[13]_i_1_n_0 ;
  wire \bank13/grn25/grn[14]_i_1_n_0 ;
  wire \bank13/grn25/grn[15]_i_2_n_0 ;
  wire \bank13/grn25/grn[1]_i_1_n_0 ;
  wire \bank13/grn25/grn[2]_i_1_n_0 ;
  wire \bank13/grn25/grn[3]_i_1_n_0 ;
  wire \bank13/grn25/grn[4]_i_1_n_0 ;
  wire \bank13/grn25/grn[5]_i_1_n_0 ;
  wire \bank13/grn25/grn[6]_i_1_n_0 ;
  wire \bank13/grn25/grn[7]_i_1_n_0 ;
  wire \bank13/grn25/grn[8]_i_1_n_0 ;
  wire \bank13/grn25/grn[9]_i_1_n_0 ;
  wire \bank13/grn26/grn[0]_i_1_n_0 ;
  wire \bank13/grn26/grn[10]_i_1_n_0 ;
  wire \bank13/grn26/grn[11]_i_1_n_0 ;
  wire \bank13/grn26/grn[12]_i_1_n_0 ;
  wire \bank13/grn26/grn[13]_i_1_n_0 ;
  wire \bank13/grn26/grn[14]_i_1_n_0 ;
  wire \bank13/grn26/grn[15]_i_2_n_0 ;
  wire \bank13/grn26/grn[1]_i_1_n_0 ;
  wire \bank13/grn26/grn[2]_i_1_n_0 ;
  wire \bank13/grn26/grn[3]_i_1_n_0 ;
  wire \bank13/grn26/grn[4]_i_1_n_0 ;
  wire \bank13/grn26/grn[5]_i_1_n_0 ;
  wire \bank13/grn26/grn[6]_i_1_n_0 ;
  wire \bank13/grn26/grn[7]_i_1_n_0 ;
  wire \bank13/grn26/grn[8]_i_1_n_0 ;
  wire \bank13/grn26/grn[9]_i_1_n_0 ;
  wire \bank13/grn27/grn[0]_i_1_n_0 ;
  wire \bank13/grn27/grn[10]_i_1_n_0 ;
  wire \bank13/grn27/grn[11]_i_1_n_0 ;
  wire \bank13/grn27/grn[12]_i_1_n_0 ;
  wire \bank13/grn27/grn[13]_i_1_n_0 ;
  wire \bank13/grn27/grn[14]_i_1_n_0 ;
  wire \bank13/grn27/grn[15]_i_2_n_0 ;
  wire \bank13/grn27/grn[1]_i_1_n_0 ;
  wire \bank13/grn27/grn[2]_i_1_n_0 ;
  wire \bank13/grn27/grn[3]_i_1_n_0 ;
  wire \bank13/grn27/grn[4]_i_1_n_0 ;
  wire \bank13/grn27/grn[5]_i_1_n_0 ;
  wire \bank13/grn27/grn[6]_i_1_n_0 ;
  wire \bank13/grn27/grn[7]_i_1_n_0 ;
  wire \bank13/grn27/grn[8]_i_1_n_0 ;
  wire \bank13/grn27/grn[9]_i_1_n_0 ;
  wire [15:0]bbus_o;
  wire \bbus_o[0]_INST_0_i_15_n_0 ;
  wire \bbus_o[0]_INST_0_i_1_n_0 ;
  wire \bbus_o[0]_INST_0_i_23_n_0 ;
  wire \bbus_o[0]_INST_0_i_24_n_0 ;
  wire \bbus_o[0]_INST_0_i_2_n_0 ;
  wire \bbus_o[0]_INST_0_i_3_n_0 ;
  wire \bbus_o[0]_INST_0_i_8_n_0 ;
  wire \bbus_o[1]_INST_0_i_14_n_0 ;
  wire \bbus_o[1]_INST_0_i_1_n_0 ;
  wire \bbus_o[1]_INST_0_i_22_n_0 ;
  wire \bbus_o[1]_INST_0_i_23_n_0 ;
  wire \bbus_o[1]_INST_0_i_2_n_0 ;
  wire \bbus_o[1]_INST_0_i_7_n_0 ;
  wire \bbus_o[2]_INST_0_i_15_n_0 ;
  wire \bbus_o[2]_INST_0_i_1_n_0 ;
  wire \bbus_o[2]_INST_0_i_23_n_0 ;
  wire \bbus_o[2]_INST_0_i_24_n_0 ;
  wire \bbus_o[2]_INST_0_i_2_n_0 ;
  wire \bbus_o[2]_INST_0_i_3_n_0 ;
  wire \bbus_o[2]_INST_0_i_8_n_0 ;
  wire \bbus_o[3]_INST_0_i_15_n_0 ;
  wire \bbus_o[3]_INST_0_i_1_n_0 ;
  wire \bbus_o[3]_INST_0_i_23_n_0 ;
  wire \bbus_o[3]_INST_0_i_24_n_0 ;
  wire \bbus_o[3]_INST_0_i_2_n_0 ;
  wire \bbus_o[3]_INST_0_i_3_n_0 ;
  wire \bbus_o[3]_INST_0_i_8_n_0 ;
  wire \bbus_o[4]_INST_0_i_15_n_0 ;
  wire \bbus_o[4]_INST_0_i_1_n_0 ;
  wire \bbus_o[4]_INST_0_i_26_n_0 ;
  wire \bbus_o[4]_INST_0_i_28_n_0 ;
  wire \bbus_o[4]_INST_0_i_2_n_0 ;
  wire \bbus_o[4]_INST_0_i_3_n_0 ;
  wire \bbus_o[4]_INST_0_i_8_n_0 ;
  wire \bbus_o[5]_INST_0_i_18_n_0 ;
  wire \bbus_o[5]_INST_0_i_1_n_0 ;
  wire \bbus_o[5]_INST_0_i_2_n_0 ;
  wire \bbus_o[5]_INST_0_i_3_n_0 ;
  wire \bbus_o[5]_INST_0_i_8_n_0 ;
  wire \bbus_o[6]_INST_0_i_18_n_0 ;
  wire \bbus_o[6]_INST_0_i_1_n_0 ;
  wire \bbus_o[6]_INST_0_i_2_n_0 ;
  wire \bbus_o[6]_INST_0_i_3_n_0 ;
  wire \bbus_o[6]_INST_0_i_8_n_0 ;
  wire \bbus_o[7]_INST_0_i_18_n_0 ;
  wire \bbus_o[7]_INST_0_i_1_n_0 ;
  wire \bbus_o[7]_INST_0_i_2_n_0 ;
  wire \bbus_o[7]_INST_0_i_3_n_0 ;
  wire \bbus_o[7]_INST_0_i_8_n_0 ;
  wire [2:0]bcmd;
  wire \bcmd[0]_INST_0_i_10_n_0 ;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_13_n_0 ;
  wire \bcmd[0]_INST_0_i_14_n_0 ;
  wire \bcmd[0]_INST_0_i_15_n_0 ;
  wire \bcmd[0]_INST_0_i_16_n_0 ;
  wire \bcmd[0]_INST_0_i_17_n_0 ;
  wire \bcmd[0]_INST_0_i_18_n_0 ;
  wire \bcmd[0]_INST_0_i_19_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_20_n_0 ;
  wire \bcmd[0]_INST_0_i_21_n_0 ;
  wire \bcmd[0]_INST_0_i_22_n_0 ;
  wire \bcmd[0]_INST_0_i_23_n_0 ;
  wire \bcmd[0]_INST_0_i_24_n_0 ;
  wire \bcmd[0]_INST_0_i_25_n_0 ;
  wire \bcmd[0]_INST_0_i_26_n_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_3_n_0 ;
  wire \bcmd[0]_INST_0_i_4_n_0 ;
  wire \bcmd[0]_INST_0_i_5_n_0 ;
  wire \bcmd[0]_INST_0_i_6_n_0 ;
  wire \bcmd[0]_INST_0_i_7_n_0 ;
  wire \bcmd[0]_INST_0_i_8_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_11_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_14_n_0 ;
  wire \bcmd[1]_INST_0_i_15_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_17_n_0 ;
  wire \bcmd[1]_INST_0_i_18_n_0 ;
  wire \bcmd[1]_INST_0_i_19_n_0 ;
  wire \bcmd[1]_INST_0_i_1_n_0 ;
  wire \bcmd[1]_INST_0_i_2_n_0 ;
  wire \bcmd[1]_INST_0_i_3_n_0 ;
  wire \bcmd[1]_INST_0_i_4_n_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_6_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_8_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2]_INST_0_i_1_n_0 ;
  wire \bcmd[2]_INST_0_i_2_n_0 ;
  wire \bcmd[2]_INST_0_i_3_n_0 ;
  wire \bcmd[2]_INST_0_i_4_n_0 ;
  wire \bcmd[2]_INST_0_i_5_n_0 ;
  wire \bcmd[2]_INST_0_i_6_n_0 ;
  wire \bcmd[2]_INST_0_i_7_n_0 ;
  wire [15:0]bdatr;
  wire [15:0]bdatw;
  wire \bdatw[10]_INST_0_i_14_n_0 ;
  wire \bdatw[10]_INST_0_i_15_n_0 ;
  wire \bdatw[10]_INST_0_i_1_n_0 ;
  wire \bdatw[10]_INST_0_i_22_n_0 ;
  wire \bdatw[10]_INST_0_i_2_n_0 ;
  wire \bdatw[10]_INST_0_i_32_n_0 ;
  wire \bdatw[10]_INST_0_i_33_n_0 ;
  wire \bdatw[10]_INST_0_i_34_n_0 ;
  wire \bdatw[10]_INST_0_i_3_n_0 ;
  wire \bdatw[10]_INST_0_i_4_n_0 ;
  wire \bdatw[10]_INST_0_i_53_n_0 ;
  wire \bdatw[10]_INST_0_i_5_n_0 ;
  wire \bdatw[10]_INST_0_i_67_n_0 ;
  wire \bdatw[10]_INST_0_i_72_n_0 ;
  wire \bdatw[10]_INST_0_i_73_n_0 ;
  wire \bdatw[10]_INST_0_i_74_n_0 ;
  wire \bdatw[10]_INST_0_i_75_n_0 ;
  wire \bdatw[10]_INST_0_i_76_n_0 ;
  wire \bdatw[10]_INST_0_i_77_n_0 ;
  wire \bdatw[10]_INST_0_i_78_n_0 ;
  wire \bdatw[10]_INST_0_i_79_n_0 ;
  wire \bdatw[10]_INST_0_i_8_n_0 ;
  wire \bdatw[10]_INST_0_i_9_n_0 ;
  wire \bdatw[11]_INST_0_i_10_n_0 ;
  wire \bdatw[11]_INST_0_i_11_n_0 ;
  wire \bdatw[11]_INST_0_i_16_n_0 ;
  wire \bdatw[11]_INST_0_i_1_n_0 ;
  wire \bdatw[11]_INST_0_i_26_n_0 ;
  wire \bdatw[11]_INST_0_i_27_n_0 ;
  wire \bdatw[11]_INST_0_i_28_n_0 ;
  wire \bdatw[11]_INST_0_i_2_n_0 ;
  wire \bdatw[11]_INST_0_i_38_n_0 ;
  wire \bdatw[11]_INST_0_i_39_n_0 ;
  wire \bdatw[11]_INST_0_i_3_n_0 ;
  wire \bdatw[11]_INST_0_i_40_n_0 ;
  wire \bdatw[11]_INST_0_i_4_n_0 ;
  wire \bdatw[11]_INST_0_i_57_n_0 ;
  wire \bdatw[11]_INST_0_i_5_n_0 ;
  wire \bdatw[11]_INST_0_i_71_n_0 ;
  wire \bdatw[11]_INST_0_i_72_n_0 ;
  wire \bdatw[11]_INST_0_i_73_n_0 ;
  wire \bdatw[11]_INST_0_i_74_n_0 ;
  wire \bdatw[11]_INST_0_i_75_n_0 ;
  wire \bdatw[11]_INST_0_i_76_n_0 ;
  wire \bdatw[11]_INST_0_i_77_n_0 ;
  wire \bdatw[11]_INST_0_i_78_n_0 ;
  wire \bdatw[11]_INST_0_i_79_n_0 ;
  wire \bdatw[12]_INST_0_i_10_n_0 ;
  wire \bdatw[12]_INST_0_i_11_n_0 ;
  wire \bdatw[12]_INST_0_i_16_n_0 ;
  wire \bdatw[12]_INST_0_i_17_n_0 ;
  wire \bdatw[12]_INST_0_i_1_n_0 ;
  wire \bdatw[12]_INST_0_i_27_n_0 ;
  wire \bdatw[12]_INST_0_i_2_n_0 ;
  wire \bdatw[12]_INST_0_i_37_n_0 ;
  wire \bdatw[12]_INST_0_i_38_n_0 ;
  wire \bdatw[12]_INST_0_i_39_n_0 ;
  wire \bdatw[12]_INST_0_i_3_n_0 ;
  wire \bdatw[12]_INST_0_i_4_n_0 ;
  wire \bdatw[12]_INST_0_i_56_n_0 ;
  wire \bdatw[12]_INST_0_i_5_n_0 ;
  wire \bdatw[12]_INST_0_i_70_n_0 ;
  wire \bdatw[12]_INST_0_i_71_n_0 ;
  wire \bdatw[12]_INST_0_i_72_n_0 ;
  wire \bdatw[12]_INST_0_i_73_n_0 ;
  wire \bdatw[12]_INST_0_i_74_n_0 ;
  wire \bdatw[12]_INST_0_i_75_n_0 ;
  wire \bdatw[12]_INST_0_i_76_n_0 ;
  wire \bdatw[12]_INST_0_i_77_n_0 ;
  wire \bdatw[12]_INST_0_i_78_n_0 ;
  wire \bdatw[12]_INST_0_i_79_n_0 ;
  wire \bdatw[12]_INST_0_i_80_n_0 ;
  wire \bdatw[12]_INST_0_i_81_n_0 ;
  wire \bdatw[12]_INST_0_i_82_n_0 ;
  wire \bdatw[12]_INST_0_i_83_n_0 ;
  wire \bdatw[12]_INST_0_i_84_n_0 ;
  wire \bdatw[12]_INST_0_i_85_n_0 ;
  wire \bdatw[12]_INST_0_i_86_n_0 ;
  wire \bdatw[12]_INST_0_i_87_n_0 ;
  wire \bdatw[12]_INST_0_i_88_n_0 ;
  wire \bdatw[12]_INST_0_i_89_n_0 ;
  wire \bdatw[12]_INST_0_i_90_n_0 ;
  wire \bdatw[12]_INST_0_i_91_n_0 ;
  wire \bdatw[12]_INST_0_i_92_n_0 ;
  wire \bdatw[12]_INST_0_i_93_n_0 ;
  wire \bdatw[12]_INST_0_i_94_n_0 ;
  wire \bdatw[12]_INST_0_i_95_n_0 ;
  wire \bdatw[12]_INST_0_i_96_n_0 ;
  wire \bdatw[12]_INST_0_i_97_n_0 ;
  wire \bdatw[12]_INST_0_i_98_n_0 ;
  wire \bdatw[13]_INST_0_i_10_n_0 ;
  wire \bdatw[13]_INST_0_i_11_n_0 ;
  wire \bdatw[13]_INST_0_i_16_n_0 ;
  wire \bdatw[13]_INST_0_i_17_n_0 ;
  wire \bdatw[13]_INST_0_i_1_n_0 ;
  wire \bdatw[13]_INST_0_i_27_n_0 ;
  wire \bdatw[13]_INST_0_i_28_n_0 ;
  wire \bdatw[13]_INST_0_i_2_n_0 ;
  wire \bdatw[13]_INST_0_i_38_n_0 ;
  wire \bdatw[13]_INST_0_i_39_n_0 ;
  wire \bdatw[13]_INST_0_i_3_n_0 ;
  wire \bdatw[13]_INST_0_i_40_n_0 ;
  wire \bdatw[13]_INST_0_i_4_n_0 ;
  wire \bdatw[13]_INST_0_i_57_n_0 ;
  wire \bdatw[13]_INST_0_i_5_n_0 ;
  wire \bdatw[13]_INST_0_i_67_n_0 ;
  wire \bdatw[14]_INST_0_i_10_n_0 ;
  wire \bdatw[14]_INST_0_i_11_n_0 ;
  wire \bdatw[14]_INST_0_i_16_n_0 ;
  wire \bdatw[14]_INST_0_i_17_n_0 ;
  wire \bdatw[14]_INST_0_i_18_n_0 ;
  wire \bdatw[14]_INST_0_i_1_n_0 ;
  wire \bdatw[14]_INST_0_i_28_n_0 ;
  wire \bdatw[14]_INST_0_i_29_n_0 ;
  wire \bdatw[14]_INST_0_i_2_n_0 ;
  wire \bdatw[14]_INST_0_i_30_n_0 ;
  wire \bdatw[14]_INST_0_i_3_n_0 ;
  wire \bdatw[14]_INST_0_i_40_n_0 ;
  wire \bdatw[14]_INST_0_i_41_n_0 ;
  wire \bdatw[14]_INST_0_i_42_n_0 ;
  wire \bdatw[14]_INST_0_i_4_n_0 ;
  wire \bdatw[14]_INST_0_i_59_n_0 ;
  wire \bdatw[14]_INST_0_i_5_n_0 ;
  wire \bdatw[14]_INST_0_i_69_n_0 ;
  wire \bdatw[15]_INST_0_i_102_n_0 ;
  wire \bdatw[15]_INST_0_i_103_n_0 ;
  wire \bdatw[15]_INST_0_i_104_n_0 ;
  wire \bdatw[15]_INST_0_i_105_n_0 ;
  wire \bdatw[15]_INST_0_i_106_n_0 ;
  wire \bdatw[15]_INST_0_i_107_n_0 ;
  wire \bdatw[15]_INST_0_i_108_n_0 ;
  wire \bdatw[15]_INST_0_i_112_n_0 ;
  wire \bdatw[15]_INST_0_i_116_n_0 ;
  wire \bdatw[15]_INST_0_i_117_n_0 ;
  wire \bdatw[15]_INST_0_i_123_n_0 ;
  wire \bdatw[15]_INST_0_i_12_n_0 ;
  wire \bdatw[15]_INST_0_i_13_n_0 ;
  wire \bdatw[15]_INST_0_i_142_n_0 ;
  wire \bdatw[15]_INST_0_i_152_n_0 ;
  wire \bdatw[15]_INST_0_i_153_n_0 ;
  wire \bdatw[15]_INST_0_i_154_n_0 ;
  wire \bdatw[15]_INST_0_i_155_n_0 ;
  wire \bdatw[15]_INST_0_i_156_n_0 ;
  wire \bdatw[15]_INST_0_i_157_n_0 ;
  wire \bdatw[15]_INST_0_i_158_n_0 ;
  wire \bdatw[15]_INST_0_i_159_n_0 ;
  wire \bdatw[15]_INST_0_i_160_n_0 ;
  wire \bdatw[15]_INST_0_i_161_n_0 ;
  wire \bdatw[15]_INST_0_i_162_n_0 ;
  wire \bdatw[15]_INST_0_i_163_n_0 ;
  wire \bdatw[15]_INST_0_i_164_n_0 ;
  wire \bdatw[15]_INST_0_i_165_n_0 ;
  wire \bdatw[15]_INST_0_i_166_n_0 ;
  wire \bdatw[15]_INST_0_i_167_n_0 ;
  wire \bdatw[15]_INST_0_i_168_n_0 ;
  wire \bdatw[15]_INST_0_i_169_n_0 ;
  wire \bdatw[15]_INST_0_i_170_n_0 ;
  wire \bdatw[15]_INST_0_i_171_n_0 ;
  wire \bdatw[15]_INST_0_i_172_n_0 ;
  wire \bdatw[15]_INST_0_i_173_n_0 ;
  wire \bdatw[15]_INST_0_i_174_n_0 ;
  wire \bdatw[15]_INST_0_i_175_n_0 ;
  wire \bdatw[15]_INST_0_i_176_n_0 ;
  wire \bdatw[15]_INST_0_i_177_n_0 ;
  wire \bdatw[15]_INST_0_i_178_n_0 ;
  wire \bdatw[15]_INST_0_i_179_n_0 ;
  wire \bdatw[15]_INST_0_i_180_n_0 ;
  wire \bdatw[15]_INST_0_i_181_n_0 ;
  wire \bdatw[15]_INST_0_i_182_n_0 ;
  wire \bdatw[15]_INST_0_i_183_n_0 ;
  wire \bdatw[15]_INST_0_i_184_n_0 ;
  wire \bdatw[15]_INST_0_i_185_n_0 ;
  wire \bdatw[15]_INST_0_i_186_n_0 ;
  wire \bdatw[15]_INST_0_i_187_n_0 ;
  wire \bdatw[15]_INST_0_i_188_n_0 ;
  wire \bdatw[15]_INST_0_i_189_n_0 ;
  wire \bdatw[15]_INST_0_i_18_n_0 ;
  wire \bdatw[15]_INST_0_i_190_n_0 ;
  wire \bdatw[15]_INST_0_i_191_n_0 ;
  wire \bdatw[15]_INST_0_i_192_n_0 ;
  wire \bdatw[15]_INST_0_i_19_n_0 ;
  wire \bdatw[15]_INST_0_i_1_n_0 ;
  wire \bdatw[15]_INST_0_i_202_n_0 ;
  wire \bdatw[15]_INST_0_i_203_n_0 ;
  wire \bdatw[15]_INST_0_i_204_n_0 ;
  wire \bdatw[15]_INST_0_i_205_n_0 ;
  wire \bdatw[15]_INST_0_i_206_n_0 ;
  wire \bdatw[15]_INST_0_i_207_n_0 ;
  wire \bdatw[15]_INST_0_i_208_n_0 ;
  wire \bdatw[15]_INST_0_i_209_n_0 ;
  wire \bdatw[15]_INST_0_i_20_n_0 ;
  wire \bdatw[15]_INST_0_i_210_n_0 ;
  wire \bdatw[15]_INST_0_i_211_n_0 ;
  wire \bdatw[15]_INST_0_i_212_n_0 ;
  wire \bdatw[15]_INST_0_i_213_n_0 ;
  wire \bdatw[15]_INST_0_i_214_n_0 ;
  wire \bdatw[15]_INST_0_i_215_n_0 ;
  wire \bdatw[15]_INST_0_i_216_n_0 ;
  wire \bdatw[15]_INST_0_i_217_n_0 ;
  wire \bdatw[15]_INST_0_i_218_n_0 ;
  wire \bdatw[15]_INST_0_i_219_n_0 ;
  wire \bdatw[15]_INST_0_i_21_n_0 ;
  wire \bdatw[15]_INST_0_i_220_n_0 ;
  wire \bdatw[15]_INST_0_i_221_n_0 ;
  wire \bdatw[15]_INST_0_i_222_n_0 ;
  wire \bdatw[15]_INST_0_i_223_n_0 ;
  wire \bdatw[15]_INST_0_i_224_n_0 ;
  wire \bdatw[15]_INST_0_i_225_n_0 ;
  wire \bdatw[15]_INST_0_i_226_n_0 ;
  wire \bdatw[15]_INST_0_i_227_n_0 ;
  wire \bdatw[15]_INST_0_i_228_n_0 ;
  wire \bdatw[15]_INST_0_i_229_n_0 ;
  wire \bdatw[15]_INST_0_i_22_n_0 ;
  wire \bdatw[15]_INST_0_i_230_n_0 ;
  wire \bdatw[15]_INST_0_i_231_n_0 ;
  wire \bdatw[15]_INST_0_i_232_n_0 ;
  wire \bdatw[15]_INST_0_i_233_n_0 ;
  wire \bdatw[15]_INST_0_i_238_n_0 ;
  wire \bdatw[15]_INST_0_i_253_n_0 ;
  wire \bdatw[15]_INST_0_i_254_n_0 ;
  wire \bdatw[15]_INST_0_i_255_n_0 ;
  wire \bdatw[15]_INST_0_i_256_n_0 ;
  wire \bdatw[15]_INST_0_i_257_n_0 ;
  wire \bdatw[15]_INST_0_i_258_n_0 ;
  wire \bdatw[15]_INST_0_i_259_n_0 ;
  wire \bdatw[15]_INST_0_i_260_n_0 ;
  wire \bdatw[15]_INST_0_i_261_n_0 ;
  wire \bdatw[15]_INST_0_i_262_n_0 ;
  wire \bdatw[15]_INST_0_i_263_n_0 ;
  wire \bdatw[15]_INST_0_i_264_n_0 ;
  wire \bdatw[15]_INST_0_i_265_n_0 ;
  wire \bdatw[15]_INST_0_i_266_n_0 ;
  wire \bdatw[15]_INST_0_i_267_n_0 ;
  wire \bdatw[15]_INST_0_i_268_n_0 ;
  wire \bdatw[15]_INST_0_i_269_n_0 ;
  wire \bdatw[15]_INST_0_i_270_n_0 ;
  wire \bdatw[15]_INST_0_i_271_n_0 ;
  wire \bdatw[15]_INST_0_i_272_n_0 ;
  wire \bdatw[15]_INST_0_i_273_n_0 ;
  wire \bdatw[15]_INST_0_i_274_n_0 ;
  wire \bdatw[15]_INST_0_i_275_n_0 ;
  wire \bdatw[15]_INST_0_i_276_n_0 ;
  wire \bdatw[15]_INST_0_i_277_n_0 ;
  wire \bdatw[15]_INST_0_i_278_n_0 ;
  wire \bdatw[15]_INST_0_i_279_n_0 ;
  wire \bdatw[15]_INST_0_i_280_n_0 ;
  wire \bdatw[15]_INST_0_i_281_n_0 ;
  wire \bdatw[15]_INST_0_i_282_n_0 ;
  wire \bdatw[15]_INST_0_i_283_n_0 ;
  wire \bdatw[15]_INST_0_i_284_n_0 ;
  wire \bdatw[15]_INST_0_i_285_n_0 ;
  wire \bdatw[15]_INST_0_i_286_n_0 ;
  wire \bdatw[15]_INST_0_i_287_n_0 ;
  wire \bdatw[15]_INST_0_i_288_n_0 ;
  wire \bdatw[15]_INST_0_i_289_n_0 ;
  wire \bdatw[15]_INST_0_i_290_n_0 ;
  wire \bdatw[15]_INST_0_i_291_n_0 ;
  wire \bdatw[15]_INST_0_i_292_n_0 ;
  wire \bdatw[15]_INST_0_i_293_n_0 ;
  wire \bdatw[15]_INST_0_i_294_n_0 ;
  wire \bdatw[15]_INST_0_i_295_n_0 ;
  wire \bdatw[15]_INST_0_i_296_n_0 ;
  wire \bdatw[15]_INST_0_i_297_n_0 ;
  wire \bdatw[15]_INST_0_i_298_n_0 ;
  wire \bdatw[15]_INST_0_i_2_n_0 ;
  wire \bdatw[15]_INST_0_i_38_n_0 ;
  wire \bdatw[15]_INST_0_i_39_n_0 ;
  wire \bdatw[15]_INST_0_i_3_n_0 ;
  wire \bdatw[15]_INST_0_i_40_n_0 ;
  wire \bdatw[15]_INST_0_i_41_n_0 ;
  wire \bdatw[15]_INST_0_i_42_n_0 ;
  wire \bdatw[15]_INST_0_i_4_n_0 ;
  wire \bdatw[15]_INST_0_i_59_n_0 ;
  wire \bdatw[15]_INST_0_i_5_n_0 ;
  wire \bdatw[15]_INST_0_i_60_n_0 ;
  wire \bdatw[15]_INST_0_i_61_n_0 ;
  wire \bdatw[15]_INST_0_i_66_n_0 ;
  wire \bdatw[15]_INST_0_i_67_n_0 ;
  wire \bdatw[15]_INST_0_i_68_n_0 ;
  wire \bdatw[15]_INST_0_i_69_n_0 ;
  wire \bdatw[15]_INST_0_i_6_n_0 ;
  wire \bdatw[15]_INST_0_i_70_n_0 ;
  wire \bdatw[15]_INST_0_i_71_n_0 ;
  wire \bdatw[15]_INST_0_i_72_n_0 ;
  wire \bdatw[15]_INST_0_i_73_n_0 ;
  wire \bdatw[15]_INST_0_i_76_n_0 ;
  wire \bdatw[15]_INST_0_i_77_n_0 ;
  wire \bdatw[15]_INST_0_i_7_n_0 ;
  wire \bdatw[15]_INST_0_i_80_n_0 ;
  wire \bdatw[15]_INST_0_i_81_n_0 ;
  wire \bdatw[8]_INST_0_i_14_n_0 ;
  wire \bdatw[8]_INST_0_i_15_n_0 ;
  wire \bdatw[8]_INST_0_i_16_n_0 ;
  wire \bdatw[8]_INST_0_i_17_n_0 ;
  wire \bdatw[8]_INST_0_i_18_n_0 ;
  wire \bdatw[8]_INST_0_i_19_n_0 ;
  wire \bdatw[8]_INST_0_i_1_n_0 ;
  wire \bdatw[8]_INST_0_i_2_n_0 ;
  wire \bdatw[8]_INST_0_i_34_n_0 ;
  wire \bdatw[8]_INST_0_i_35_n_0 ;
  wire \bdatw[8]_INST_0_i_36_n_0 ;
  wire \bdatw[8]_INST_0_i_3_n_0 ;
  wire \bdatw[8]_INST_0_i_41_n_0 ;
  wire \bdatw[8]_INST_0_i_42_n_0 ;
  wire \bdatw[8]_INST_0_i_43_n_0 ;
  wire \bdatw[8]_INST_0_i_44_n_0 ;
  wire \bdatw[8]_INST_0_i_4_n_0 ;
  wire \bdatw[8]_INST_0_i_59_n_0 ;
  wire \bdatw[8]_INST_0_i_5_n_0 ;
  wire \bdatw[8]_INST_0_i_73_n_0 ;
  wire \bdatw[8]_INST_0_i_78_n_0 ;
  wire \bdatw[8]_INST_0_i_79_n_0 ;
  wire \bdatw[8]_INST_0_i_80_n_0 ;
  wire \bdatw[8]_INST_0_i_81_n_0 ;
  wire \bdatw[8]_INST_0_i_82_n_0 ;
  wire \bdatw[8]_INST_0_i_83_n_0 ;
  wire \bdatw[8]_INST_0_i_84_n_0 ;
  wire \bdatw[8]_INST_0_i_85_n_0 ;
  wire \bdatw[8]_INST_0_i_8_n_0 ;
  wire \bdatw[8]_INST_0_i_9_n_0 ;
  wire \bdatw[9]_INST_0_i_13_n_0 ;
  wire \bdatw[9]_INST_0_i_14_n_0 ;
  wire \bdatw[9]_INST_0_i_1_n_0 ;
  wire \bdatw[9]_INST_0_i_20_n_0 ;
  wire \bdatw[9]_INST_0_i_2_n_0 ;
  wire \bdatw[9]_INST_0_i_30_n_0 ;
  wire \bdatw[9]_INST_0_i_31_n_0 ;
  wire \bdatw[9]_INST_0_i_36_n_0 ;
  wire \bdatw[9]_INST_0_i_3_n_0 ;
  wire \bdatw[9]_INST_0_i_4_n_0 ;
  wire \bdatw[9]_INST_0_i_64_n_0 ;
  wire \bdatw[9]_INST_0_i_65_n_0 ;
  wire \bdatw[9]_INST_0_i_70_n_0 ;
  wire \bdatw[9]_INST_0_i_71_n_0 ;
  wire \bdatw[9]_INST_0_i_72_n_0 ;
  wire \bdatw[9]_INST_0_i_73_n_0 ;
  wire \bdatw[9]_INST_0_i_74_n_0 ;
  wire \bdatw[9]_INST_0_i_75_n_0 ;
  wire \bdatw[9]_INST_0_i_76_n_0 ;
  wire \bdatw[9]_INST_0_i_77_n_0 ;
  wire \bdatw[9]_INST_0_i_7_n_0 ;
  wire \bdatw[9]_INST_0_i_8_n_0 ;
  wire brdy;
  wire [15:0]c0bus;
  wire [15:0]c1bus;
  wire [15:0]cbus_i;
  wire [4:0]ccmd;
  wire \ccmd[0]_INST_0_i_10_n_0 ;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_13_n_0 ;
  wire \ccmd[0]_INST_0_i_14_n_0 ;
  wire \ccmd[0]_INST_0_i_15_n_0 ;
  wire \ccmd[0]_INST_0_i_16_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_19_n_0 ;
  wire \ccmd[0]_INST_0_i_1_n_0 ;
  wire \ccmd[0]_INST_0_i_20_n_0 ;
  wire \ccmd[0]_INST_0_i_21_n_0 ;
  wire \ccmd[0]_INST_0_i_22_n_0 ;
  wire \ccmd[0]_INST_0_i_23_n_0 ;
  wire \ccmd[0]_INST_0_i_24_n_0 ;
  wire \ccmd[0]_INST_0_i_25_n_0 ;
  wire \ccmd[0]_INST_0_i_26_n_0 ;
  wire \ccmd[0]_INST_0_i_27_n_0 ;
  wire \ccmd[0]_INST_0_i_28_n_0 ;
  wire \ccmd[0]_INST_0_i_29_n_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_30_n_0 ;
  wire \ccmd[0]_INST_0_i_31_n_0 ;
  wire \ccmd[0]_INST_0_i_32_n_0 ;
  wire \ccmd[0]_INST_0_i_33_n_0 ;
  wire \ccmd[0]_INST_0_i_34_n_0 ;
  wire \ccmd[0]_INST_0_i_35_n_0 ;
  wire \ccmd[0]_INST_0_i_36_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_6_n_0 ;
  wire \ccmd[0]_INST_0_i_7_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1]_INST_0_i_10_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_12_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_15_n_0 ;
  wire \ccmd[1]_INST_0_i_16_n_0 ;
  wire \ccmd[1]_INST_0_i_17_n_0 ;
  wire \ccmd[1]_INST_0_i_18_n_0 ;
  wire \ccmd[1]_INST_0_i_19_n_0 ;
  wire \ccmd[1]_INST_0_i_1_n_0 ;
  wire \ccmd[1]_INST_0_i_20_n_0 ;
  wire \ccmd[1]_INST_0_i_21_n_0 ;
  wire \ccmd[1]_INST_0_i_22_n_0 ;
  wire \ccmd[1]_INST_0_i_23_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_6_n_0 ;
  wire \ccmd[1]_INST_0_i_7_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_10_n_0 ;
  wire \ccmd[2]_INST_0_i_11_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_13_n_0 ;
  wire \ccmd[2]_INST_0_i_14_n_0 ;
  wire \ccmd[2]_INST_0_i_15_n_0 ;
  wire \ccmd[2]_INST_0_i_16_n_0 ;
  wire \ccmd[2]_INST_0_i_17_n_0 ;
  wire \ccmd[2]_INST_0_i_18_n_0 ;
  wire \ccmd[2]_INST_0_i_19_n_0 ;
  wire \ccmd[2]_INST_0_i_1_n_0 ;
  wire \ccmd[2]_INST_0_i_20_n_0 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_3_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[2]_INST_0_i_7_n_0 ;
  wire \ccmd[2]_INST_0_i_8_n_0 ;
  wire \ccmd[2]_INST_0_i_9_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_12_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_14_n_0 ;
  wire \ccmd[3]_INST_0_i_15_n_0 ;
  wire \ccmd[3]_INST_0_i_16_n_0 ;
  wire \ccmd[3]_INST_0_i_1_n_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_8_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire \ccmd[4]_INST_0_i_10_n_0 ;
  wire \ccmd[4]_INST_0_i_11_n_0 ;
  wire \ccmd[4]_INST_0_i_12_n_0 ;
  wire \ccmd[4]_INST_0_i_13_n_0 ;
  wire \ccmd[4]_INST_0_i_14_n_0 ;
  wire \ccmd[4]_INST_0_i_15_n_0 ;
  wire \ccmd[4]_INST_0_i_16_n_0 ;
  wire \ccmd[4]_INST_0_i_17_n_0 ;
  wire \ccmd[4]_INST_0_i_18_n_0 ;
  wire \ccmd[4]_INST_0_i_19_n_0 ;
  wire \ccmd[4]_INST_0_i_1_n_0 ;
  wire \ccmd[4]_INST_0_i_20_n_0 ;
  wire \ccmd[4]_INST_0_i_21_n_0 ;
  wire \ccmd[4]_INST_0_i_22_n_0 ;
  wire \ccmd[4]_INST_0_i_2_n_0 ;
  wire \ccmd[4]_INST_0_i_3_n_0 ;
  wire \ccmd[4]_INST_0_i_4_n_0 ;
  wire \ccmd[4]_INST_0_i_5_n_0 ;
  wire \ccmd[4]_INST_0_i_6_n_0 ;
  wire \ccmd[4]_INST_0_i_7_n_0 ;
  wire \ccmd[4]_INST_0_i_8_n_0 ;
  wire \ccmd[4]_INST_0_i_9_n_0 ;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire [2:0]\ctl0/stat ;
  wire [2:0]\ctl0/stat_nx ;
  wire [2:0]\ctl1/stat ;
  wire [2:0]\ctl1/stat_nx ;
  wire ctl_bcc_take0_fl_i_1_n_0;
  wire ctl_bcc_take1;
  wire ctl_bcc_take1_fl_i_1_n_0;
  wire ctl_fetch0;
  wire ctl_fetch0_fl_i_10_n_0;
  wire ctl_fetch0_fl_i_11_n_0;
  wire ctl_fetch0_fl_i_12_n_0;
  wire ctl_fetch0_fl_i_13_n_0;
  wire ctl_fetch0_fl_i_14_n_0;
  wire ctl_fetch0_fl_i_15_n_0;
  wire ctl_fetch0_fl_i_16_n_0;
  wire ctl_fetch0_fl_i_17_n_0;
  wire ctl_fetch0_fl_i_18_n_0;
  wire ctl_fetch0_fl_i_19_n_0;
  wire ctl_fetch0_fl_i_20_n_0;
  wire ctl_fetch0_fl_i_21_n_0;
  wire ctl_fetch0_fl_i_22_n_0;
  wire ctl_fetch0_fl_i_23_n_0;
  wire ctl_fetch0_fl_i_24_n_0;
  wire ctl_fetch0_fl_i_25_n_0;
  wire ctl_fetch0_fl_i_26_n_0;
  wire ctl_fetch0_fl_i_27_n_0;
  wire ctl_fetch0_fl_i_28_n_0;
  wire ctl_fetch0_fl_i_29_n_0;
  wire ctl_fetch0_fl_i_2_n_0;
  wire ctl_fetch0_fl_i_30_n_0;
  wire ctl_fetch0_fl_i_31_n_0;
  wire ctl_fetch0_fl_i_32_n_0;
  wire ctl_fetch0_fl_i_33_n_0;
  wire ctl_fetch0_fl_i_34_n_0;
  wire ctl_fetch0_fl_i_35_n_0;
  wire ctl_fetch0_fl_i_36_n_0;
  wire ctl_fetch0_fl_i_37_n_0;
  wire ctl_fetch0_fl_i_38_n_0;
  wire ctl_fetch0_fl_i_39_n_0;
  wire ctl_fetch0_fl_i_3_n_0;
  wire ctl_fetch0_fl_i_40_n_0;
  wire ctl_fetch0_fl_i_4_n_0;
  wire ctl_fetch0_fl_i_5_n_0;
  wire ctl_fetch0_fl_i_6_n_0;
  wire ctl_fetch0_fl_i_7_n_0;
  wire ctl_fetch0_fl_i_8_n_0;
  wire ctl_fetch0_fl_i_9_n_0;
  wire ctl_fetch1;
  wire ctl_fetch1_fl_i_10_n_0;
  wire ctl_fetch1_fl_i_11_n_0;
  wire ctl_fetch1_fl_i_12_n_0;
  wire ctl_fetch1_fl_i_13_n_0;
  wire ctl_fetch1_fl_i_14_n_0;
  wire ctl_fetch1_fl_i_15_n_0;
  wire ctl_fetch1_fl_i_16_n_0;
  wire ctl_fetch1_fl_i_17_n_0;
  wire ctl_fetch1_fl_i_18_n_0;
  wire ctl_fetch1_fl_i_19_n_0;
  wire ctl_fetch1_fl_i_20_n_0;
  wire ctl_fetch1_fl_i_21_n_0;
  wire ctl_fetch1_fl_i_22_n_0;
  wire ctl_fetch1_fl_i_23_n_0;
  wire ctl_fetch1_fl_i_24_n_0;
  wire ctl_fetch1_fl_i_25_n_0;
  wire ctl_fetch1_fl_i_26_n_0;
  wire ctl_fetch1_fl_i_27_n_0;
  wire ctl_fetch1_fl_i_28_n_0;
  wire ctl_fetch1_fl_i_29_n_0;
  wire ctl_fetch1_fl_i_2_n_0;
  wire ctl_fetch1_fl_i_30_n_0;
  wire ctl_fetch1_fl_i_31_n_0;
  wire ctl_fetch1_fl_i_32_n_0;
  wire ctl_fetch1_fl_i_33_n_0;
  wire ctl_fetch1_fl_i_34_n_0;
  wire ctl_fetch1_fl_i_35_n_0;
  wire ctl_fetch1_fl_i_36_n_0;
  wire ctl_fetch1_fl_i_37_n_0;
  wire ctl_fetch1_fl_i_38_n_0;
  wire ctl_fetch1_fl_i_39_n_0;
  wire ctl_fetch1_fl_i_3_n_0;
  wire ctl_fetch1_fl_i_40_n_0;
  wire ctl_fetch1_fl_i_41_n_0;
  wire ctl_fetch1_fl_i_42_n_0;
  wire ctl_fetch1_fl_i_43_n_0;
  wire ctl_fetch1_fl_i_4_n_0;
  wire ctl_fetch1_fl_i_5_n_0;
  wire ctl_fetch1_fl_i_6_n_0;
  wire ctl_fetch1_fl_i_7_n_0;
  wire ctl_fetch1_fl_i_8_n_0;
  wire ctl_fetch1_fl_i_9_n_0;
  wire ctl_fetch_ext1;
  wire ctl_fetch_ext_fl_i_1_n_0;
  wire [0:0]ctl_sela0;
  wire [2:0]ctl_sela0_rn;
  wire [0:0]ctl_sela1;
  wire [0:0]ctl_sela1_rn;
  wire [1:0]ctl_selb0_rn;
  wire [0:0]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [1:1]ctl_selc0;
  wire [1:1]ctl_selc0_rn;
  wire [1:1]ctl_selc1;
  wire [2:0]ctl_selc1_rn;
  wire ctl_sp_dec1;
  wire ctl_sp_inc1;
  wire ctl_sr_ldie0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  wire \eir_fl[15]_i_1_n_0 ;
  wire \eir_fl[1]_i_1_n_0 ;
  wire \eir_fl[2]_i_1_n_0 ;
  wire \eir_fl[3]_i_1_n_0 ;
  wire \eir_fl[4]_i_1_n_0 ;
  wire \eir_fl[5]_i_1_n_0 ;
  wire \eir_fl[6]_i_1_n_0 ;
  wire \eir_fl[6]_i_2_n_0 ;
  wire eir_inferred_i_17_n_0;
  wire eir_inferred_i_18_n_0;
  wire eir_inferred_i_19_n_0;
  wire eir_inferred_i_20_n_0;
  wire eir_inferred_i_21_n_0;
  wire eir_inferred_i_22_n_0;
  wire eir_inferred_i_23_n_0;
  wire eir_inferred_i_24_n_0;
  wire eir_inferred_i_25_n_0;
  wire eir_inferred_i_26_n_0;
  wire eir_inferred_i_27_n_0;
  wire eir_inferred_i_28_n_0;
  wire eir_inferred_i_29_n_0;
  wire eir_inferred_i_30_n_0;
  wire eir_inferred_i_31_n_0;
  wire eir_inferred_i_32_n_0;
  wire [15:0]fadr;
  wire \fadr[15]_INST_0_i_10_n_0 ;
  wire \fadr[15]_INST_0_i_11_n_0 ;
  wire \fadr[15]_INST_0_i_12_n_0 ;
  wire \fadr[15]_INST_0_i_14_n_0 ;
  wire \fadr[15]_INST_0_i_15_n_0 ;
  wire \fadr[15]_INST_0_i_17_n_0 ;
  wire \fadr[15]_INST_0_i_18_n_0 ;
  wire \fadr[15]_INST_0_i_19_n_0 ;
  wire \fadr[15]_INST_0_i_1_n_0 ;
  wire \fadr[15]_INST_0_i_20_n_0 ;
  wire \fadr[15]_INST_0_i_21_n_0 ;
  wire \fadr[15]_INST_0_i_2_n_0 ;
  wire \fadr[15]_INST_0_i_3_n_0 ;
  wire \fadr[15]_INST_0_i_4_n_0 ;
  wire \fadr[15]_INST_0_i_5_n_0 ;
  wire \fadr[15]_INST_0_i_6_n_0 ;
  wire \fadr[15]_INST_0_i_7_n_0 ;
  wire \fadr[15]_INST_0_i_8_n_0 ;
  wire \fadr[15]_INST_0_i_9_n_0 ;
  wire \fch/ctl_bcc_take0_fl ;
  wire \fch/ctl_bcc_take1_fl ;
  wire \fch/ctl_fetch0_fl ;
  wire \fch/ctl_fetch1_fl ;
  wire \fch/ctl_fetch_ext_fl ;
  (* DONT_TOUCH *) wire [15:0]\fch/eir ;
  wire \fch/eir_fl_reg_n_0_[0] ;
  wire \fch/eir_fl_reg_n_0_[10] ;
  wire \fch/eir_fl_reg_n_0_[11] ;
  wire \fch/eir_fl_reg_n_0_[12] ;
  wire \fch/eir_fl_reg_n_0_[13] ;
  wire \fch/eir_fl_reg_n_0_[14] ;
  wire \fch/eir_fl_reg_n_0_[15] ;
  wire \fch/eir_fl_reg_n_0_[1] ;
  wire \fch/eir_fl_reg_n_0_[2] ;
  wire \fch/eir_fl_reg_n_0_[3] ;
  wire \fch/eir_fl_reg_n_0_[4] ;
  wire \fch/eir_fl_reg_n_0_[5] ;
  wire \fch/eir_fl_reg_n_0_[6] ;
  wire \fch/eir_fl_reg_n_0_[7] ;
  wire \fch/eir_fl_reg_n_0_[8] ;
  wire \fch/eir_fl_reg_n_0_[9] ;
  wire \fch/fadr_1_fl ;
  wire \fch/fch_irq_req_fl ;
  (* DONT_TOUCH *) wire \fch/fch_issu1 ;
  wire \fch/fch_issu1_fl ;
  wire \fch/fch_issu1_ir ;
  wire \fch/fch_leir_hir ;
  wire \fch/fch_leir_lir ;
  wire \fch/fch_leir_nir ;
  wire \fch/fch_pc_nx2_carry__0_n_0 ;
  wire \fch/fch_pc_nx2_carry__0_n_1 ;
  wire \fch/fch_pc_nx2_carry__0_n_2 ;
  wire \fch/fch_pc_nx2_carry__0_n_3 ;
  wire \fch/fch_pc_nx2_carry__1_n_0 ;
  wire \fch/fch_pc_nx2_carry__1_n_1 ;
  wire \fch/fch_pc_nx2_carry__1_n_2 ;
  wire \fch/fch_pc_nx2_carry__1_n_3 ;
  wire \fch/fch_pc_nx2_carry__2_n_1 ;
  wire \fch/fch_pc_nx2_carry__2_n_2 ;
  wire \fch/fch_pc_nx2_carry__2_n_3 ;
  wire \fch/fch_pc_nx2_carry_n_0 ;
  wire \fch/fch_pc_nx2_carry_n_1 ;
  wire \fch/fch_pc_nx2_carry_n_2 ;
  wire \fch/fch_pc_nx2_carry_n_3 ;
  wire \fch/fch_pc_nx4_carry__0_n_0 ;
  wire \fch/fch_pc_nx4_carry__0_n_1 ;
  wire \fch/fch_pc_nx4_carry__0_n_2 ;
  wire \fch/fch_pc_nx4_carry__0_n_3 ;
  wire \fch/fch_pc_nx4_carry__0_n_4 ;
  wire \fch/fch_pc_nx4_carry__0_n_5 ;
  wire \fch/fch_pc_nx4_carry__0_n_6 ;
  wire \fch/fch_pc_nx4_carry__0_n_7 ;
  wire \fch/fch_pc_nx4_carry__1_n_0 ;
  wire \fch/fch_pc_nx4_carry__1_n_1 ;
  wire \fch/fch_pc_nx4_carry__1_n_2 ;
  wire \fch/fch_pc_nx4_carry__1_n_3 ;
  wire \fch/fch_pc_nx4_carry__1_n_4 ;
  wire \fch/fch_pc_nx4_carry__1_n_5 ;
  wire \fch/fch_pc_nx4_carry__1_n_6 ;
  wire \fch/fch_pc_nx4_carry__1_n_7 ;
  wire \fch/fch_pc_nx4_carry__2_n_2 ;
  wire \fch/fch_pc_nx4_carry__2_n_3 ;
  wire \fch/fch_pc_nx4_carry__2_n_5 ;
  wire \fch/fch_pc_nx4_carry__2_n_6 ;
  wire \fch/fch_pc_nx4_carry__2_n_7 ;
  wire \fch/fch_pc_nx4_carry_n_0 ;
  wire \fch/fch_pc_nx4_carry_n_1 ;
  wire \fch/fch_pc_nx4_carry_n_2 ;
  wire \fch/fch_pc_nx4_carry_n_3 ;
  wire \fch/fch_pc_nx4_carry_n_4 ;
  wire \fch/fch_pc_nx4_carry_n_5 ;
  wire \fch/fch_pc_nx4_carry_n_6 ;
  wire \fch/fch_pc_nx4_carry_n_7 ;
  wire \fch/fch_term_fl ;
  wire \fch/fctl/fch_leir_hir_t ;
  wire \fch/fctl/fch_leir_lir_t ;
  wire \fch/fctl/fch_leir_nir_t ;
  wire \fch/fctl/fch_nir_lir ;
  wire [2:0]\fch/fctl/stat_nx ;
  (* DONT_TOUCH *) wire [15:0]\fch/ir0 ;
  wire [15:0]\fch/ir0_fl ;
  wire [21:21]\fch/ir0_id ;
  wire [21:20]\fch/ir0_id_fl ;
  (* DONT_TOUCH *) wire [15:0]\fch/ir1 ;
  wire [15:0]\fch/ir1_fl ;
  wire [21:20]\fch/ir1_id_fl ;
  wire [24:12]\fch/lir_id_0 ;
  wire [15:0]\fch/nir ;
  wire [24:12]\fch/nir_id ;
  wire \fch/p_0_in ;
  wire [15:0]\fch/p_2_in ;
  wire \fch/pc10_carry__0_n_0 ;
  wire \fch/pc10_carry__0_n_1 ;
  wire \fch/pc10_carry__0_n_2 ;
  wire \fch/pc10_carry__0_n_3 ;
  wire \fch/pc10_carry__0_n_4 ;
  wire \fch/pc10_carry__0_n_5 ;
  wire \fch/pc10_carry__0_n_6 ;
  wire \fch/pc10_carry__0_n_7 ;
  wire \fch/pc10_carry__1_n_0 ;
  wire \fch/pc10_carry__1_n_1 ;
  wire \fch/pc10_carry__1_n_2 ;
  wire \fch/pc10_carry__1_n_3 ;
  wire \fch/pc10_carry__1_n_4 ;
  wire \fch/pc10_carry__1_n_5 ;
  wire \fch/pc10_carry__1_n_6 ;
  wire \fch/pc10_carry__1_n_7 ;
  wire \fch/pc10_carry__2_n_1 ;
  wire \fch/pc10_carry__2_n_2 ;
  wire \fch/pc10_carry__2_n_3 ;
  wire \fch/pc10_carry__2_n_4 ;
  wire \fch/pc10_carry__2_n_5 ;
  wire \fch/pc10_carry__2_n_6 ;
  wire \fch/pc10_carry__2_n_7 ;
  wire \fch/pc10_carry_n_0 ;
  wire \fch/pc10_carry_n_1 ;
  wire \fch/pc10_carry_n_2 ;
  wire \fch/pc10_carry_n_3 ;
  wire \fch/pc10_carry_n_4 ;
  wire \fch/pc10_carry_n_5 ;
  wire \fch/pc10_carry_n_6 ;
  wire \fch/pc10_carry_n_7 ;
  wire \fch/rst_n_fl ;
  wire [2:0]\fch/stat ;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[0]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_2_n_0 ;
  wire \fch_irq_lev[1]_i_3_n_0 ;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev[1]_i_5_n_0 ;
  wire fch_irq_req;
  wire fch_issu1_inferred_i_100_n_0;
  wire fch_issu1_inferred_i_101_n_0;
  wire fch_issu1_inferred_i_102_n_0;
  wire fch_issu1_inferred_i_103_n_0;
  wire fch_issu1_inferred_i_104_n_0;
  wire fch_issu1_inferred_i_105_n_0;
  wire fch_issu1_inferred_i_106_n_0;
  wire fch_issu1_inferred_i_107_n_0;
  wire fch_issu1_inferred_i_108_n_0;
  wire fch_issu1_inferred_i_109_n_0;
  wire fch_issu1_inferred_i_10_n_0;
  wire fch_issu1_inferred_i_110_n_0;
  wire fch_issu1_inferred_i_111_n_0;
  wire fch_issu1_inferred_i_112_n_0;
  wire fch_issu1_inferred_i_113_n_0;
  wire fch_issu1_inferred_i_114_n_0;
  wire fch_issu1_inferred_i_115_n_0;
  wire fch_issu1_inferred_i_116_n_0;
  wire fch_issu1_inferred_i_117_n_0;
  wire fch_issu1_inferred_i_118_n_0;
  wire fch_issu1_inferred_i_119_n_0;
  wire fch_issu1_inferred_i_11_n_0;
  wire fch_issu1_inferred_i_120_n_0;
  wire fch_issu1_inferred_i_121_n_0;
  wire fch_issu1_inferred_i_122_n_0;
  wire fch_issu1_inferred_i_123_n_0;
  wire fch_issu1_inferred_i_124_n_0;
  wire fch_issu1_inferred_i_125_n_0;
  wire fch_issu1_inferred_i_126_n_0;
  wire fch_issu1_inferred_i_127_n_0;
  wire fch_issu1_inferred_i_128_n_0;
  wire fch_issu1_inferred_i_129_n_0;
  wire fch_issu1_inferred_i_12_n_0;
  wire fch_issu1_inferred_i_130_n_0;
  wire fch_issu1_inferred_i_131_n_0;
  wire fch_issu1_inferred_i_132_n_0;
  wire fch_issu1_inferred_i_133_n_0;
  wire fch_issu1_inferred_i_134_n_0;
  wire fch_issu1_inferred_i_135_n_0;
  wire fch_issu1_inferred_i_136_n_0;
  wire fch_issu1_inferred_i_137_n_0;
  wire fch_issu1_inferred_i_138_n_0;
  wire fch_issu1_inferred_i_139_n_0;
  wire fch_issu1_inferred_i_13_n_0;
  wire fch_issu1_inferred_i_140_n_0;
  wire fch_issu1_inferred_i_141_n_0;
  wire fch_issu1_inferred_i_142_n_0;
  wire fch_issu1_inferred_i_143_n_0;
  wire fch_issu1_inferred_i_144_n_0;
  wire fch_issu1_inferred_i_145_n_0;
  wire fch_issu1_inferred_i_146_n_0;
  wire fch_issu1_inferred_i_147_n_0;
  wire fch_issu1_inferred_i_148_n_0;
  wire fch_issu1_inferred_i_149_n_0;
  wire fch_issu1_inferred_i_14_n_0;
  wire fch_issu1_inferred_i_150_n_0;
  wire fch_issu1_inferred_i_151_n_0;
  wire fch_issu1_inferred_i_152_n_0;
  wire fch_issu1_inferred_i_153_n_0;
  wire fch_issu1_inferred_i_154_n_0;
  wire fch_issu1_inferred_i_155_n_0;
  wire fch_issu1_inferred_i_156_n_0;
  wire fch_issu1_inferred_i_157_n_0;
  wire fch_issu1_inferred_i_158_n_0;
  wire fch_issu1_inferred_i_159_n_0;
  wire fch_issu1_inferred_i_15_n_0;
  wire fch_issu1_inferred_i_160_n_0;
  wire fch_issu1_inferred_i_161_n_0;
  wire fch_issu1_inferred_i_162_n_0;
  wire fch_issu1_inferred_i_163_n_0;
  wire fch_issu1_inferred_i_164_n_0;
  wire fch_issu1_inferred_i_165_n_0;
  wire fch_issu1_inferred_i_166_n_0;
  wire fch_issu1_inferred_i_167_n_0;
  wire fch_issu1_inferred_i_168_n_0;
  wire fch_issu1_inferred_i_169_n_0;
  wire fch_issu1_inferred_i_16_n_0;
  wire fch_issu1_inferred_i_170_n_0;
  wire fch_issu1_inferred_i_171_n_0;
  wire fch_issu1_inferred_i_172_n_0;
  wire fch_issu1_inferred_i_173_n_0;
  wire fch_issu1_inferred_i_174_n_0;
  wire fch_issu1_inferred_i_175_n_0;
  wire fch_issu1_inferred_i_176_n_0;
  wire fch_issu1_inferred_i_177_n_0;
  wire fch_issu1_inferred_i_178_n_0;
  wire fch_issu1_inferred_i_179_n_0;
  wire fch_issu1_inferred_i_17_n_0;
  wire fch_issu1_inferred_i_180_n_0;
  wire fch_issu1_inferred_i_181_n_0;
  wire fch_issu1_inferred_i_182_n_0;
  wire fch_issu1_inferred_i_183_n_0;
  wire fch_issu1_inferred_i_184_n_0;
  wire fch_issu1_inferred_i_185_n_0;
  wire fch_issu1_inferred_i_186_n_0;
  wire fch_issu1_inferred_i_187_n_0;
  wire fch_issu1_inferred_i_188_n_0;
  wire fch_issu1_inferred_i_189_n_0;
  wire fch_issu1_inferred_i_18_n_0;
  wire fch_issu1_inferred_i_190_n_0;
  wire fch_issu1_inferred_i_191_n_0;
  wire fch_issu1_inferred_i_192_n_0;
  wire fch_issu1_inferred_i_193_n_0;
  wire fch_issu1_inferred_i_194_n_0;
  wire fch_issu1_inferred_i_195_n_0;
  wire fch_issu1_inferred_i_196_n_0;
  wire fch_issu1_inferred_i_197_n_0;
  wire fch_issu1_inferred_i_198_n_0;
  wire fch_issu1_inferred_i_199_n_0;
  wire fch_issu1_inferred_i_19_n_0;
  wire fch_issu1_inferred_i_200_n_0;
  wire fch_issu1_inferred_i_201_n_0;
  wire fch_issu1_inferred_i_20_n_0;
  wire fch_issu1_inferred_i_21_n_0;
  wire fch_issu1_inferred_i_22_n_0;
  wire fch_issu1_inferred_i_23_n_0;
  wire fch_issu1_inferred_i_24_n_0;
  wire fch_issu1_inferred_i_25_n_0;
  wire fch_issu1_inferred_i_26_n_0;
  wire fch_issu1_inferred_i_27_n_0;
  wire fch_issu1_inferred_i_28_n_0;
  wire fch_issu1_inferred_i_29_n_0;
  wire fch_issu1_inferred_i_2_n_0;
  wire fch_issu1_inferred_i_30_n_0;
  wire fch_issu1_inferred_i_31_n_0;
  wire fch_issu1_inferred_i_32_n_0;
  wire fch_issu1_inferred_i_33_n_0;
  wire fch_issu1_inferred_i_34_n_0;
  wire fch_issu1_inferred_i_35_n_0;
  wire fch_issu1_inferred_i_36_n_0;
  wire fch_issu1_inferred_i_37_n_0;
  wire fch_issu1_inferred_i_38_n_0;
  wire fch_issu1_inferred_i_39_n_0;
  wire fch_issu1_inferred_i_3_n_0;
  wire fch_issu1_inferred_i_40_n_0;
  wire fch_issu1_inferred_i_41_n_0;
  wire fch_issu1_inferred_i_42_n_0;
  wire fch_issu1_inferred_i_43_n_0;
  wire fch_issu1_inferred_i_44_n_0;
  wire fch_issu1_inferred_i_45_n_0;
  wire fch_issu1_inferred_i_46_n_0;
  wire fch_issu1_inferred_i_47_n_0;
  wire fch_issu1_inferred_i_48_n_0;
  wire fch_issu1_inferred_i_49_n_0;
  wire fch_issu1_inferred_i_4_n_0;
  wire fch_issu1_inferred_i_50_n_0;
  wire fch_issu1_inferred_i_51_n_0;
  wire fch_issu1_inferred_i_52_n_0;
  wire fch_issu1_inferred_i_53_n_0;
  wire fch_issu1_inferred_i_54_n_0;
  wire fch_issu1_inferred_i_55_n_0;
  wire fch_issu1_inferred_i_56_n_0;
  wire fch_issu1_inferred_i_57_n_0;
  wire fch_issu1_inferred_i_58_n_0;
  wire fch_issu1_inferred_i_59_n_0;
  wire fch_issu1_inferred_i_5_n_0;
  wire fch_issu1_inferred_i_60_n_0;
  wire fch_issu1_inferred_i_61_n_0;
  wire fch_issu1_inferred_i_62_n_0;
  wire fch_issu1_inferred_i_63_n_0;
  wire fch_issu1_inferred_i_64_n_0;
  wire fch_issu1_inferred_i_65_n_0;
  wire fch_issu1_inferred_i_66_n_0;
  wire fch_issu1_inferred_i_67_n_0;
  wire fch_issu1_inferred_i_68_n_0;
  wire fch_issu1_inferred_i_69_n_0;
  wire fch_issu1_inferred_i_6_n_0;
  wire fch_issu1_inferred_i_70_n_0;
  wire fch_issu1_inferred_i_71_n_0;
  wire fch_issu1_inferred_i_72_n_0;
  wire fch_issu1_inferred_i_73_n_0;
  wire fch_issu1_inferred_i_74_n_0;
  wire fch_issu1_inferred_i_75_n_0;
  wire fch_issu1_inferred_i_76_n_0;
  wire fch_issu1_inferred_i_77_n_0;
  wire fch_issu1_inferred_i_78_n_0;
  wire fch_issu1_inferred_i_79_n_0;
  wire fch_issu1_inferred_i_7_n_0;
  wire fch_issu1_inferred_i_80_n_0;
  wire fch_issu1_inferred_i_81_n_0;
  wire fch_issu1_inferred_i_82_n_0;
  wire fch_issu1_inferred_i_83_n_0;
  wire fch_issu1_inferred_i_84_n_0;
  wire fch_issu1_inferred_i_85_n_0;
  wire fch_issu1_inferred_i_86_n_0;
  wire fch_issu1_inferred_i_87_n_0;
  wire fch_issu1_inferred_i_88_n_0;
  wire fch_issu1_inferred_i_89_n_0;
  wire fch_issu1_inferred_i_8_n_0;
  wire fch_issu1_inferred_i_90_n_0;
  wire fch_issu1_inferred_i_91_n_0;
  wire fch_issu1_inferred_i_92_n_0;
  wire fch_issu1_inferred_i_93_n_0;
  wire fch_issu1_inferred_i_94_n_0;
  wire fch_issu1_inferred_i_95_n_0;
  wire fch_issu1_inferred_i_96_n_0;
  wire fch_issu1_inferred_i_97_n_0;
  wire fch_issu1_inferred_i_98_n_0;
  wire fch_issu1_inferred_i_99_n_0;
  wire fch_issu1_inferred_i_9_n_0;
  wire fch_leir_hir_i_2_n_0;
  wire fch_leir_nir_i_2_n_0;
  wire fch_memacc1;
  wire [15:0]fch_pc;
  wire [15:0]fch_pc0;
  wire [15:0]fch_pc1;
  wire fch_pc_nx2_carry_i_1_n_0;
  wire fch_pc_nx4_carry_i_1_n_0;
  (* DONT_TOUCH *) wire fch_term;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire [15:0]fdat;
  wire [15:0]fdatx;
  wire \grn[15]_i_1__0_n_0 ;
  wire \grn[15]_i_1__10_n_0 ;
  wire \grn[15]_i_1__11_n_0 ;
  wire \grn[15]_i_1__12_n_0 ;
  wire \grn[15]_i_1__13_n_0 ;
  wire \grn[15]_i_1__14_n_0 ;
  wire \grn[15]_i_1__15_n_0 ;
  wire \grn[15]_i_1__16_n_0 ;
  wire \grn[15]_i_1__17_n_0 ;
  wire \grn[15]_i_1__18_n_0 ;
  wire \grn[15]_i_1__19_n_0 ;
  wire \grn[15]_i_1__1_n_0 ;
  wire \grn[15]_i_1__20_n_0 ;
  wire \grn[15]_i_1__21_n_0 ;
  wire \grn[15]_i_1__22_n_0 ;
  wire \grn[15]_i_1__23_n_0 ;
  wire \grn[15]_i_1__24_n_0 ;
  wire \grn[15]_i_1__25_n_0 ;
  wire \grn[15]_i_1__26_n_0 ;
  wire \grn[15]_i_1__27_n_0 ;
  wire \grn[15]_i_1__28_n_0 ;
  wire \grn[15]_i_1__29_n_0 ;
  wire \grn[15]_i_1__2_n_0 ;
  wire \grn[15]_i_1__30_n_0 ;
  wire \grn[15]_i_1__3_n_0 ;
  wire \grn[15]_i_1__4_n_0 ;
  wire \grn[15]_i_1__5_n_0 ;
  wire \grn[15]_i_1__6_n_0 ;
  wire \grn[15]_i_1__7_n_0 ;
  wire \grn[15]_i_1__8_n_0 ;
  wire \grn[15]_i_1__9_n_0 ;
  wire \grn[15]_i_1_n_0 ;
  wire \grn[15]_i_3__1_n_0 ;
  wire \grn[15]_i_3__5_n_0 ;
  wire \grn[15]_i_3_n_0 ;
  wire \grn[15]_i_5__0_n_0 ;
  wire \grn[15]_i_7_n_0 ;
  wire \ir0_id_fl[20]_i_2_n_0 ;
  wire \ir0_id_fl[20]_i_3_n_0 ;
  wire \ir0_id_fl[20]_i_4_n_0 ;
  wire \ir0_id_fl[20]_i_5_n_0 ;
  wire \ir0_id_fl[20]_i_6_n_0 ;
  wire \ir0_id_fl[20]_i_7_n_0 ;
  wire \ir0_id_fl[20]_i_8_n_0 ;
  wire \ir0_id_fl[21]_i_10_n_0 ;
  wire \ir0_id_fl[21]_i_2_n_0 ;
  wire \ir0_id_fl[21]_i_3_n_0 ;
  wire \ir0_id_fl[21]_i_4_n_0 ;
  wire \ir0_id_fl[21]_i_5_n_0 ;
  wire \ir0_id_fl[21]_i_6_n_0 ;
  wire \ir0_id_fl[21]_i_7_n_0 ;
  wire \ir0_id_fl[21]_i_8_n_0 ;
  wire \ir0_id_fl[21]_i_9_n_0 ;
  wire ir0_inferred_i_17_n_0;
  wire ir0_inferred_i_18_n_0;
  wire ir0_inferred_i_19_n_0;
  wire ir0_inferred_i_20_n_0;
  wire ir0_inferred_i_21_n_0;
  wire ir0_inferred_i_22_n_0;
  wire ir0_inferred_i_23_n_0;
  wire ir0_inferred_i_24_n_0;
  wire ir0_inferred_i_25_n_0;
  wire ir0_inferred_i_26_n_0;
  wire ir0_inferred_i_27_n_0;
  wire ir0_inferred_i_28_n_0;
  wire ir0_inferred_i_29_n_0;
  wire ir0_inferred_i_30_n_0;
  wire ir0_inferred_i_31_n_0;
  wire ir0_inferred_i_32_n_0;
  wire ir0_inferred_i_33_n_0;
  wire \ir1_id_fl[20]_i_2_n_0 ;
  wire \ir1_id_fl[21]_i_2_n_0 ;
  wire ir1_inferred_i_17_n_0;
  wire ir1_inferred_i_18_n_0;
  wire ir1_inferred_i_19_n_0;
  wire ir1_inferred_i_20_n_0;
  wire ir1_inferred_i_21_n_0;
  wire ir1_inferred_i_22_n_0;
  wire ir1_inferred_i_23_n_0;
  wire ir1_inferred_i_24_n_0;
  wire ir1_inferred_i_25_n_0;
  wire ir1_inferred_i_26_n_0;
  wire ir1_inferred_i_27_n_0;
  wire ir1_inferred_i_28_n_0;
  wire ir1_inferred_i_29_n_0;
  wire ir1_inferred_i_30_n_0;
  wire ir1_inferred_i_31_n_0;
  wire ir1_inferred_i_32_n_0;
  wire ir1_inferred_i_33_n_0;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [5:4]\mem/bctl/ctl/p_0_in ;
  wire [1:0]\mem/bctl/ctl/stat_nx ;
  wire \mem/bctl/fch_term_fl ;
  wire \mem/mem_accslot ;
  wire [3:0]\mem/read_cyc ;
  wire \nir_id[12]_i_2_n_0 ;
  wire \nir_id[12]_i_3_n_0 ;
  wire \nir_id[12]_i_4_n_0 ;
  wire \nir_id[13]_i_2_n_0 ;
  wire \nir_id[13]_i_3_n_0 ;
  wire \nir_id[13]_i_4_n_0 ;
  wire \nir_id[13]_i_5_n_0 ;
  wire \nir_id[13]_i_6_n_0 ;
  wire \nir_id[13]_i_7_n_0 ;
  wire \nir_id[14]_i_10_n_0 ;
  wire \nir_id[14]_i_11_n_0 ;
  wire \nir_id[14]_i_12_n_0 ;
  wire \nir_id[14]_i_13_n_0 ;
  wire \nir_id[14]_i_2_n_0 ;
  wire \nir_id[14]_i_3_n_0 ;
  wire \nir_id[14]_i_4_n_0 ;
  wire \nir_id[14]_i_5_n_0 ;
  wire \nir_id[14]_i_6_n_0 ;
  wire \nir_id[14]_i_7_n_0 ;
  wire \nir_id[14]_i_8_n_0 ;
  wire \nir_id[14]_i_9_n_0 ;
  wire \nir_id[15]_i_2_n_0 ;
  wire \nir_id[16]_i_2_n_0 ;
  wire \nir_id[16]_i_3_n_0 ;
  wire \nir_id[17]_i_2_n_0 ;
  wire \nir_id[17]_i_3_n_0 ;
  wire \nir_id[17]_i_4_n_0 ;
  wire \nir_id[17]_i_5_n_0 ;
  wire \nir_id[18]_i_2_n_0 ;
  wire \nir_id[18]_i_3_n_0 ;
  wire \nir_id[18]_i_4_n_0 ;
  wire \nir_id[19]_i_10_n_0 ;
  wire \nir_id[19]_i_11_n_0 ;
  wire \nir_id[19]_i_12_n_0 ;
  wire \nir_id[19]_i_2_n_0 ;
  wire \nir_id[19]_i_3_n_0 ;
  wire \nir_id[19]_i_4_n_0 ;
  wire \nir_id[19]_i_5_n_0 ;
  wire \nir_id[19]_i_6_n_0 ;
  wire \nir_id[19]_i_7_n_0 ;
  wire \nir_id[19]_i_8_n_0 ;
  wire \nir_id[19]_i_9_n_0 ;
  wire \nir_id[20]_i_1_n_0 ;
  wire \nir_id[20]_i_2_n_0 ;
  wire \nir_id[20]_i_3_n_0 ;
  wire \nir_id[20]_i_4_n_0 ;
  wire \nir_id[20]_i_5_n_0 ;
  wire \nir_id[21]_i_2_n_0 ;
  wire \nir_id[21]_i_3_n_0 ;
  wire \nir_id[21]_i_4_n_0 ;
  wire \nir_id[21]_i_5_n_0 ;
  wire \nir_id[21]_i_6_n_0 ;
  wire \nir_id[21]_i_7_n_0 ;
  wire \nir_id[21]_i_8_n_0 ;
  wire \nir_id[24]_i_10_n_0 ;
  wire \nir_id[24]_i_11_n_0 ;
  wire \nir_id[24]_i_12_n_0 ;
  wire \nir_id[24]_i_13_n_0 ;
  wire \nir_id[24]_i_14_n_0 ;
  wire \nir_id[24]_i_3_n_0 ;
  wire \nir_id[24]_i_4_n_0 ;
  wire \nir_id[24]_i_5_n_0 ;
  wire \nir_id[24]_i_6_n_0 ;
  wire \nir_id[24]_i_7_n_0 ;
  wire \nir_id[24]_i_8_n_0 ;
  wire \nir_id[24]_i_9_n_0 ;
  wire \pc0[15]_i_2_n_0 ;
  wire \pc0[15]_i_3_n_0 ;
  wire \pc0[15]_i_4_n_0 ;
  wire pc10_carry__0_i_1_n_0;
  wire pc10_carry__0_i_2_n_0;
  wire pc10_carry__0_i_3_n_0;
  wire pc10_carry__0_i_4_n_0;
  wire pc10_carry__1_i_1_n_0;
  wire pc10_carry__1_i_2_n_0;
  wire pc10_carry__1_i_3_n_0;
  wire pc10_carry__1_i_4_n_0;
  wire pc10_carry__2_i_1_n_0;
  wire pc10_carry__2_i_2_n_0;
  wire pc10_carry__2_i_3_n_0;
  wire pc10_carry__2_i_4_n_0;
  wire pc10_carry_i_1_n_0;
  wire pc10_carry_i_2_n_0;
  wire pc10_carry_i_3_n_0;
  wire pc10_carry_i_4_n_0;
  wire \pc[0]_i_2_n_0 ;
  wire \pc[10]_i_2_n_0 ;
  wire \pc[11]_i_2_n_0 ;
  wire \pc[12]_i_4_n_0 ;
  wire \pc[13]_i_4_n_0 ;
  wire \pc[14]_i_4_n_0 ;
  wire \pc[15]_i_6_n_0 ;
  wire \pc[15]_i_7_n_0 ;
  wire \pc[15]_i_8_n_0 ;
  wire \pc[1]_i_2_n_0 ;
  wire \pc[2]_i_2_n_0 ;
  wire \pc[3]_i_2_n_0 ;
  wire \pc[4]_i_4_n_0 ;
  wire \pc[5]_i_3_n_0 ;
  wire \pc[6]_i_3_n_0 ;
  wire \pc[7]_i_3_n_0 ;
  wire \pc[8]_i_4_n_0 ;
  wire \pc[8]_i_5_n_0 ;
  wire \pc[8]_i_6_n_0 ;
  wire \pc[9]_i_2_n_0 ;
  wire [15:0]\rgf/a0bus_b13 ;
  wire \rgf/a0bus_out/badr[0]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[10]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[11]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[12]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[13]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[14]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[15]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[1]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[2]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[3]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[4]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[5]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[6]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[7]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[8]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/badr[9]_INST_0_i_8_n_0 ;
  wire \rgf/a0bus_out/rgf_c0bus_wb[12]_i_35_n_0 ;
  wire [5:1]\rgf/a0bus_sel_cr ;
  wire [15:0]\rgf/a1bus_b13 ;
  wire \rgf/a1bus_out/badr[0]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[10]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[11]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[12]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[13]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[14]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[15]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[1]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[2]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[3]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[4]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[5]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[6]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[7]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[8]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/badr[9]_INST_0_i_14_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[10]_i_25_n_0 ;
  wire [5:1]\rgf/a1bus_sel_cr ;
  wire [4:0]\rgf/b0bus_b02 ;
  wire \rgf/b0bus_out/bbus_o[0]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bbus_o[0]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bbus_o[1]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[1]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bbus_o[1]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bbus_o[2]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[2]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bbus_o[2]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bbus_o[3]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[3]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bbus_o[3]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bbus_o[4]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[4]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bbus_o[4]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bbus_o[5]_INST_0_i_13_n_0 ;
  wire \rgf/b0bus_out/bbus_o[5]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[5]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bbus_o[6]_INST_0_i_13_n_0 ;
  wire \rgf/b0bus_out/bbus_o[6]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[6]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bbus_o[7]_INST_0_i_13_n_0 ;
  wire \rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[7]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bdatw[10]_INST_0_i_18_n_0 ;
  wire \rgf/b0bus_out/bdatw[10]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bdatw[10]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bdatw[11]_INST_0_i_21_n_0 ;
  wire \rgf/b0bus_out/bdatw[11]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bdatw[11]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/bdatw[12]_INST_0_i_22_n_0 ;
  wire \rgf/b0bus_out/bdatw[12]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bdatw[12]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/bdatw[13]_INST_0_i_22_n_0 ;
  wire \rgf/b0bus_out/bdatw[13]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bdatw[13]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/bdatw[14]_INST_0_i_23_n_0 ;
  wire \rgf/b0bus_out/bdatw[14]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bdatw[14]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/bdatw[15]_INST_0_i_11_n_0 ;
  wire \rgf/b0bus_out/bdatw[15]_INST_0_i_33_n_0 ;
  wire \rgf/b0bus_out/bdatw[15]_INST_0_i_8_n_0 ;
  wire \rgf/b0bus_out/bdatw[8]_INST_0_i_22_n_0 ;
  wire \rgf/b0bus_out/bdatw[8]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bdatw[8]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bdatw[9]_INST_0_i_17_n_0 ;
  wire \rgf/b0bus_out/bdatw[9]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bdatw[9]_INST_0_i_6_n_0 ;
  wire [5:0]\rgf/b0bus_sel_cr ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_10_n_0 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_13_n_0 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_27_n_0 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_35_n_0 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_38_n_0 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_62_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_12_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_15_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_33_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_41_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_44_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_66_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_12_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_15_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_32_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_40_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_43_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_65_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_12_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_15_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_33_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_41_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_44_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_62_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_12_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_15_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_35_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_43_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_46_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_64_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_147_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_14_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_17_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_54_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_62_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_65_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_10_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_13_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_29_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_37_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_40_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_68_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_12_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_25_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_32_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_35_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_59_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_9_n_0 ;
  wire [5:1]\rgf/b1bus_sel_cr ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_47_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_48_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_49_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_50_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_69_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_47_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_84_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_47_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_48_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_75_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_67_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_68_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_48_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_89_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_74_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_38_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_66_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_47_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_54_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_55_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_56_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_57_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_51_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_58_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_59_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_60_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_61_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_50_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_57_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_58_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_59_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_60_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_51_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_58_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_59_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_68_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_53_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_60_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_61_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_70_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_120_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_143_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_144_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_247_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_49_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_63_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_38_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_53_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_60_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_61_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_62_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_63_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_51_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_52_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_53_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_54_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_48_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_58_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_59_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_60_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_61_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_52_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_62_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_63_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_64_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_65_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_51_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_61_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_62_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_63_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_64_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_52_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_60_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_61_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_69_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_54_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_62_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_63_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_71_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_126_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_145_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_146_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_248_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_50_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_53_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_64_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_54_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_64_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_65_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_66_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_67_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_55_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_56_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_57_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_58_n_0 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr00 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr01 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr02 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr03 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr04 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr05 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr06 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr07 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr20 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr21 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr22 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr23 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr24 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr25 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr26 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr27 ;
  wire \rgf/bank02/grn00/grn1 ;
  wire \rgf/bank02/grn01/grn1 ;
  wire \rgf/bank02/grn02/grn1 ;
  wire \rgf/bank02/grn03/grn1 ;
  wire \rgf/bank02/grn04/grn1 ;
  wire \rgf/bank02/grn05/grn1 ;
  wire \rgf/bank02/grn06/grn1 ;
  wire \rgf/bank02/grn07/grn1 ;
  wire \rgf/bank02/grn20/grn1 ;
  wire \rgf/bank02/grn21/grn1 ;
  wire \rgf/bank02/grn22/grn1 ;
  wire \rgf/bank02/grn23/grn1 ;
  wire \rgf/bank02/grn24/grn1 ;
  wire \rgf/bank02/grn25/grn1 ;
  wire \rgf/bank02/grn26/grn1 ;
  wire \rgf/bank02/grn27/grn1 ;
  wire [15:0]\rgf/bank02/p_0_in ;
  wire [15:0]\rgf/bank02/p_0_in0_in ;
  wire [15:5]\rgf/bank02/p_0_in2_in ;
  wire [15:0]\rgf/bank02/p_1_in ;
  wire [15:0]\rgf/bank02/p_1_in1_in ;
  wire [15:5]\rgf/bank02/p_1_in3_in ;
  wire \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_37_n_0 ;
  wire \rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_38_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_53_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_54_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_55_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_26_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_57_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_58_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_70_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_46_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_92_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_95_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_76_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_68_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_45_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_46_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_71_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_51_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_52_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_101_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_98_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_51_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_52_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_77_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_69_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_63_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_64_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_53_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_54_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_67_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_68_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_52_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_53_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_66_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_67_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_53_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_54_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_63_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_64_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_70_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_71_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_55_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_65_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_66_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_72_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_73_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_132_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_135_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_148_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_149_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_249_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_250_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_55_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_55_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_69_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_70_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_60_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_61_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_51_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_52_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_65_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_66_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_55_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_69_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_70_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_54_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_55_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_68_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_69_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_55_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_65_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_66_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_72_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_73_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_57_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_58_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_67_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_68_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_74_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_75_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_138_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_141_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_150_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_151_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_251_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_252_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_57_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_58_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_57_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_58_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_71_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_72_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_62_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_63_n_0 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr00 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr01 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr02 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr03 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr04 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr05 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr06 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr07 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr20 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr21 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr22 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr23 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr24 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr25 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr26 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr27 ;
  wire \rgf/bank13/grn00/grn1 ;
  wire \rgf/bank13/grn01/grn1 ;
  wire \rgf/bank13/grn02/grn1 ;
  wire \rgf/bank13/grn03/grn1 ;
  wire \rgf/bank13/grn04/grn1 ;
  wire \rgf/bank13/grn05/grn1 ;
  wire \rgf/bank13/grn06/grn1 ;
  wire \rgf/bank13/grn07/grn1 ;
  wire \rgf/bank13/grn20/grn1 ;
  wire \rgf/bank13/grn21/grn1 ;
  wire \rgf/bank13/grn22/grn1 ;
  wire \rgf/bank13/grn23/grn1 ;
  wire \rgf/bank13/grn24/grn1 ;
  wire \rgf/bank13/grn25/grn1 ;
  wire \rgf/bank13/grn26/grn1 ;
  wire \rgf/bank13/grn27/grn1 ;
  wire [10:8]\rgf/bank13/p_0_in2_in ;
  wire [10:8]\rgf/bank13/p_1_in3_in ;
  wire [3:0]\rgf/bank_sel ;
  wire [5:5]\rgf/c0bus_sel_0 ;
  wire [5:0]\rgf/c0bus_sel_cr ;
  wire [4:1]\rgf/c1bus_sel_cr ;
  (* DONT_TOUCH *) wire [15:0]\rgf/ivec/iv ;
  wire [15:0]\rgf/ivec/p_1_in ;
  wire [15:0]\rgf/p_2_in ;
  wire [15:0]\rgf/pcnt/p_1_in ;
  (* DONT_TOUCH *) wire [15:0]\rgf/pcnt/pc ;
  wire [4:0]\rgf/rctl/p_0_in ;
  wire \rgf/rctl/p_2_in ;
  wire [15:0]\rgf/rctl/rgf_c0bus_wb ;
  wire [15:0]\rgf/rctl/rgf_c1bus_wb ;
  wire [2:0]\rgf/rctl/rgf_selc0_rn_wb ;
  wire \rgf/rctl/rgf_selc0_stat ;
  wire [1:0]\rgf/rctl/rgf_selc0_wb ;
  wire [1:0]\rgf/rctl/rgf_selc1 ;
  wire [2:0]\rgf/rctl/rgf_selc1_rn ;
  wire [2:0]\rgf/rctl/rgf_selc1_rn_wb ;
  wire \rgf/rctl/rgf_selc1_stat ;
  wire [1:0]\rgf/rctl/rgf_selc1_wb ;
  wire [15:0]\rgf/rgf_c0bus_0 ;
  wire [15:0]\rgf/rgf_c1bus_0 ;
  wire [15:1]\rgf/sptr/data2 ;
  wire [15:0]\rgf/sptr/data3 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/sptr/sp ;
  wire [15:0]\rgf/sreg/p_0_in ;
  (* DONT_TOUCH *) wire [15:0]\rgf/sreg/sr ;
  wire \rgf/treg/p_0_in ;
  wire [15:0]\rgf/treg/p_1_in ;
  (* DONT_TOUCH *) wire [15:0]\rgf/treg/tr ;
  wire \rgf_c0bus_wb[0]_i_10_n_0 ;
  wire \rgf_c0bus_wb[0]_i_11_n_0 ;
  wire \rgf_c0bus_wb[0]_i_12_n_0 ;
  wire \rgf_c0bus_wb[0]_i_13_n_0 ;
  wire \rgf_c0bus_wb[0]_i_14_n_0 ;
  wire \rgf_c0bus_wb[0]_i_15_n_0 ;
  wire \rgf_c0bus_wb[0]_i_16_n_0 ;
  wire \rgf_c0bus_wb[0]_i_17_n_0 ;
  wire \rgf_c0bus_wb[0]_i_2_n_0 ;
  wire \rgf_c0bus_wb[0]_i_4_n_0 ;
  wire \rgf_c0bus_wb[0]_i_5_n_0 ;
  wire \rgf_c0bus_wb[0]_i_6_n_0 ;
  wire \rgf_c0bus_wb[0]_i_7_n_0 ;
  wire \rgf_c0bus_wb[0]_i_8_n_0 ;
  wire \rgf_c0bus_wb[0]_i_9_n_0 ;
  wire \rgf_c0bus_wb[10]_i_10_n_0 ;
  wire \rgf_c0bus_wb[10]_i_11_n_0 ;
  wire \rgf_c0bus_wb[10]_i_12_n_0 ;
  wire \rgf_c0bus_wb[10]_i_13_n_0 ;
  wire \rgf_c0bus_wb[10]_i_14_n_0 ;
  wire \rgf_c0bus_wb[10]_i_15_n_0 ;
  wire \rgf_c0bus_wb[10]_i_16_n_0 ;
  wire \rgf_c0bus_wb[10]_i_17_n_0 ;
  wire \rgf_c0bus_wb[10]_i_18_n_0 ;
  wire \rgf_c0bus_wb[10]_i_19_n_0 ;
  wire \rgf_c0bus_wb[10]_i_20_n_0 ;
  wire \rgf_c0bus_wb[10]_i_21_n_0 ;
  wire \rgf_c0bus_wb[10]_i_22_n_0 ;
  wire \rgf_c0bus_wb[10]_i_23_n_0 ;
  wire \rgf_c0bus_wb[10]_i_2_n_0 ;
  wire \rgf_c0bus_wb[10]_i_4_n_0 ;
  wire \rgf_c0bus_wb[10]_i_5_n_0 ;
  wire \rgf_c0bus_wb[10]_i_6_n_0 ;
  wire \rgf_c0bus_wb[10]_i_7_n_0 ;
  wire \rgf_c0bus_wb[10]_i_8_n_0 ;
  wire \rgf_c0bus_wb[10]_i_9_n_0 ;
  wire \rgf_c0bus_wb[11]_i_10_n_0 ;
  wire \rgf_c0bus_wb[11]_i_11_n_0 ;
  wire \rgf_c0bus_wb[11]_i_12_n_0 ;
  wire \rgf_c0bus_wb[11]_i_13_n_0 ;
  wire \rgf_c0bus_wb[11]_i_14_n_0 ;
  wire \rgf_c0bus_wb[11]_i_15_n_0 ;
  wire \rgf_c0bus_wb[11]_i_16_n_0 ;
  wire \rgf_c0bus_wb[11]_i_17_n_0 ;
  wire \rgf_c0bus_wb[11]_i_18_n_0 ;
  wire \rgf_c0bus_wb[11]_i_2_n_0 ;
  wire \rgf_c0bus_wb[11]_i_3_n_0 ;
  wire \rgf_c0bus_wb[11]_i_4_n_0 ;
  wire \rgf_c0bus_wb[11]_i_5_n_0 ;
  wire \rgf_c0bus_wb[11]_i_6_n_0 ;
  wire \rgf_c0bus_wb[11]_i_7_n_0 ;
  wire \rgf_c0bus_wb[11]_i_8_n_0 ;
  wire \rgf_c0bus_wb[11]_i_9_n_0 ;
  wire \rgf_c0bus_wb[12]_i_10_n_0 ;
  wire \rgf_c0bus_wb[12]_i_11_n_0 ;
  wire \rgf_c0bus_wb[12]_i_12_n_0 ;
  wire \rgf_c0bus_wb[12]_i_13_n_0 ;
  wire \rgf_c0bus_wb[12]_i_14_n_0 ;
  wire \rgf_c0bus_wb[12]_i_15_n_0 ;
  wire \rgf_c0bus_wb[12]_i_16_n_0 ;
  wire \rgf_c0bus_wb[12]_i_17_n_0 ;
  wire \rgf_c0bus_wb[12]_i_18_n_0 ;
  wire \rgf_c0bus_wb[12]_i_19_n_0 ;
  wire \rgf_c0bus_wb[12]_i_20_n_0 ;
  wire \rgf_c0bus_wb[12]_i_21_n_0 ;
  wire \rgf_c0bus_wb[12]_i_22_n_0 ;
  wire \rgf_c0bus_wb[12]_i_23_n_0 ;
  wire \rgf_c0bus_wb[12]_i_24_n_0 ;
  wire \rgf_c0bus_wb[12]_i_25_n_0 ;
  wire \rgf_c0bus_wb[12]_i_26_n_0 ;
  wire \rgf_c0bus_wb[12]_i_27_n_0 ;
  wire \rgf_c0bus_wb[12]_i_28_n_0 ;
  wire \rgf_c0bus_wb[12]_i_29_n_0 ;
  wire \rgf_c0bus_wb[12]_i_2_n_0 ;
  wire \rgf_c0bus_wb[12]_i_30_n_0 ;
  wire \rgf_c0bus_wb[12]_i_31_n_0 ;
  wire \rgf_c0bus_wb[12]_i_32_n_0 ;
  wire \rgf_c0bus_wb[12]_i_33_n_0 ;
  wire \rgf_c0bus_wb[12]_i_34_n_0 ;
  wire \rgf_c0bus_wb[12]_i_36_n_0 ;
  wire \rgf_c0bus_wb[12]_i_39_n_0 ;
  wire \rgf_c0bus_wb[12]_i_3_n_0 ;
  wire \rgf_c0bus_wb[12]_i_40_n_0 ;
  wire \rgf_c0bus_wb[12]_i_41_n_0 ;
  wire \rgf_c0bus_wb[12]_i_42_n_0 ;
  wire \rgf_c0bus_wb[12]_i_4_n_0 ;
  wire \rgf_c0bus_wb[12]_i_5_n_0 ;
  wire \rgf_c0bus_wb[12]_i_6_n_0 ;
  wire \rgf_c0bus_wb[12]_i_7_n_0 ;
  wire \rgf_c0bus_wb[12]_i_8_n_0 ;
  wire \rgf_c0bus_wb[12]_i_9_n_0 ;
  wire \rgf_c0bus_wb[13]_i_10_n_0 ;
  wire \rgf_c0bus_wb[13]_i_11_n_0 ;
  wire \rgf_c0bus_wb[13]_i_12_n_0 ;
  wire \rgf_c0bus_wb[13]_i_13_n_0 ;
  wire \rgf_c0bus_wb[13]_i_14_n_0 ;
  wire \rgf_c0bus_wb[13]_i_15_n_0 ;
  wire \rgf_c0bus_wb[13]_i_16_n_0 ;
  wire \rgf_c0bus_wb[13]_i_17_n_0 ;
  wire \rgf_c0bus_wb[13]_i_18_n_0 ;
  wire \rgf_c0bus_wb[13]_i_19_n_0 ;
  wire \rgf_c0bus_wb[13]_i_20_n_0 ;
  wire \rgf_c0bus_wb[13]_i_21_n_0 ;
  wire \rgf_c0bus_wb[13]_i_22_n_0 ;
  wire \rgf_c0bus_wb[13]_i_23_n_0 ;
  wire \rgf_c0bus_wb[13]_i_24_n_0 ;
  wire \rgf_c0bus_wb[13]_i_25_n_0 ;
  wire \rgf_c0bus_wb[13]_i_26_n_0 ;
  wire \rgf_c0bus_wb[13]_i_27_n_0 ;
  wire \rgf_c0bus_wb[13]_i_28_n_0 ;
  wire \rgf_c0bus_wb[13]_i_29_n_0 ;
  wire \rgf_c0bus_wb[13]_i_2_n_0 ;
  wire \rgf_c0bus_wb[13]_i_3_n_0 ;
  wire \rgf_c0bus_wb[13]_i_4_n_0 ;
  wire \rgf_c0bus_wb[13]_i_5_n_0 ;
  wire \rgf_c0bus_wb[13]_i_6_n_0 ;
  wire \rgf_c0bus_wb[13]_i_7_n_0 ;
  wire \rgf_c0bus_wb[13]_i_9_n_0 ;
  wire \rgf_c0bus_wb[14]_i_10_n_0 ;
  wire \rgf_c0bus_wb[14]_i_11_n_0 ;
  wire \rgf_c0bus_wb[14]_i_12_n_0 ;
  wire \rgf_c0bus_wb[14]_i_13_n_0 ;
  wire \rgf_c0bus_wb[14]_i_14_n_0 ;
  wire \rgf_c0bus_wb[14]_i_15_n_0 ;
  wire \rgf_c0bus_wb[14]_i_16_n_0 ;
  wire \rgf_c0bus_wb[14]_i_17_n_0 ;
  wire \rgf_c0bus_wb[14]_i_18_n_0 ;
  wire \rgf_c0bus_wb[14]_i_19_n_0 ;
  wire \rgf_c0bus_wb[14]_i_20_n_0 ;
  wire \rgf_c0bus_wb[14]_i_21_n_0 ;
  wire \rgf_c0bus_wb[14]_i_22_n_0 ;
  wire \rgf_c0bus_wb[14]_i_23_n_0 ;
  wire \rgf_c0bus_wb[14]_i_24_n_0 ;
  wire \rgf_c0bus_wb[14]_i_25_n_0 ;
  wire \rgf_c0bus_wb[14]_i_26_n_0 ;
  wire \rgf_c0bus_wb[14]_i_27_n_0 ;
  wire \rgf_c0bus_wb[14]_i_28_n_0 ;
  wire \rgf_c0bus_wb[14]_i_29_n_0 ;
  wire \rgf_c0bus_wb[14]_i_2_n_0 ;
  wire \rgf_c0bus_wb[14]_i_30_n_0 ;
  wire \rgf_c0bus_wb[14]_i_31_n_0 ;
  wire \rgf_c0bus_wb[14]_i_32_n_0 ;
  wire \rgf_c0bus_wb[14]_i_33_n_0 ;
  wire \rgf_c0bus_wb[14]_i_34_n_0 ;
  wire \rgf_c0bus_wb[14]_i_35_n_0 ;
  wire \rgf_c0bus_wb[14]_i_3_n_0 ;
  wire \rgf_c0bus_wb[14]_i_4_n_0 ;
  wire \rgf_c0bus_wb[14]_i_5_n_0 ;
  wire \rgf_c0bus_wb[14]_i_6_n_0 ;
  wire \rgf_c0bus_wb[14]_i_7_n_0 ;
  wire \rgf_c0bus_wb[14]_i_8_n_0 ;
  wire \rgf_c0bus_wb[14]_i_9_n_0 ;
  wire \rgf_c0bus_wb[15]_i_10_n_0 ;
  wire \rgf_c0bus_wb[15]_i_11_n_0 ;
  wire \rgf_c0bus_wb[15]_i_12_n_0 ;
  wire \rgf_c0bus_wb[15]_i_13_n_0 ;
  wire \rgf_c0bus_wb[15]_i_14_n_0 ;
  wire \rgf_c0bus_wb[15]_i_15_n_0 ;
  wire \rgf_c0bus_wb[15]_i_16_n_0 ;
  wire \rgf_c0bus_wb[15]_i_17_n_0 ;
  wire \rgf_c0bus_wb[15]_i_18_n_0 ;
  wire \rgf_c0bus_wb[15]_i_19_n_0 ;
  wire \rgf_c0bus_wb[15]_i_20_n_0 ;
  wire \rgf_c0bus_wb[15]_i_21_n_0 ;
  wire \rgf_c0bus_wb[15]_i_22_n_0 ;
  wire \rgf_c0bus_wb[15]_i_23_n_0 ;
  wire \rgf_c0bus_wb[15]_i_24_n_0 ;
  wire \rgf_c0bus_wb[15]_i_25_n_0 ;
  wire \rgf_c0bus_wb[15]_i_26_n_0 ;
  wire \rgf_c0bus_wb[15]_i_27_n_0 ;
  wire \rgf_c0bus_wb[15]_i_28_n_0 ;
  wire \rgf_c0bus_wb[15]_i_29_n_0 ;
  wire \rgf_c0bus_wb[15]_i_2_n_0 ;
  wire \rgf_c0bus_wb[15]_i_30_n_0 ;
  wire \rgf_c0bus_wb[15]_i_31_n_0 ;
  wire \rgf_c0bus_wb[15]_i_32_n_0 ;
  wire \rgf_c0bus_wb[15]_i_33_n_0 ;
  wire \rgf_c0bus_wb[15]_i_34_n_0 ;
  wire \rgf_c0bus_wb[15]_i_35_n_0 ;
  wire \rgf_c0bus_wb[15]_i_36_n_0 ;
  wire \rgf_c0bus_wb[15]_i_37_n_0 ;
  wire \rgf_c0bus_wb[15]_i_38_n_0 ;
  wire \rgf_c0bus_wb[15]_i_39_n_0 ;
  wire \rgf_c0bus_wb[15]_i_3_n_0 ;
  wire \rgf_c0bus_wb[15]_i_40_n_0 ;
  wire \rgf_c0bus_wb[15]_i_41_n_0 ;
  wire \rgf_c0bus_wb[15]_i_42_n_0 ;
  wire \rgf_c0bus_wb[15]_i_43_n_0 ;
  wire \rgf_c0bus_wb[15]_i_4_n_0 ;
  wire \rgf_c0bus_wb[15]_i_5_n_0 ;
  wire \rgf_c0bus_wb[15]_i_6_n_0 ;
  wire \rgf_c0bus_wb[15]_i_7_n_0 ;
  wire \rgf_c0bus_wb[15]_i_8_n_0 ;
  wire \rgf_c0bus_wb[15]_i_9_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10_n_0 ;
  wire \rgf_c0bus_wb[1]_i_11_n_0 ;
  wire \rgf_c0bus_wb[1]_i_12_n_0 ;
  wire \rgf_c0bus_wb[1]_i_13_n_0 ;
  wire \rgf_c0bus_wb[1]_i_14_n_0 ;
  wire \rgf_c0bus_wb[1]_i_15_n_0 ;
  wire \rgf_c0bus_wb[1]_i_16_n_0 ;
  wire \rgf_c0bus_wb[1]_i_17_n_0 ;
  wire \rgf_c0bus_wb[1]_i_18_n_0 ;
  wire \rgf_c0bus_wb[1]_i_19_n_0 ;
  wire \rgf_c0bus_wb[1]_i_20_n_0 ;
  wire \rgf_c0bus_wb[1]_i_2_n_0 ;
  wire \rgf_c0bus_wb[1]_i_3_n_0 ;
  wire \rgf_c0bus_wb[1]_i_4_n_0 ;
  wire \rgf_c0bus_wb[1]_i_5_n_0 ;
  wire \rgf_c0bus_wb[1]_i_6_n_0 ;
  wire \rgf_c0bus_wb[1]_i_7_n_0 ;
  wire \rgf_c0bus_wb[1]_i_8_n_0 ;
  wire \rgf_c0bus_wb[1]_i_9_n_0 ;
  wire \rgf_c0bus_wb[2]_i_10_n_0 ;
  wire \rgf_c0bus_wb[2]_i_11_n_0 ;
  wire \rgf_c0bus_wb[2]_i_12_n_0 ;
  wire \rgf_c0bus_wb[2]_i_2_n_0 ;
  wire \rgf_c0bus_wb[2]_i_3_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4_n_0 ;
  wire \rgf_c0bus_wb[2]_i_5_n_0 ;
  wire \rgf_c0bus_wb[2]_i_6_n_0 ;
  wire \rgf_c0bus_wb[2]_i_7_n_0 ;
  wire \rgf_c0bus_wb[2]_i_8_n_0 ;
  wire \rgf_c0bus_wb[2]_i_9_n_0 ;
  wire \rgf_c0bus_wb[3]_i_10_n_0 ;
  wire \rgf_c0bus_wb[3]_i_11_n_0 ;
  wire \rgf_c0bus_wb[3]_i_12_n_0 ;
  wire \rgf_c0bus_wb[3]_i_13_n_0 ;
  wire \rgf_c0bus_wb[3]_i_14_n_0 ;
  wire \rgf_c0bus_wb[3]_i_15_n_0 ;
  wire \rgf_c0bus_wb[3]_i_16_n_0 ;
  wire \rgf_c0bus_wb[3]_i_17_n_0 ;
  wire \rgf_c0bus_wb[3]_i_18_n_0 ;
  wire \rgf_c0bus_wb[3]_i_2_n_0 ;
  wire \rgf_c0bus_wb[3]_i_3_n_0 ;
  wire \rgf_c0bus_wb[3]_i_4_n_0 ;
  wire \rgf_c0bus_wb[3]_i_5_n_0 ;
  wire \rgf_c0bus_wb[3]_i_6_n_0 ;
  wire \rgf_c0bus_wb[3]_i_7_n_0 ;
  wire \rgf_c0bus_wb[3]_i_8_n_0 ;
  wire \rgf_c0bus_wb[3]_i_9_n_0 ;
  wire \rgf_c0bus_wb[4]_i_10_n_0 ;
  wire \rgf_c0bus_wb[4]_i_11_n_0 ;
  wire \rgf_c0bus_wb[4]_i_12_n_0 ;
  wire \rgf_c0bus_wb[4]_i_13_n_0 ;
  wire \rgf_c0bus_wb[4]_i_14_n_0 ;
  wire \rgf_c0bus_wb[4]_i_15_n_0 ;
  wire \rgf_c0bus_wb[4]_i_16_n_0 ;
  wire \rgf_c0bus_wb[4]_i_17_n_0 ;
  wire \rgf_c0bus_wb[4]_i_2_n_0 ;
  wire \rgf_c0bus_wb[4]_i_3_n_0 ;
  wire \rgf_c0bus_wb[4]_i_4_n_0 ;
  wire \rgf_c0bus_wb[4]_i_5_n_0 ;
  wire \rgf_c0bus_wb[4]_i_6_n_0 ;
  wire \rgf_c0bus_wb[4]_i_7_n_0 ;
  wire \rgf_c0bus_wb[4]_i_8_n_0 ;
  wire \rgf_c0bus_wb[4]_i_9_n_0 ;
  wire \rgf_c0bus_wb[5]_i_10_n_0 ;
  wire \rgf_c0bus_wb[5]_i_11_n_0 ;
  wire \rgf_c0bus_wb[5]_i_12_n_0 ;
  wire \rgf_c0bus_wb[5]_i_13_n_0 ;
  wire \rgf_c0bus_wb[5]_i_14_n_0 ;
  wire \rgf_c0bus_wb[5]_i_15_n_0 ;
  wire \rgf_c0bus_wb[5]_i_2_n_0 ;
  wire \rgf_c0bus_wb[5]_i_3_n_0 ;
  wire \rgf_c0bus_wb[5]_i_4_n_0 ;
  wire \rgf_c0bus_wb[5]_i_5_n_0 ;
  wire \rgf_c0bus_wb[5]_i_6_n_0 ;
  wire \rgf_c0bus_wb[5]_i_7_n_0 ;
  wire \rgf_c0bus_wb[5]_i_8_n_0 ;
  wire \rgf_c0bus_wb[5]_i_9_n_0 ;
  wire \rgf_c0bus_wb[6]_i_10_n_0 ;
  wire \rgf_c0bus_wb[6]_i_11_n_0 ;
  wire \rgf_c0bus_wb[6]_i_12_n_0 ;
  wire \rgf_c0bus_wb[6]_i_13_n_0 ;
  wire \rgf_c0bus_wb[6]_i_14_n_0 ;
  wire \rgf_c0bus_wb[6]_i_15_n_0 ;
  wire \rgf_c0bus_wb[6]_i_16_n_0 ;
  wire \rgf_c0bus_wb[6]_i_2_n_0 ;
  wire \rgf_c0bus_wb[6]_i_3_n_0 ;
  wire \rgf_c0bus_wb[6]_i_4_n_0 ;
  wire \rgf_c0bus_wb[6]_i_5_n_0 ;
  wire \rgf_c0bus_wb[6]_i_6_n_0 ;
  wire \rgf_c0bus_wb[6]_i_7_n_0 ;
  wire \rgf_c0bus_wb[6]_i_8_n_0 ;
  wire \rgf_c0bus_wb[6]_i_9_n_0 ;
  wire \rgf_c0bus_wb[7]_i_10_n_0 ;
  wire \rgf_c0bus_wb[7]_i_11_n_0 ;
  wire \rgf_c0bus_wb[7]_i_12_n_0 ;
  wire \rgf_c0bus_wb[7]_i_13_n_0 ;
  wire \rgf_c0bus_wb[7]_i_14_n_0 ;
  wire \rgf_c0bus_wb[7]_i_15_n_0 ;
  wire \rgf_c0bus_wb[7]_i_16_n_0 ;
  wire \rgf_c0bus_wb[7]_i_17_n_0 ;
  wire \rgf_c0bus_wb[7]_i_18_n_0 ;
  wire \rgf_c0bus_wb[7]_i_19_n_0 ;
  wire \rgf_c0bus_wb[7]_i_2_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3_n_0 ;
  wire \rgf_c0bus_wb[7]_i_4_n_0 ;
  wire \rgf_c0bus_wb[7]_i_5_n_0 ;
  wire \rgf_c0bus_wb[7]_i_6_n_0 ;
  wire \rgf_c0bus_wb[7]_i_7_n_0 ;
  wire \rgf_c0bus_wb[7]_i_8_n_0 ;
  wire \rgf_c0bus_wb[7]_i_9_n_0 ;
  wire \rgf_c0bus_wb[8]_i_10_n_0 ;
  wire \rgf_c0bus_wb[8]_i_11_n_0 ;
  wire \rgf_c0bus_wb[8]_i_12_n_0 ;
  wire \rgf_c0bus_wb[8]_i_13_n_0 ;
  wire \rgf_c0bus_wb[8]_i_14_n_0 ;
  wire \rgf_c0bus_wb[8]_i_15_n_0 ;
  wire \rgf_c0bus_wb[8]_i_16_n_0 ;
  wire \rgf_c0bus_wb[8]_i_2_n_0 ;
  wire \rgf_c0bus_wb[8]_i_4_n_0 ;
  wire \rgf_c0bus_wb[8]_i_5_n_0 ;
  wire \rgf_c0bus_wb[8]_i_6_n_0 ;
  wire \rgf_c0bus_wb[8]_i_7_n_0 ;
  wire \rgf_c0bus_wb[8]_i_8_n_0 ;
  wire \rgf_c0bus_wb[8]_i_9_n_0 ;
  wire \rgf_c0bus_wb[9]_i_10_n_0 ;
  wire \rgf_c0bus_wb[9]_i_11_n_0 ;
  wire \rgf_c0bus_wb[9]_i_12_n_0 ;
  wire \rgf_c0bus_wb[9]_i_13_n_0 ;
  wire \rgf_c0bus_wb[9]_i_14_n_0 ;
  wire \rgf_c0bus_wb[9]_i_15_n_0 ;
  wire \rgf_c0bus_wb[9]_i_16_n_0 ;
  wire \rgf_c0bus_wb[9]_i_17_n_0 ;
  wire \rgf_c0bus_wb[9]_i_18_n_0 ;
  wire \rgf_c0bus_wb[9]_i_19_n_0 ;
  wire \rgf_c0bus_wb[9]_i_20_n_0 ;
  wire \rgf_c0bus_wb[9]_i_21_n_0 ;
  wire \rgf_c0bus_wb[9]_i_22_n_0 ;
  wire \rgf_c0bus_wb[9]_i_2_n_0 ;
  wire \rgf_c0bus_wb[9]_i_4_n_0 ;
  wire \rgf_c0bus_wb[9]_i_5_n_0 ;
  wire \rgf_c0bus_wb[9]_i_6_n_0 ;
  wire \rgf_c0bus_wb[9]_i_7_n_0 ;
  wire \rgf_c0bus_wb[9]_i_8_n_0 ;
  wire \rgf_c0bus_wb[9]_i_9_n_0 ;
  wire \rgf_c0bus_wb_reg[0]_i_3_n_0 ;
  wire \rgf_c0bus_wb_reg[10]_i_3_n_0 ;
  wire \rgf_c0bus_wb_reg[13]_i_8_n_0 ;
  wire \rgf_c0bus_wb_reg[8]_i_3_n_0 ;
  wire \rgf_c0bus_wb_reg[9]_i_3_n_0 ;
  wire \rgf_c1bus_wb[0]_i_10_n_0 ;
  wire \rgf_c1bus_wb[0]_i_11_n_0 ;
  wire \rgf_c1bus_wb[0]_i_12_n_0 ;
  wire \rgf_c1bus_wb[0]_i_13_n_0 ;
  wire \rgf_c1bus_wb[0]_i_14_n_0 ;
  wire \rgf_c1bus_wb[0]_i_15_n_0 ;
  wire \rgf_c1bus_wb[0]_i_16_n_0 ;
  wire \rgf_c1bus_wb[0]_i_2_n_0 ;
  wire \rgf_c1bus_wb[0]_i_3_n_0 ;
  wire \rgf_c1bus_wb[0]_i_5_n_0 ;
  wire \rgf_c1bus_wb[0]_i_6_n_0 ;
  wire \rgf_c1bus_wb[0]_i_7_n_0 ;
  wire \rgf_c1bus_wb[0]_i_8_n_0 ;
  wire \rgf_c1bus_wb[0]_i_9_n_0 ;
  wire \rgf_c1bus_wb[10]_i_10_n_0 ;
  wire \rgf_c1bus_wb[10]_i_11_n_0 ;
  wire \rgf_c1bus_wb[10]_i_12_n_0 ;
  wire \rgf_c1bus_wb[10]_i_13_n_0 ;
  wire \rgf_c1bus_wb[10]_i_14_n_0 ;
  wire \rgf_c1bus_wb[10]_i_15_n_0 ;
  wire \rgf_c1bus_wb[10]_i_16_n_0 ;
  wire \rgf_c1bus_wb[10]_i_17_n_0 ;
  wire \rgf_c1bus_wb[10]_i_18_n_0 ;
  wire \rgf_c1bus_wb[10]_i_19_n_0 ;
  wire \rgf_c1bus_wb[10]_i_20_n_0 ;
  wire \rgf_c1bus_wb[10]_i_21_n_0 ;
  wire \rgf_c1bus_wb[10]_i_22_n_0 ;
  wire \rgf_c1bus_wb[10]_i_23_n_0 ;
  wire \rgf_c1bus_wb[10]_i_24_n_0 ;
  wire \rgf_c1bus_wb[10]_i_28_n_0 ;
  wire \rgf_c1bus_wb[10]_i_29_n_0 ;
  wire \rgf_c1bus_wb[10]_i_2_n_0 ;
  wire \rgf_c1bus_wb[10]_i_30_n_0 ;
  wire \rgf_c1bus_wb[10]_i_31_n_0 ;
  wire \rgf_c1bus_wb[10]_i_3_n_0 ;
  wire \rgf_c1bus_wb[10]_i_4_n_0 ;
  wire \rgf_c1bus_wb[10]_i_5_n_0 ;
  wire \rgf_c1bus_wb[10]_i_6_n_0 ;
  wire \rgf_c1bus_wb[10]_i_7_n_0 ;
  wire \rgf_c1bus_wb[10]_i_8_n_0 ;
  wire \rgf_c1bus_wb[10]_i_9_n_0 ;
  wire \rgf_c1bus_wb[11]_i_10_n_0 ;
  wire \rgf_c1bus_wb[11]_i_11_n_0 ;
  wire \rgf_c1bus_wb[11]_i_12_n_0 ;
  wire \rgf_c1bus_wb[11]_i_13_n_0 ;
  wire \rgf_c1bus_wb[11]_i_14_n_0 ;
  wire \rgf_c1bus_wb[11]_i_15_n_0 ;
  wire \rgf_c1bus_wb[11]_i_16_n_0 ;
  wire \rgf_c1bus_wb[11]_i_17_n_0 ;
  wire \rgf_c1bus_wb[11]_i_18_n_0 ;
  wire \rgf_c1bus_wb[11]_i_19_n_0 ;
  wire \rgf_c1bus_wb[11]_i_2_n_0 ;
  wire \rgf_c1bus_wb[11]_i_3_n_0 ;
  wire \rgf_c1bus_wb[11]_i_4_n_0 ;
  wire \rgf_c1bus_wb[11]_i_5_n_0 ;
  wire \rgf_c1bus_wb[11]_i_6_n_0 ;
  wire \rgf_c1bus_wb[11]_i_7_n_0 ;
  wire \rgf_c1bus_wb[11]_i_8_n_0 ;
  wire \rgf_c1bus_wb[11]_i_9_n_0 ;
  wire \rgf_c1bus_wb[12]_i_10_n_0 ;
  wire \rgf_c1bus_wb[12]_i_11_n_0 ;
  wire \rgf_c1bus_wb[12]_i_12_n_0 ;
  wire \rgf_c1bus_wb[12]_i_13_n_0 ;
  wire \rgf_c1bus_wb[12]_i_14_n_0 ;
  wire \rgf_c1bus_wb[12]_i_15_n_0 ;
  wire \rgf_c1bus_wb[12]_i_16_n_0 ;
  wire \rgf_c1bus_wb[12]_i_17_n_0 ;
  wire \rgf_c1bus_wb[12]_i_18_n_0 ;
  wire \rgf_c1bus_wb[12]_i_19_n_0 ;
  wire \rgf_c1bus_wb[12]_i_20_n_0 ;
  wire \rgf_c1bus_wb[12]_i_21_n_0 ;
  wire \rgf_c1bus_wb[12]_i_22_n_0 ;
  wire \rgf_c1bus_wb[12]_i_23_n_0 ;
  wire \rgf_c1bus_wb[12]_i_24_n_0 ;
  wire \rgf_c1bus_wb[12]_i_25_n_0 ;
  wire \rgf_c1bus_wb[12]_i_26_n_0 ;
  wire \rgf_c1bus_wb[12]_i_27_n_0 ;
  wire \rgf_c1bus_wb[12]_i_28_n_0 ;
  wire \rgf_c1bus_wb[12]_i_2_n_0 ;
  wire \rgf_c1bus_wb[12]_i_3_n_0 ;
  wire \rgf_c1bus_wb[12]_i_4_n_0 ;
  wire \rgf_c1bus_wb[12]_i_5_n_0 ;
  wire \rgf_c1bus_wb[12]_i_6_n_0 ;
  wire \rgf_c1bus_wb[12]_i_7_n_0 ;
  wire \rgf_c1bus_wb[12]_i_8_n_0 ;
  wire \rgf_c1bus_wb[12]_i_9_n_0 ;
  wire \rgf_c1bus_wb[13]_i_10_n_0 ;
  wire \rgf_c1bus_wb[13]_i_11_n_0 ;
  wire \rgf_c1bus_wb[13]_i_12_n_0 ;
  wire \rgf_c1bus_wb[13]_i_13_n_0 ;
  wire \rgf_c1bus_wb[13]_i_14_n_0 ;
  wire \rgf_c1bus_wb[13]_i_15_n_0 ;
  wire \rgf_c1bus_wb[13]_i_16_n_0 ;
  wire \rgf_c1bus_wb[13]_i_17_n_0 ;
  wire \rgf_c1bus_wb[13]_i_18_n_0 ;
  wire \rgf_c1bus_wb[13]_i_19_n_0 ;
  wire \rgf_c1bus_wb[13]_i_20_n_0 ;
  wire \rgf_c1bus_wb[13]_i_21_n_0 ;
  wire \rgf_c1bus_wb[13]_i_22_n_0 ;
  wire \rgf_c1bus_wb[13]_i_23_n_0 ;
  wire \rgf_c1bus_wb[13]_i_24_n_0 ;
  wire \rgf_c1bus_wb[13]_i_25_n_0 ;
  wire \rgf_c1bus_wb[13]_i_2_n_0 ;
  wire \rgf_c1bus_wb[13]_i_3_n_0 ;
  wire \rgf_c1bus_wb[13]_i_4_n_0 ;
  wire \rgf_c1bus_wb[13]_i_5_n_0 ;
  wire \rgf_c1bus_wb[13]_i_6_n_0 ;
  wire \rgf_c1bus_wb[13]_i_7_n_0 ;
  wire \rgf_c1bus_wb[13]_i_8_n_0 ;
  wire \rgf_c1bus_wb[13]_i_9_n_0 ;
  wire \rgf_c1bus_wb[14]_i_10_n_0 ;
  wire \rgf_c1bus_wb[14]_i_11_n_0 ;
  wire \rgf_c1bus_wb[14]_i_12_n_0 ;
  wire \rgf_c1bus_wb[14]_i_13_n_0 ;
  wire \rgf_c1bus_wb[14]_i_14_n_0 ;
  wire \rgf_c1bus_wb[14]_i_15_n_0 ;
  wire \rgf_c1bus_wb[14]_i_16_n_0 ;
  wire \rgf_c1bus_wb[14]_i_17_n_0 ;
  wire \rgf_c1bus_wb[14]_i_18_n_0 ;
  wire \rgf_c1bus_wb[14]_i_19_n_0 ;
  wire \rgf_c1bus_wb[14]_i_20_n_0 ;
  wire \rgf_c1bus_wb[14]_i_21_n_0 ;
  wire \rgf_c1bus_wb[14]_i_22_n_0 ;
  wire \rgf_c1bus_wb[14]_i_23_n_0 ;
  wire \rgf_c1bus_wb[14]_i_24_n_0 ;
  wire \rgf_c1bus_wb[14]_i_25_n_0 ;
  wire \rgf_c1bus_wb[14]_i_26_n_0 ;
  wire \rgf_c1bus_wb[14]_i_27_n_0 ;
  wire \rgf_c1bus_wb[14]_i_28_n_0 ;
  wire \rgf_c1bus_wb[14]_i_29_n_0 ;
  wire \rgf_c1bus_wb[14]_i_2_n_0 ;
  wire \rgf_c1bus_wb[14]_i_30_n_0 ;
  wire \rgf_c1bus_wb[14]_i_31_n_0 ;
  wire \rgf_c1bus_wb[14]_i_32_n_0 ;
  wire \rgf_c1bus_wb[14]_i_3_n_0 ;
  wire \rgf_c1bus_wb[14]_i_4_n_0 ;
  wire \rgf_c1bus_wb[14]_i_5_n_0 ;
  wire \rgf_c1bus_wb[14]_i_6_n_0 ;
  wire \rgf_c1bus_wb[14]_i_7_n_0 ;
  wire \rgf_c1bus_wb[14]_i_8_n_0 ;
  wire \rgf_c1bus_wb[14]_i_9_n_0 ;
  wire \rgf_c1bus_wb[15]_i_100_n_0 ;
  wire \rgf_c1bus_wb[15]_i_101_n_0 ;
  wire \rgf_c1bus_wb[15]_i_102_n_0 ;
  wire \rgf_c1bus_wb[15]_i_103_n_0 ;
  wire \rgf_c1bus_wb[15]_i_10_n_0 ;
  wire \rgf_c1bus_wb[15]_i_11_n_0 ;
  wire \rgf_c1bus_wb[15]_i_12_n_0 ;
  wire \rgf_c1bus_wb[15]_i_13_n_0 ;
  wire \rgf_c1bus_wb[15]_i_14_n_0 ;
  wire \rgf_c1bus_wb[15]_i_15_n_0 ;
  wire \rgf_c1bus_wb[15]_i_16_n_0 ;
  wire \rgf_c1bus_wb[15]_i_17_n_0 ;
  wire \rgf_c1bus_wb[15]_i_18_n_0 ;
  wire \rgf_c1bus_wb[15]_i_19_n_0 ;
  wire \rgf_c1bus_wb[15]_i_20_n_0 ;
  wire \rgf_c1bus_wb[15]_i_21_n_0 ;
  wire \rgf_c1bus_wb[15]_i_22_n_0 ;
  wire \rgf_c1bus_wb[15]_i_23_n_0 ;
  wire \rgf_c1bus_wb[15]_i_24_n_0 ;
  wire \rgf_c1bus_wb[15]_i_25_n_0 ;
  wire \rgf_c1bus_wb[15]_i_26_n_0 ;
  wire \rgf_c1bus_wb[15]_i_27_n_0 ;
  wire \rgf_c1bus_wb[15]_i_28_n_0 ;
  wire \rgf_c1bus_wb[15]_i_29_n_0 ;
  wire \rgf_c1bus_wb[15]_i_2_n_0 ;
  wire \rgf_c1bus_wb[15]_i_30_n_0 ;
  wire \rgf_c1bus_wb[15]_i_31_n_0 ;
  wire \rgf_c1bus_wb[15]_i_32_n_0 ;
  wire \rgf_c1bus_wb[15]_i_33_n_0 ;
  wire \rgf_c1bus_wb[15]_i_34_n_0 ;
  wire \rgf_c1bus_wb[15]_i_35_n_0 ;
  wire \rgf_c1bus_wb[15]_i_36_n_0 ;
  wire \rgf_c1bus_wb[15]_i_37_n_0 ;
  wire \rgf_c1bus_wb[15]_i_38_n_0 ;
  wire \rgf_c1bus_wb[15]_i_39_n_0 ;
  wire \rgf_c1bus_wb[15]_i_3_n_0 ;
  wire \rgf_c1bus_wb[15]_i_40_n_0 ;
  wire \rgf_c1bus_wb[15]_i_41_n_0 ;
  wire \rgf_c1bus_wb[15]_i_42_n_0 ;
  wire \rgf_c1bus_wb[15]_i_43_n_0 ;
  wire \rgf_c1bus_wb[15]_i_44_n_0 ;
  wire \rgf_c1bus_wb[15]_i_45_n_0 ;
  wire \rgf_c1bus_wb[15]_i_46_n_0 ;
  wire \rgf_c1bus_wb[15]_i_47_n_0 ;
  wire \rgf_c1bus_wb[15]_i_48_n_0 ;
  wire \rgf_c1bus_wb[15]_i_49_n_0 ;
  wire \rgf_c1bus_wb[15]_i_4_n_0 ;
  wire \rgf_c1bus_wb[15]_i_50_n_0 ;
  wire \rgf_c1bus_wb[15]_i_51_n_0 ;
  wire \rgf_c1bus_wb[15]_i_52_n_0 ;
  wire \rgf_c1bus_wb[15]_i_53_n_0 ;
  wire \rgf_c1bus_wb[15]_i_54_n_0 ;
  wire \rgf_c1bus_wb[15]_i_55_n_0 ;
  wire \rgf_c1bus_wb[15]_i_56_n_0 ;
  wire \rgf_c1bus_wb[15]_i_57_n_0 ;
  wire \rgf_c1bus_wb[15]_i_58_n_0 ;
  wire \rgf_c1bus_wb[15]_i_59_n_0 ;
  wire \rgf_c1bus_wb[15]_i_5_n_0 ;
  wire \rgf_c1bus_wb[15]_i_60_n_0 ;
  wire \rgf_c1bus_wb[15]_i_61_n_0 ;
  wire \rgf_c1bus_wb[15]_i_62_n_0 ;
  wire \rgf_c1bus_wb[15]_i_63_n_0 ;
  wire \rgf_c1bus_wb[15]_i_64_n_0 ;
  wire \rgf_c1bus_wb[15]_i_65_n_0 ;
  wire \rgf_c1bus_wb[15]_i_66_n_0 ;
  wire \rgf_c1bus_wb[15]_i_67_n_0 ;
  wire \rgf_c1bus_wb[15]_i_68_n_0 ;
  wire \rgf_c1bus_wb[15]_i_69_n_0 ;
  wire \rgf_c1bus_wb[15]_i_6_n_0 ;
  wire \rgf_c1bus_wb[15]_i_70_n_0 ;
  wire \rgf_c1bus_wb[15]_i_71_n_0 ;
  wire \rgf_c1bus_wb[15]_i_72_n_0 ;
  wire \rgf_c1bus_wb[15]_i_73_n_0 ;
  wire \rgf_c1bus_wb[15]_i_74_n_0 ;
  wire \rgf_c1bus_wb[15]_i_75_n_0 ;
  wire \rgf_c1bus_wb[15]_i_76_n_0 ;
  wire \rgf_c1bus_wb[15]_i_77_n_0 ;
  wire \rgf_c1bus_wb[15]_i_78_n_0 ;
  wire \rgf_c1bus_wb[15]_i_79_n_0 ;
  wire \rgf_c1bus_wb[15]_i_7_n_0 ;
  wire \rgf_c1bus_wb[15]_i_80_n_0 ;
  wire \rgf_c1bus_wb[15]_i_81_n_0 ;
  wire \rgf_c1bus_wb[15]_i_82_n_0 ;
  wire \rgf_c1bus_wb[15]_i_83_n_0 ;
  wire \rgf_c1bus_wb[15]_i_84_n_0 ;
  wire \rgf_c1bus_wb[15]_i_85_n_0 ;
  wire \rgf_c1bus_wb[15]_i_86_n_0 ;
  wire \rgf_c1bus_wb[15]_i_87_n_0 ;
  wire \rgf_c1bus_wb[15]_i_88_n_0 ;
  wire \rgf_c1bus_wb[15]_i_89_n_0 ;
  wire \rgf_c1bus_wb[15]_i_8_n_0 ;
  wire \rgf_c1bus_wb[15]_i_90_n_0 ;
  wire \rgf_c1bus_wb[15]_i_91_n_0 ;
  wire \rgf_c1bus_wb[15]_i_92_n_0 ;
  wire \rgf_c1bus_wb[15]_i_93_n_0 ;
  wire \rgf_c1bus_wb[15]_i_94_n_0 ;
  wire \rgf_c1bus_wb[15]_i_95_n_0 ;
  wire \rgf_c1bus_wb[15]_i_96_n_0 ;
  wire \rgf_c1bus_wb[15]_i_97_n_0 ;
  wire \rgf_c1bus_wb[15]_i_98_n_0 ;
  wire \rgf_c1bus_wb[15]_i_99_n_0 ;
  wire \rgf_c1bus_wb[15]_i_9_n_0 ;
  wire \rgf_c1bus_wb[1]_i_10_n_0 ;
  wire \rgf_c1bus_wb[1]_i_11_n_0 ;
  wire \rgf_c1bus_wb[1]_i_12_n_0 ;
  wire \rgf_c1bus_wb[1]_i_13_n_0 ;
  wire \rgf_c1bus_wb[1]_i_14_n_0 ;
  wire \rgf_c1bus_wb[1]_i_15_n_0 ;
  wire \rgf_c1bus_wb[1]_i_16_n_0 ;
  wire \rgf_c1bus_wb[1]_i_17_n_0 ;
  wire \rgf_c1bus_wb[1]_i_18_n_0 ;
  wire \rgf_c1bus_wb[1]_i_19_n_0 ;
  wire \rgf_c1bus_wb[1]_i_20_n_0 ;
  wire \rgf_c1bus_wb[1]_i_2_n_0 ;
  wire \rgf_c1bus_wb[1]_i_3_n_0 ;
  wire \rgf_c1bus_wb[1]_i_4_n_0 ;
  wire \rgf_c1bus_wb[1]_i_5_n_0 ;
  wire \rgf_c1bus_wb[1]_i_6_n_0 ;
  wire \rgf_c1bus_wb[1]_i_7_n_0 ;
  wire \rgf_c1bus_wb[1]_i_8_n_0 ;
  wire \rgf_c1bus_wb[1]_i_9_n_0 ;
  wire \rgf_c1bus_wb[2]_i_10_n_0 ;
  wire \rgf_c1bus_wb[2]_i_11_n_0 ;
  wire \rgf_c1bus_wb[2]_i_12_n_0 ;
  wire \rgf_c1bus_wb[2]_i_13_n_0 ;
  wire \rgf_c1bus_wb[2]_i_14_n_0 ;
  wire \rgf_c1bus_wb[2]_i_15_n_0 ;
  wire \rgf_c1bus_wb[2]_i_16_n_0 ;
  wire \rgf_c1bus_wb[2]_i_17_n_0 ;
  wire \rgf_c1bus_wb[2]_i_2_n_0 ;
  wire \rgf_c1bus_wb[2]_i_3_n_0 ;
  wire \rgf_c1bus_wb[2]_i_4_n_0 ;
  wire \rgf_c1bus_wb[2]_i_5_n_0 ;
  wire \rgf_c1bus_wb[2]_i_6_n_0 ;
  wire \rgf_c1bus_wb[2]_i_7_n_0 ;
  wire \rgf_c1bus_wb[2]_i_8_n_0 ;
  wire \rgf_c1bus_wb[2]_i_9_n_0 ;
  wire \rgf_c1bus_wb[3]_i_10_n_0 ;
  wire \rgf_c1bus_wb[3]_i_11_n_0 ;
  wire \rgf_c1bus_wb[3]_i_12_n_0 ;
  wire \rgf_c1bus_wb[3]_i_13_n_0 ;
  wire \rgf_c1bus_wb[3]_i_14_n_0 ;
  wire \rgf_c1bus_wb[3]_i_15_n_0 ;
  wire \rgf_c1bus_wb[3]_i_16_n_0 ;
  wire \rgf_c1bus_wb[3]_i_17_n_0 ;
  wire \rgf_c1bus_wb[3]_i_18_n_0 ;
  wire \rgf_c1bus_wb[3]_i_19_n_0 ;
  wire \rgf_c1bus_wb[3]_i_20_n_0 ;
  wire \rgf_c1bus_wb[3]_i_21_n_0 ;
  wire \rgf_c1bus_wb[3]_i_22_n_0 ;
  wire \rgf_c1bus_wb[3]_i_2_n_0 ;
  wire \rgf_c1bus_wb[3]_i_3_n_0 ;
  wire \rgf_c1bus_wb[3]_i_4_n_0 ;
  wire \rgf_c1bus_wb[3]_i_5_n_0 ;
  wire \rgf_c1bus_wb[3]_i_6_n_0 ;
  wire \rgf_c1bus_wb[3]_i_7_n_0 ;
  wire \rgf_c1bus_wb[3]_i_8_n_0 ;
  wire \rgf_c1bus_wb[3]_i_9_n_0 ;
  wire \rgf_c1bus_wb[4]_i_10_n_0 ;
  wire \rgf_c1bus_wb[4]_i_11_n_0 ;
  wire \rgf_c1bus_wb[4]_i_12_n_0 ;
  wire \rgf_c1bus_wb[4]_i_13_n_0 ;
  wire \rgf_c1bus_wb[4]_i_14_n_0 ;
  wire \rgf_c1bus_wb[4]_i_15_n_0 ;
  wire \rgf_c1bus_wb[4]_i_16_n_0 ;
  wire \rgf_c1bus_wb[4]_i_17_n_0 ;
  wire \rgf_c1bus_wb[4]_i_2_n_0 ;
  wire \rgf_c1bus_wb[4]_i_3_n_0 ;
  wire \rgf_c1bus_wb[4]_i_4_n_0 ;
  wire \rgf_c1bus_wb[4]_i_5_n_0 ;
  wire \rgf_c1bus_wb[4]_i_6_n_0 ;
  wire \rgf_c1bus_wb[4]_i_7_n_0 ;
  wire \rgf_c1bus_wb[4]_i_8_n_0 ;
  wire \rgf_c1bus_wb[4]_i_9_n_0 ;
  wire \rgf_c1bus_wb[5]_i_10_n_0 ;
  wire \rgf_c1bus_wb[5]_i_11_n_0 ;
  wire \rgf_c1bus_wb[5]_i_12_n_0 ;
  wire \rgf_c1bus_wb[5]_i_13_n_0 ;
  wire \rgf_c1bus_wb[5]_i_14_n_0 ;
  wire \rgf_c1bus_wb[5]_i_15_n_0 ;
  wire \rgf_c1bus_wb[5]_i_16_n_0 ;
  wire \rgf_c1bus_wb[5]_i_17_n_0 ;
  wire \rgf_c1bus_wb[5]_i_18_n_0 ;
  wire \rgf_c1bus_wb[5]_i_19_n_0 ;
  wire \rgf_c1bus_wb[5]_i_2_n_0 ;
  wire \rgf_c1bus_wb[5]_i_3_n_0 ;
  wire \rgf_c1bus_wb[5]_i_4_n_0 ;
  wire \rgf_c1bus_wb[5]_i_5_n_0 ;
  wire \rgf_c1bus_wb[5]_i_6_n_0 ;
  wire \rgf_c1bus_wb[5]_i_7_n_0 ;
  wire \rgf_c1bus_wb[5]_i_8_n_0 ;
  wire \rgf_c1bus_wb[5]_i_9_n_0 ;
  wire \rgf_c1bus_wb[6]_i_10_n_0 ;
  wire \rgf_c1bus_wb[6]_i_11_n_0 ;
  wire \rgf_c1bus_wb[6]_i_12_n_0 ;
  wire \rgf_c1bus_wb[6]_i_13_n_0 ;
  wire \rgf_c1bus_wb[6]_i_14_n_0 ;
  wire \rgf_c1bus_wb[6]_i_15_n_0 ;
  wire \rgf_c1bus_wb[6]_i_16_n_0 ;
  wire \rgf_c1bus_wb[6]_i_17_n_0 ;
  wire \rgf_c1bus_wb[6]_i_18_n_0 ;
  wire \rgf_c1bus_wb[6]_i_2_n_0 ;
  wire \rgf_c1bus_wb[6]_i_3_n_0 ;
  wire \rgf_c1bus_wb[6]_i_4_n_0 ;
  wire \rgf_c1bus_wb[6]_i_5_n_0 ;
  wire \rgf_c1bus_wb[6]_i_6_n_0 ;
  wire \rgf_c1bus_wb[6]_i_7_n_0 ;
  wire \rgf_c1bus_wb[6]_i_8_n_0 ;
  wire \rgf_c1bus_wb[6]_i_9_n_0 ;
  wire \rgf_c1bus_wb[7]_i_10_n_0 ;
  wire \rgf_c1bus_wb[7]_i_11_n_0 ;
  wire \rgf_c1bus_wb[7]_i_12_n_0 ;
  wire \rgf_c1bus_wb[7]_i_13_n_0 ;
  wire \rgf_c1bus_wb[7]_i_14_n_0 ;
  wire \rgf_c1bus_wb[7]_i_15_n_0 ;
  wire \rgf_c1bus_wb[7]_i_16_n_0 ;
  wire \rgf_c1bus_wb[7]_i_17_n_0 ;
  wire \rgf_c1bus_wb[7]_i_18_n_0 ;
  wire \rgf_c1bus_wb[7]_i_19_n_0 ;
  wire \rgf_c1bus_wb[7]_i_20_n_0 ;
  wire \rgf_c1bus_wb[7]_i_21_n_0 ;
  wire \rgf_c1bus_wb[7]_i_22_n_0 ;
  wire \rgf_c1bus_wb[7]_i_2_n_0 ;
  wire \rgf_c1bus_wb[7]_i_3_n_0 ;
  wire \rgf_c1bus_wb[7]_i_4_n_0 ;
  wire \rgf_c1bus_wb[7]_i_5_n_0 ;
  wire \rgf_c1bus_wb[7]_i_6_n_0 ;
  wire \rgf_c1bus_wb[7]_i_7_n_0 ;
  wire \rgf_c1bus_wb[7]_i_8_n_0 ;
  wire \rgf_c1bus_wb[7]_i_9_n_0 ;
  wire \rgf_c1bus_wb[8]_i_10_n_0 ;
  wire \rgf_c1bus_wb[8]_i_11_n_0 ;
  wire \rgf_c1bus_wb[8]_i_12_n_0 ;
  wire \rgf_c1bus_wb[8]_i_13_n_0 ;
  wire \rgf_c1bus_wb[8]_i_14_n_0 ;
  wire \rgf_c1bus_wb[8]_i_15_n_0 ;
  wire \rgf_c1bus_wb[8]_i_16_n_0 ;
  wire \rgf_c1bus_wb[8]_i_17_n_0 ;
  wire \rgf_c1bus_wb[8]_i_18_n_0 ;
  wire \rgf_c1bus_wb[8]_i_19_n_0 ;
  wire \rgf_c1bus_wb[8]_i_20_n_0 ;
  wire \rgf_c1bus_wb[8]_i_2_n_0 ;
  wire \rgf_c1bus_wb[8]_i_3_n_0 ;
  wire \rgf_c1bus_wb[8]_i_4_n_0 ;
  wire \rgf_c1bus_wb[8]_i_5_n_0 ;
  wire \rgf_c1bus_wb[8]_i_6_n_0 ;
  wire \rgf_c1bus_wb[8]_i_7_n_0 ;
  wire \rgf_c1bus_wb[8]_i_8_n_0 ;
  wire \rgf_c1bus_wb[8]_i_9_n_0 ;
  wire \rgf_c1bus_wb[9]_i_10_n_0 ;
  wire \rgf_c1bus_wb[9]_i_11_n_0 ;
  wire \rgf_c1bus_wb[9]_i_12_n_0 ;
  wire \rgf_c1bus_wb[9]_i_13_n_0 ;
  wire \rgf_c1bus_wb[9]_i_14_n_0 ;
  wire \rgf_c1bus_wb[9]_i_15_n_0 ;
  wire \rgf_c1bus_wb[9]_i_16_n_0 ;
  wire \rgf_c1bus_wb[9]_i_17_n_0 ;
  wire \rgf_c1bus_wb[9]_i_18_n_0 ;
  wire \rgf_c1bus_wb[9]_i_19_n_0 ;
  wire \rgf_c1bus_wb[9]_i_20_n_0 ;
  wire \rgf_c1bus_wb[9]_i_21_n_0 ;
  wire \rgf_c1bus_wb[9]_i_22_n_0 ;
  wire \rgf_c1bus_wb[9]_i_23_n_0 ;
  wire \rgf_c1bus_wb[9]_i_2_n_0 ;
  wire \rgf_c1bus_wb[9]_i_3_n_0 ;
  wire \rgf_c1bus_wb[9]_i_4_n_0 ;
  wire \rgf_c1bus_wb[9]_i_5_n_0 ;
  wire \rgf_c1bus_wb[9]_i_6_n_0 ;
  wire \rgf_c1bus_wb[9]_i_7_n_0 ;
  wire \rgf_c1bus_wb[9]_i_8_n_0 ;
  wire \rgf_c1bus_wb[9]_i_9_n_0 ;
  wire \rgf_c1bus_wb_reg[0]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_1_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_33_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_34_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_1_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_9_n_0 ;
  wire rgf_selc0_stat_i_1_n_0;
  wire rgf_selc0_stat_i_2_n_0;
  wire \rgf_selc0_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_wb[0]_i_1_n_0 ;
  wire \rgf_selc0_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_wb[1]_i_25_n_0 ;
  wire \rgf_selc0_wb[1]_i_26_n_0 ;
  wire \rgf_selc0_wb[1]_i_27_n_0 ;
  wire \rgf_selc0_wb[1]_i_28_n_0 ;
  wire \rgf_selc0_wb[1]_i_29_n_0 ;
  wire \rgf_selc0_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_wb[1]_i_30_n_0 ;
  wire \rgf_selc0_wb[1]_i_31_n_0 ;
  wire \rgf_selc0_wb[1]_i_32_n_0 ;
  wire \rgf_selc0_wb[1]_i_33_n_0 ;
  wire \rgf_selc0_wb[1]_i_34_n_0 ;
  wire \rgf_selc0_wb[1]_i_35_n_0 ;
  wire \rgf_selc0_wb[1]_i_36_n_0 ;
  wire \rgf_selc0_wb[1]_i_37_n_0 ;
  wire \rgf_selc0_wb[1]_i_38_n_0 ;
  wire \rgf_selc0_wb[1]_i_39_n_0 ;
  wire \rgf_selc0_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_1_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_9_n_0 ;
  wire rgf_selc1_stat_i_1_n_0;
  wire rgf_selc1_stat_i_2_n_0;
  wire \rgf_selc1_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_wb[0]_i_1_n_0 ;
  wire \rgf_selc1_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_wb[1]_i_21_n_0 ;
  wire \rgf_selc1_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_wb[1]_i_25_n_0 ;
  wire \rgf_selc1_wb[1]_i_26_n_0 ;
  wire \rgf_selc1_wb[1]_i_27_n_0 ;
  wire \rgf_selc1_wb[1]_i_28_n_0 ;
  wire \rgf_selc1_wb[1]_i_29_n_0 ;
  wire \rgf_selc1_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_wb[1]_i_30_n_0 ;
  wire \rgf_selc1_wb[1]_i_31_n_0 ;
  wire \rgf_selc1_wb[1]_i_32_n_0 ;
  wire \rgf_selc1_wb[1]_i_33_n_0 ;
  wire \rgf_selc1_wb[1]_i_34_n_0 ;
  wire \rgf_selc1_wb[1]_i_35_n_0 ;
  wire \rgf_selc1_wb[1]_i_36_n_0 ;
  wire \rgf_selc1_wb[1]_i_37_n_0 ;
  wire \rgf_selc1_wb[1]_i_38_n_0 ;
  wire \rgf_selc1_wb[1]_i_39_n_0 ;
  wire \rgf_selc1_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_wb[1]_i_40_n_0 ;
  wire \rgf_selc1_wb[1]_i_41_n_0 ;
  wire \rgf_selc1_wb[1]_i_42_n_0 ;
  wire \rgf_selc1_wb[1]_i_43_n_0 ;
  wire \rgf_selc1_wb[1]_i_44_n_0 ;
  wire \rgf_selc1_wb[1]_i_45_n_0 ;
  wire \rgf_selc1_wb[1]_i_46_n_0 ;
  wire \rgf_selc1_wb[1]_i_47_n_0 ;
  wire \rgf_selc1_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_wb[1]_i_9_n_0 ;
  wire rst_n;
  wire \sp[0]_i_1_n_0 ;
  wire \sp[0]_i_2_n_0 ;
  wire \sp[10]_i_1_n_0 ;
  wire \sp[10]_i_2_n_0 ;
  wire \sp[11]_i_1_n_0 ;
  wire \sp[11]_i_2_n_0 ;
  wire \sp[12]_i_1_n_0 ;
  wire \sp[12]_i_2_n_0 ;
  wire \sp[13]_i_1_n_0 ;
  wire \sp[13]_i_2_n_0 ;
  wire \sp[14]_i_1_n_0 ;
  wire \sp[14]_i_2_n_0 ;
  wire \sp[15]_i_10_n_0 ;
  wire \sp[15]_i_11_n_0 ;
  wire \sp[15]_i_12_n_0 ;
  wire \sp[15]_i_14_n_0 ;
  wire \sp[15]_i_15_n_0 ;
  wire \sp[15]_i_16_n_0 ;
  wire \sp[15]_i_17_n_0 ;
  wire \sp[15]_i_18_n_0 ;
  wire \sp[15]_i_19_n_0 ;
  wire \sp[15]_i_1_n_0 ;
  wire \sp[15]_i_20_n_0 ;
  wire \sp[15]_i_21_n_0 ;
  wire \sp[15]_i_22_n_0 ;
  wire \sp[15]_i_23_n_0 ;
  wire \sp[15]_i_24_n_0 ;
  wire \sp[15]_i_25_n_0 ;
  wire \sp[15]_i_26_n_0 ;
  wire \sp[15]_i_2_n_0 ;
  wire \sp[15]_i_5_n_0 ;
  wire \sp[15]_i_6_n_0 ;
  wire \sp[15]_i_8_n_0 ;
  wire \sp[1]_i_1_n_0 ;
  wire \sp[1]_i_2_n_0 ;
  wire \sp[2]_i_1_n_0 ;
  wire \sp[2]_i_2_n_0 ;
  wire \sp[3]_i_1_n_0 ;
  wire \sp[3]_i_2_n_0 ;
  wire \sp[4]_i_1_n_0 ;
  wire \sp[4]_i_2_n_0 ;
  wire \sp[5]_i_1_n_0 ;
  wire \sp[5]_i_2_n_0 ;
  wire \sp[6]_i_1_n_0 ;
  wire \sp[6]_i_2_n_0 ;
  wire \sp[7]_i_1_n_0 ;
  wire \sp[7]_i_2_n_0 ;
  wire \sp[8]_i_1_n_0 ;
  wire \sp[8]_i_2_n_0 ;
  wire \sp[9]_i_1_n_0 ;
  wire \sp[9]_i_2_n_0 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[15]_i_7_n_1 ;
  wire \sp_reg[15]_i_7_n_2 ;
  wire \sp_reg[15]_i_7_n_3 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sr[11]_i_11_n_0 ;
  wire \sr[11]_i_12_n_0 ;
  wire \sr[11]_i_13_n_0 ;
  wire \sr[11]_i_14_n_0 ;
  wire \sr[11]_i_15_n_0 ;
  wire \sr[11]_i_2_n_0 ;
  wire \sr[11]_i_5_n_0 ;
  wire \sr[11]_i_9_n_0 ;
  wire \sr[13]_i_11_n_0 ;
  wire \sr[13]_i_12_n_0 ;
  wire \sr[13]_i_13_n_0 ;
  wire \sr[13]_i_14_n_0 ;
  wire \sr[13]_i_15_n_0 ;
  wire \sr[13]_i_16_n_0 ;
  wire \sr[13]_i_3_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire \sr[13]_i_5_n_0 ;
  wire \sr[13]_i_6_n_0 ;
  wire \sr[13]_i_7_n_0 ;
  wire \sr[13]_i_8_n_0 ;
  wire \sr[15]_i_2_n_0 ;
  wire \sr[15]_i_4_n_0 ;
  wire \sr[15]_i_6_n_0 ;
  wire \sr[15]_i_7_n_0 ;
  wire \sr[15]_i_8_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[3]_i_5_n_0 ;
  wire \sr[3]_i_6_n_0 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_11_n_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_14_n_0 ;
  wire \sr[4]_i_15_n_0 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_17_n_0 ;
  wire \sr[4]_i_18_n_0 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_25_n_0 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_29_n_0 ;
  wire \sr[4]_i_2_n_0 ;
  wire \sr[4]_i_30_n_0 ;
  wire \sr[4]_i_31_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_35_n_0 ;
  wire \sr[4]_i_36_n_0 ;
  wire \sr[4]_i_37_n_0 ;
  wire \sr[4]_i_38_n_0 ;
  wire \sr[4]_i_39_n_0 ;
  wire \sr[4]_i_3_n_0 ;
  wire \sr[4]_i_40_n_0 ;
  wire \sr[4]_i_41_n_0 ;
  wire \sr[4]_i_42_n_0 ;
  wire \sr[4]_i_43_n_0 ;
  wire \sr[4]_i_44_n_0 ;
  wire \sr[4]_i_45_n_0 ;
  wire \sr[4]_i_46_n_0 ;
  wire \sr[4]_i_47_n_0 ;
  wire \sr[4]_i_48_n_0 ;
  wire \sr[4]_i_49_n_0 ;
  wire \sr[4]_i_4_n_0 ;
  wire \sr[4]_i_50_n_0 ;
  wire \sr[4]_i_51_n_0 ;
  wire \sr[4]_i_52_n_0 ;
  wire \sr[4]_i_53_n_0 ;
  wire \sr[4]_i_54_n_0 ;
  wire \sr[4]_i_55_n_0 ;
  wire \sr[4]_i_56_n_0 ;
  wire \sr[4]_i_57_n_0 ;
  wire \sr[4]_i_58_n_0 ;
  wire \sr[4]_i_59_n_0 ;
  wire \sr[4]_i_5_n_0 ;
  wire \sr[4]_i_60_n_0 ;
  wire \sr[4]_i_61_n_0 ;
  wire \sr[4]_i_62_n_0 ;
  wire \sr[4]_i_63_n_0 ;
  wire \sr[4]_i_64_n_0 ;
  wire \sr[4]_i_65_n_0 ;
  wire \sr[4]_i_66_n_0 ;
  wire \sr[4]_i_67_n_0 ;
  wire \sr[4]_i_68_n_0 ;
  wire \sr[4]_i_69_n_0 ;
  wire \sr[4]_i_70_n_0 ;
  wire \sr[4]_i_71_n_0 ;
  wire \sr[4]_i_72_n_0 ;
  wire \sr[4]_i_73_n_0 ;
  wire \sr[4]_i_74_n_0 ;
  wire \sr[4]_i_75_n_0 ;
  wire \sr[4]_i_76_n_0 ;
  wire \sr[4]_i_77_n_0 ;
  wire \sr[4]_i_78_n_0 ;
  wire \sr[4]_i_79_n_0 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[4]_i_80_n_0 ;
  wire \sr[4]_i_81_n_0 ;
  wire \sr[4]_i_82_n_0 ;
  wire \sr[4]_i_83_n_0 ;
  wire \sr[4]_i_84_n_0 ;
  wire \sr[4]_i_85_n_0 ;
  wire \sr[4]_i_86_n_0 ;
  wire \sr[4]_i_87_n_0 ;
  wire \sr[4]_i_8_n_0 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_10_n_0 ;
  wire \sr[5]_i_11_n_0 ;
  wire \sr[5]_i_12_n_0 ;
  wire \sr[5]_i_2_n_0 ;
  wire \sr[5]_i_3_n_0 ;
  wire \sr[5]_i_4_n_0 ;
  wire \sr[5]_i_5_n_0 ;
  wire \sr[5]_i_7_n_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[5]_i_9_n_0 ;
  wire \sr[6]_i_10_n_0 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_12_n_0 ;
  wire \sr[6]_i_13_n_0 ;
  wire \sr[6]_i_14_n_0 ;
  wire \sr[6]_i_15_n_0 ;
  wire \sr[6]_i_16_n_0 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr[6]_i_18_n_0 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_20_n_0 ;
  wire \sr[6]_i_21_n_0 ;
  wire \sr[6]_i_22_n_0 ;
  wire \sr[6]_i_23_n_0 ;
  wire \sr[6]_i_24_n_0 ;
  wire \sr[6]_i_2_n_0 ;
  wire \sr[6]_i_4_n_0 ;
  wire \sr[6]_i_5_n_0 ;
  wire \sr[6]_i_6_n_0 ;
  wire \sr[6]_i_7_n_0 ;
  wire \sr[6]_i_8_n_0 ;
  wire \sr[6]_i_9_n_0 ;
  wire \sr[7]_i_2_n_0 ;
  wire \sr[7]_i_3_n_0 ;
  wire \sr[7]_i_5_n_0 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_7_n_0 ;
  wire \sr[7]_i_8_n_0 ;
  wire \sr[7]_i_9_n_0 ;
  wire \stat[0]_i_10__0_n_0 ;
  wire \stat[0]_i_10__1_n_0 ;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_11__0_n_0 ;
  wire \stat[0]_i_11__1_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12__0_n_0 ;
  wire \stat[0]_i_12__1_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13__0_n_0 ;
  wire \stat[0]_i_13__1_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14__0_n_0 ;
  wire \stat[0]_i_14__1_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15__0_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16__0_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_17__0_n_0 ;
  wire \stat[0]_i_17_n_0 ;
  wire \stat[0]_i_18__0_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_19__0_n_0 ;
  wire \stat[0]_i_19_n_0 ;
  wire \stat[0]_i_20__0_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21__0_n_0 ;
  wire \stat[0]_i_21_n_0 ;
  wire \stat[0]_i_22__0_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23__0_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24__0_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25__0_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26__0_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_27__0_n_0 ;
  wire \stat[0]_i_27_n_0 ;
  wire \stat[0]_i_28__0_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29__0_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2__0_n_0 ;
  wire \stat[0]_i_2__1_n_0 ;
  wire \stat[0]_i_2__2_n_0 ;
  wire \stat[0]_i_2_n_0 ;
  wire \stat[0]_i_30__0_n_0 ;
  wire \stat[0]_i_30_n_0 ;
  wire \stat[0]_i_31__0_n_0 ;
  wire \stat[0]_i_31_n_0 ;
  wire \stat[0]_i_32__0_n_0 ;
  wire \stat[0]_i_32_n_0 ;
  wire \stat[0]_i_33__0_n_0 ;
  wire \stat[0]_i_33_n_0 ;
  wire \stat[0]_i_34__0_n_0 ;
  wire \stat[0]_i_34_n_0 ;
  wire \stat[0]_i_35__0_n_0 ;
  wire \stat[0]_i_35_n_0 ;
  wire \stat[0]_i_36__0_n_0 ;
  wire \stat[0]_i_36_n_0 ;
  wire \stat[0]_i_37_n_0 ;
  wire \stat[0]_i_38_n_0 ;
  wire \stat[0]_i_3__0_n_0 ;
  wire \stat[0]_i_3__1_n_0 ;
  wire \stat[0]_i_3__2_n_0 ;
  wire \stat[0]_i_3_n_0 ;
  wire \stat[0]_i_4__0_n_0 ;
  wire \stat[0]_i_4__1_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5__0_n_0 ;
  wire \stat[0]_i_5__1_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6__0_n_0 ;
  wire \stat[0]_i_6__1_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7__0_n_0 ;
  wire \stat[0]_i_7__1_n_0 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8__0_n_0 ;
  wire \stat[0]_i_8__1_n_0 ;
  wire \stat[0]_i_8_n_0 ;
  wire \stat[0]_i_9__0_n_0 ;
  wire \stat[0]_i_9__1_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_10__0_n_0 ;
  wire \stat[1]_i_10_n_0 ;
  wire \stat[1]_i_11__0_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_12__0_n_0 ;
  wire \stat[1]_i_12_n_0 ;
  wire \stat[1]_i_13__0_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_14__0_n_0 ;
  wire \stat[1]_i_14_n_0 ;
  wire \stat[1]_i_15__0_n_0 ;
  wire \stat[1]_i_15_n_0 ;
  wire \stat[1]_i_16__0_n_0 ;
  wire \stat[1]_i_16_n_0 ;
  wire \stat[1]_i_17__0_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18__0_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_19__0_n_0 ;
  wire \stat[1]_i_19_n_0 ;
  wire \stat[1]_i_20__0_n_0 ;
  wire \stat[1]_i_20_n_0 ;
  wire \stat[1]_i_21_n_0 ;
  wire \stat[1]_i_22_n_0 ;
  wire \stat[1]_i_23_n_0 ;
  wire \stat[1]_i_24_n_0 ;
  wire \stat[1]_i_2__0_n_0 ;
  wire \stat[1]_i_2__1_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3__0_n_0 ;
  wire \stat[1]_i_3__1_n_0 ;
  wire \stat[1]_i_3_n_0 ;
  wire \stat[1]_i_4_n_0 ;
  wire \stat[1]_i_5__0_n_0 ;
  wire \stat[1]_i_5_n_0 ;
  wire \stat[1]_i_6_n_0 ;
  wire \stat[1]_i_7__0_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8__0_n_0 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[1]_i_9__0_n_0 ;
  wire \stat[1]_i_9_n_0 ;
  wire \stat[2]_i_10__0_n_0 ;
  wire \stat[2]_i_10_n_0 ;
  wire \stat[2]_i_11__0_n_0 ;
  wire \stat[2]_i_11_n_0 ;
  wire \stat[2]_i_12__0_n_0 ;
  wire \stat[2]_i_12_n_0 ;
  wire \stat[2]_i_13__0_n_0 ;
  wire \stat[2]_i_13_n_0 ;
  wire \stat[2]_i_14_n_0 ;
  wire \stat[2]_i_1__1_n_0 ;
  wire \stat[2]_i_2__1_n_0 ;
  wire \stat[2]_i_3__0_n_0 ;
  wire \stat[2]_i_3__1_n_0 ;
  wire \stat[2]_i_3_n_0 ;
  wire \stat[2]_i_4__0_n_0 ;
  wire \stat[2]_i_4_n_0 ;
  wire \stat[2]_i_5__0_n_0 ;
  wire \stat[2]_i_5_n_0 ;
  wire \stat[2]_i_6__0_n_0 ;
  wire \stat[2]_i_6_n_0 ;
  wire \stat[2]_i_7__0_n_0 ;
  wire \stat[2]_i_7_n_0 ;
  wire \stat[2]_i_8__0_n_0 ;
  wire \stat[2]_i_8_n_0 ;
  wire \stat[2]_i_9__0_n_0 ;
  wire \stat[2]_i_9_n_0 ;
  wire \stat_reg[1]_i_4__0_n_0 ;
  wire \stat_reg[1]_i_4_n_0 ;
  wire \stat_reg[1]_i_6_n_0 ;
  wire tout__1_carry__0_i_1__0_n_0;
  wire tout__1_carry__0_i_1_n_0;
  wire tout__1_carry__0_i_2__0_n_0;
  wire tout__1_carry__0_i_2_n_0;
  wire tout__1_carry__0_i_3__0_n_0;
  wire tout__1_carry__0_i_3_n_0;
  wire tout__1_carry__0_i_4__0_n_0;
  wire tout__1_carry__0_i_4_n_0;
  wire tout__1_carry__0_i_5__0_n_0;
  wire tout__1_carry__0_i_5_n_0;
  wire tout__1_carry__0_i_6__0_n_0;
  wire tout__1_carry__0_i_6_n_0;
  wire tout__1_carry__0_i_7__0_n_0;
  wire tout__1_carry__0_i_7_n_0;
  wire tout__1_carry__0_i_8__0_n_0;
  wire tout__1_carry__0_i_8_n_0;
  wire tout__1_carry__1_i_1__0_n_0;
  wire tout__1_carry__1_i_1_n_0;
  wire tout__1_carry__1_i_2__0_n_0;
  wire tout__1_carry__1_i_2_n_0;
  wire tout__1_carry__1_i_3__0_n_0;
  wire tout__1_carry__1_i_3_n_0;
  wire tout__1_carry__1_i_4__0_n_0;
  wire tout__1_carry__1_i_4_n_0;
  wire tout__1_carry__1_i_5__0_n_0;
  wire tout__1_carry__1_i_5_n_0;
  wire tout__1_carry__1_i_6__0_n_0;
  wire tout__1_carry__1_i_6_n_0;
  wire tout__1_carry__1_i_7__0_n_0;
  wire tout__1_carry__1_i_7_n_0;
  wire tout__1_carry__1_i_8__0_n_0;
  wire tout__1_carry__1_i_8_n_0;
  wire tout__1_carry__2_i_1__0_n_0;
  wire tout__1_carry__2_i_1_n_0;
  wire tout__1_carry__2_i_2__0_n_0;
  wire tout__1_carry__2_i_2_n_0;
  wire tout__1_carry__2_i_3__0_n_0;
  wire tout__1_carry__2_i_3_n_0;
  wire tout__1_carry__2_i_4__0_n_0;
  wire tout__1_carry__2_i_4_n_0;
  wire tout__1_carry__2_i_5__0_n_0;
  wire tout__1_carry__2_i_5_n_0;
  wire tout__1_carry__2_i_6__0_n_0;
  wire tout__1_carry__2_i_6_n_0;
  wire tout__1_carry__2_i_7__0_n_0;
  wire tout__1_carry__2_i_7_n_0;
  wire tout__1_carry__2_i_8__0_n_0;
  wire tout__1_carry__2_i_8_n_0;
  wire tout__1_carry__3_i_1__0_n_0;
  wire tout__1_carry__3_i_1_n_0;
  wire tout__1_carry__3_i_2__0_n_0;
  wire tout__1_carry__3_i_2_n_0;
  wire tout__1_carry__3_i_3__0_n_0;
  wire tout__1_carry__3_i_3_n_0;
  wire tout__1_carry_i_10__0_n_0;
  wire tout__1_carry_i_10_n_0;
  wire tout__1_carry_i_11__0_n_0;
  wire tout__1_carry_i_11_n_0;
  wire tout__1_carry_i_12__0_n_0;
  wire tout__1_carry_i_12_n_0;
  wire tout__1_carry_i_13__0_n_0;
  wire tout__1_carry_i_13_n_0;
  wire tout__1_carry_i_14_n_0;
  wire tout__1_carry_i_15_n_0;
  wire tout__1_carry_i_16_n_0;
  wire tout__1_carry_i_17_n_0;
  wire tout__1_carry_i_18_n_0;
  wire tout__1_carry_i_19_n_0;
  wire tout__1_carry_i_1__0_n_0;
  wire tout__1_carry_i_1_n_0;
  wire tout__1_carry_i_20_n_0;
  wire tout__1_carry_i_2__0_n_0;
  wire tout__1_carry_i_2_n_0;
  wire tout__1_carry_i_3__0_n_0;
  wire tout__1_carry_i_3_n_0;
  wire tout__1_carry_i_4__0_n_0;
  wire tout__1_carry_i_4_n_0;
  wire tout__1_carry_i_5__0_n_0;
  wire tout__1_carry_i_5_n_0;
  wire tout__1_carry_i_6__0_n_0;
  wire tout__1_carry_i_6_n_0;
  wire tout__1_carry_i_7__0_n_0;
  wire tout__1_carry_i_7_n_0;
  wire tout__1_carry_i_8__0_n_0;
  wire tout__1_carry_i_8_n_0;
  wire tout__1_carry_i_9__0_n_0;
  wire tout__1_carry_i_9_n_0;
  wire [3:0]\NLW_alu0/art/add/tout__1_carry__3_O_UNCONNECTED ;
  wire [3:0]\NLW_alu1/art/add/tout__1_carry__3_O_UNCONNECTED ;
  wire [3:0]\NLW_badr[3]_INST_0_i_29_O_UNCONNECTED ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[0]),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[10]),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[11]),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[12]),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[13]),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[14]),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[15]),
        .O(abus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[1]),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[2]),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[3]),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[4]),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[5]),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[6]),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[7]),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[8]),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[9]),
        .O(abus_o[9]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/art/add/tout__1_carry 
       (.CI(\<const0> ),
        .CO({\alu0/art/add/tout__1_carry_n_0 ,\alu0/art/add/tout__1_carry_n_1 ,\alu0/art/add/tout__1_carry_n_2 ,\alu0/art/add/tout__1_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry_i_1_n_0,tout__1_carry_i_2_n_0,tout__1_carry_i_3__0_n_0,\<const0> }),
        .O({\alu0/art/add/tout__1_carry_n_4 ,\alu0/art/add/tout__1_carry_n_5 ,\alu0/art/add/tout__1_carry_n_6 ,\alu0/art/add/tout__1_carry_n_7 }),
        .S({tout__1_carry_i_4_n_0,tout__1_carry_i_5_n_0,tout__1_carry_i_6_n_0,tout__1_carry_i_7__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/art/add/tout__1_carry__0 
       (.CI(\alu0/art/add/tout__1_carry_n_0 ),
        .CO({\alu0/art/add/tout__1_carry__0_n_0 ,\alu0/art/add/tout__1_carry__0_n_1 ,\alu0/art/add/tout__1_carry__0_n_2 ,\alu0/art/add/tout__1_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry__0_i_1_n_0,tout__1_carry__0_i_2_n_0,tout__1_carry__0_i_3_n_0,tout__1_carry__0_i_4_n_0}),
        .O({\alu0/art/add/tout__1_carry__0_n_4 ,\alu0/art/add/tout__1_carry__0_n_5 ,\alu0/art/add/tout__1_carry__0_n_6 ,\alu0/art/add/tout__1_carry__0_n_7 }),
        .S({tout__1_carry__0_i_5_n_0,tout__1_carry__0_i_6_n_0,tout__1_carry__0_i_7_n_0,tout__1_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/art/add/tout__1_carry__1 
       (.CI(\alu0/art/add/tout__1_carry__0_n_0 ),
        .CO({\alu0/art/add/tout__1_carry__1_n_0 ,\alu0/art/add/tout__1_carry__1_n_1 ,\alu0/art/add/tout__1_carry__1_n_2 ,\alu0/art/add/tout__1_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry__1_i_1_n_0,tout__1_carry__1_i_2_n_0,tout__1_carry__1_i_3_n_0,tout__1_carry__1_i_4_n_0}),
        .O({\alu0/art/add/tout__1_carry__1_n_4 ,\alu0/art/add/tout__1_carry__1_n_5 ,\alu0/art/add/tout__1_carry__1_n_6 ,\alu0/art/add/tout__1_carry__1_n_7 }),
        .S({tout__1_carry__1_i_5_n_0,tout__1_carry__1_i_6_n_0,tout__1_carry__1_i_7_n_0,tout__1_carry__1_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/art/add/tout__1_carry__2 
       (.CI(\alu0/art/add/tout__1_carry__1_n_0 ),
        .CO({\alu0/art/add/tout__1_carry__2_n_0 ,\alu0/art/add/tout__1_carry__2_n_1 ,\alu0/art/add/tout__1_carry__2_n_2 ,\alu0/art/add/tout__1_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry__2_i_1_n_0,tout__1_carry__2_i_2_n_0,tout__1_carry__2_i_3_n_0,tout__1_carry__2_i_4_n_0}),
        .O({\alu0/art/p_0_in ,\alu0/art/add/tout__1_carry__2_n_5 ,\alu0/art/add/tout__1_carry__2_n_6 ,\alu0/art/add/tout__1_carry__2_n_7 }),
        .S({tout__1_carry__2_i_5__0_n_0,tout__1_carry__2_i_6_n_0,tout__1_carry__2_i_7_n_0,tout__1_carry__2_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/art/add/tout__1_carry__3 
       (.CI(\alu0/art/add/tout__1_carry__2_n_0 ),
        .CO(\alu0/art/add/tout__1_carry__3_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,tout__1_carry__3_i_1_n_0}),
        .O({\alu0/art/add/tout ,\NLW_alu0/art/add/tout__1_carry__3_O_UNCONNECTED [0]}),
        .S({\<const0> ,\<const0> ,tout__1_carry__3_i_2__0_n_0,tout__1_carry__3_i_3__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/art/add/tout__1_carry 
       (.CI(\<const0> ),
        .CO({\alu1/art/add/tout__1_carry_n_0 ,\alu1/art/add/tout__1_carry_n_1 ,\alu1/art/add/tout__1_carry_n_2 ,\alu1/art/add/tout__1_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry_i_1__0_n_0,tout__1_carry_i_2__0_n_0,tout__1_carry_i_3_n_0,\<const0> }),
        .O({\alu1/art/add/tout__1_carry_n_4 ,\alu1/art/add/tout__1_carry_n_5 ,\alu1/art/add/tout__1_carry_n_6 ,\alu1/art/add/tout__1_carry_n_7 }),
        .S({tout__1_carry_i_4__0_n_0,tout__1_carry_i_5__0_n_0,tout__1_carry_i_6__0_n_0,tout__1_carry_i_7_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/art/add/tout__1_carry__0 
       (.CI(\alu1/art/add/tout__1_carry_n_0 ),
        .CO({\alu1/art/add/tout__1_carry__0_n_0 ,\alu1/art/add/tout__1_carry__0_n_1 ,\alu1/art/add/tout__1_carry__0_n_2 ,\alu1/art/add/tout__1_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry__0_i_1__0_n_0,tout__1_carry__0_i_2__0_n_0,tout__1_carry__0_i_3__0_n_0,tout__1_carry__0_i_4__0_n_0}),
        .O({\alu1/art/add/tout__1_carry__0_n_4 ,\alu1/art/add/tout__1_carry__0_n_5 ,\alu1/art/add/tout__1_carry__0_n_6 ,\alu1/art/add/tout__1_carry__0_n_7 }),
        .S({tout__1_carry__0_i_5__0_n_0,tout__1_carry__0_i_6__0_n_0,tout__1_carry__0_i_7__0_n_0,tout__1_carry__0_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/art/add/tout__1_carry__1 
       (.CI(\alu1/art/add/tout__1_carry__0_n_0 ),
        .CO({\alu1/art/add/tout__1_carry__1_n_0 ,\alu1/art/add/tout__1_carry__1_n_1 ,\alu1/art/add/tout__1_carry__1_n_2 ,\alu1/art/add/tout__1_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry__1_i_1__0_n_0,tout__1_carry__1_i_2__0_n_0,tout__1_carry__1_i_3__0_n_0,tout__1_carry__1_i_4__0_n_0}),
        .O({\alu1/art/add/tout__1_carry__1_n_4 ,\alu1/art/add/tout__1_carry__1_n_5 ,\alu1/art/add/tout__1_carry__1_n_6 ,\alu1/art/add/tout__1_carry__1_n_7 }),
        .S({tout__1_carry__1_i_5__0_n_0,tout__1_carry__1_i_6__0_n_0,tout__1_carry__1_i_7__0_n_0,tout__1_carry__1_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/art/add/tout__1_carry__2 
       (.CI(\alu1/art/add/tout__1_carry__1_n_0 ),
        .CO({\alu1/art/add/tout__1_carry__2_n_0 ,\alu1/art/add/tout__1_carry__2_n_1 ,\alu1/art/add/tout__1_carry__2_n_2 ,\alu1/art/add/tout__1_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({tout__1_carry__2_i_1__0_n_0,tout__1_carry__2_i_2__0_n_0,tout__1_carry__2_i_3__0_n_0,tout__1_carry__2_i_4__0_n_0}),
        .O({\alu1/art/p_0_in ,\alu1/art/add/tout__1_carry__2_n_5 ,\alu1/art/add/tout__1_carry__2_n_6 ,\alu1/art/add/tout__1_carry__2_n_7 }),
        .S({tout__1_carry__2_i_5_n_0,tout__1_carry__2_i_6__0_n_0,tout__1_carry__2_i_7__0_n_0,tout__1_carry__2_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/art/add/tout__1_carry__3 
       (.CI(\alu1/art/add/tout__1_carry__2_n_0 ),
        .CO(\alu1/art/add/tout__1_carry__3_n_3 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,tout__1_carry__3_i_1__0_n_0}),
        .O({\alu1/art/add/tout ,\NLW_alu1/art/add/tout__1_carry__3_O_UNCONNECTED [0]}),
        .S({\<const0> ,\<const0> ,tout__1_carry__3_i_2_n_0,tout__1_carry__3_i_3_n_0}));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[0]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[0]),
        .I3(a1bus_0[0]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[0]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[0]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [0]),
        .O(\badr[0]_INST_0_i_12_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[0]_INST_0_i_29 
       (.CI(\<const0> ),
        .CO({\badr[0]_INST_0_i_29_n_0 ,\badr[0]_INST_0_i_29_n_1 ,\badr[0]_INST_0_i_29_n_2 ,\badr[0]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/sptr/sp [1],\<const0> }),
        .O({\rgf/sptr/data2 [3:1],\rgf/sptr/data3 [0]}),
        .S({\rgf/sptr/sp [3:2],\badr[0]_INST_0_i_48_n_0 ,\rgf/sptr/sp [0]}));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [0]),
        .I5(\rgf/ivec/iv [0]),
        .O(\badr[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [0]),
        .O(\badr[0]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [0]),
        .O(\badr[0]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\badr[0]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [0]),
        .O(\badr[0]_INST_0_i_47_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[0]_INST_0_i_48 
       (.I0(\rgf/sptr/sp [1]),
        .O(\badr[0]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [0]),
        .O(\badr[0]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [0]),
        .O(\badr[0]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\badr[0]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [0]),
        .O(\badr[0]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[0]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [0]),
        .O(\badr[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [0]),
        .I5(\rgf/ivec/iv [0]),
        .O(\badr[0]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[10]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[10]),
        .I3(a1bus_0[10]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[10]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[10]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [10]),
        .O(\badr[10]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [10]),
        .I5(\rgf/ivec/iv [10]),
        .O(\badr[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [10]),
        .O(\badr[10]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [10]),
        .O(\badr[10]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [10]),
        .O(\badr[10]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [10]),
        .O(\badr[10]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [10]),
        .O(\badr[10]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [10]),
        .O(\badr[10]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [10]),
        .O(\badr[10]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [10]),
        .O(\badr[10]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[10]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [10]),
        .O(\badr[10]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [10]),
        .I5(\rgf/ivec/iv [10]),
        .O(\badr[10]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[11]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[11]),
        .I3(a1bus_0[11]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[11]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[11]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [11]),
        .O(\badr[11]_INST_0_i_12_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[11]_INST_0_i_29 
       (.CI(\badr[7]_INST_0_i_29_n_0 ),
        .CO({\badr[11]_INST_0_i_29_n_0 ,\badr[11]_INST_0_i_29_n_1 ,\badr[11]_INST_0_i_29_n_2 ,\badr[11]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [11:8]),
        .O(\rgf/sptr/data3 [11:8]),
        .S({\badr[11]_INST_0_i_48_n_0 ,\badr[11]_INST_0_i_49_n_0 ,\badr[11]_INST_0_i_50_n_0 ,\badr[11]_INST_0_i_51_n_0 }));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [11]),
        .I5(\rgf/ivec/iv [11]),
        .O(\badr[11]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [11]),
        .O(\badr[11]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [11]),
        .O(\badr[11]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [11]),
        .O(\badr[11]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [11]),
        .O(\badr[11]_INST_0_i_47_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_48 
       (.I0(\rgf/sptr/sp [11]),
        .O(\badr[11]_INST_0_i_48_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_49 
       (.I0(\rgf/sptr/sp [10]),
        .O(\badr[11]_INST_0_i_49_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_50 
       (.I0(\rgf/sptr/sp [9]),
        .O(\badr[11]_INST_0_i_50_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[11]_INST_0_i_51 
       (.I0(\rgf/sptr/sp [8]),
        .O(\badr[11]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [11]),
        .O(\badr[11]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [11]),
        .O(\badr[11]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_54 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [11]),
        .O(\badr[11]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_55 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [11]),
        .O(\badr[11]_INST_0_i_55_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[11]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [11]),
        .O(\badr[11]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [11]),
        .I5(\rgf/ivec/iv [11]),
        .O(\badr[11]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[12]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[12]),
        .I3(a1bus_0[12]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[12]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[12]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [12]),
        .O(\badr[12]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [12]),
        .I5(\rgf/ivec/iv [12]),
        .O(\badr[12]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [12]),
        .O(\badr[12]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [12]),
        .O(\badr[12]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [12]),
        .O(\badr[12]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [12]),
        .O(\badr[12]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [12]),
        .O(\badr[12]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [12]),
        .O(\badr[12]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [12]),
        .O(\badr[12]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [12]),
        .O(\badr[12]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[12]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [12]),
        .O(\badr[12]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [12]),
        .I5(\rgf/ivec/iv [12]),
        .O(\badr[12]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[13]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[13]),
        .I3(a1bus_0[13]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[13]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[13]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [13]),
        .O(\badr[13]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [13]),
        .I5(\rgf/ivec/iv [13]),
        .O(\badr[13]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [13]),
        .O(\badr[13]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [13]),
        .O(\badr[13]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [13]),
        .O(\badr[13]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [13]),
        .O(\badr[13]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [13]),
        .O(\badr[13]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [13]),
        .O(\badr[13]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [13]),
        .O(\badr[13]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [13]),
        .O(\badr[13]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[13]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [13]),
        .O(\badr[13]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [13]),
        .I5(\rgf/ivec/iv [13]),
        .O(\badr[13]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[14]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[14]),
        .I3(a1bus_0[14]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[14]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[14]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [14]),
        .O(\badr[14]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [14]),
        .I5(\rgf/ivec/iv [14]),
        .O(\badr[14]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [14]),
        .O(\badr[14]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [14]),
        .O(\badr[14]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [14]),
        .O(\badr[14]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [14]),
        .O(\badr[14]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [14]),
        .O(\badr[14]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [14]),
        .O(\badr[14]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [14]),
        .O(\badr[14]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [14]),
        .O(\badr[14]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[14]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [14]),
        .O(\badr[14]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [14]),
        .I5(\rgf/ivec/iv [14]),
        .O(\badr[14]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[15]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[15]),
        .I3(a1bus_0[15]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[15]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_104 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [15]),
        .O(\badr[15]_INST_0_i_104_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_105 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [15]),
        .O(\badr[15]_INST_0_i_105_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_108 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\badr[15]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_109 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [15]),
        .O(\badr[15]_INST_0_i_109_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_110 
       (.I0(\rgf/sptr/sp [15]),
        .O(\badr[15]_INST_0_i_110_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_111 
       (.I0(\rgf/sptr/sp [14]),
        .O(\badr[15]_INST_0_i_111_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_112 
       (.I0(\rgf/sptr/sp [13]),
        .O(\badr[15]_INST_0_i_112_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[15]_INST_0_i_113 
       (.I0(\rgf/sptr/sp [12]),
        .O(\badr[15]_INST_0_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4F4F4F4F4F4F4)) 
    \badr[15]_INST_0_i_114 
       (.I0(\badr[15]_INST_0_i_210_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I2(\badr[15]_INST_0_i_211_n_0 ),
        .I3(\badr[15]_INST_0_i_212_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .I5(\badr[15]_INST_0_i_213_n_0 ),
        .O(\badr[15]_INST_0_i_114_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[15]_INST_0_i_115 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat [1]),
        .I2(\ctl1/stat [0]),
        .O(\badr[15]_INST_0_i_115_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \badr[15]_INST_0_i_116 
       (.I0(\pc0[15]_i_3_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\bdatw[9]_INST_0_i_20_n_0 ),
        .I3(\badr[15]_INST_0_i_214_n_0 ),
        .I4(\badr[15]_INST_0_i_215_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_15_n_0 ),
        .O(\badr[15]_INST_0_i_116_n_0 ));
  LUT6 #(
    .INIT(64'h55555554FFFFFFFF)) 
    \badr[15]_INST_0_i_117 
       (.I0(\badr[15]_INST_0_i_216_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [10]),
        .I4(\badr[15]_INST_0_i_217_n_0 ),
        .I5(\bcmd[1]_INST_0_i_8_n_0 ),
        .O(\badr[15]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFD0FFFF)) 
    \badr[15]_INST_0_i_118 
       (.I0(\badr[15]_INST_0_i_218_n_0 ),
        .I1(\badr[15]_INST_0_i_219_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\badr[15]_INST_0_i_220_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\badr[15]_INST_0_i_221_n_0 ),
        .O(\badr[15]_INST_0_i_118_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA200AAAAAAAA)) 
    \badr[15]_INST_0_i_119 
       (.I0(\stat[2]_i_5__0_n_0 ),
        .I1(\badr[15]_INST_0_i_222_n_0 ),
        .I2(\badr[15]_INST_0_i_223_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I4(\badr[15]_INST_0_i_224_n_0 ),
        .I5(\badr[15]_INST_0_i_225_n_0 ),
        .O(ctl_sela1));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[15]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/sreg/sr [15]),
        .O(\badr[15]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFD00)) 
    \badr[15]_INST_0_i_120 
       (.I0(\badr[15]_INST_0_i_226_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I3(ctl_fetch1_fl_i_15_n_0),
        .I4(\fch/ir1 [13]),
        .I5(\ctl1/stat [0]),
        .O(\badr[15]_INST_0_i_120_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40444040)) 
    \badr[15]_INST_0_i_121 
       (.I0(\badr[15]_INST_0_i_227_n_0 ),
        .I1(\fch/ir1 [13]),
        .I2(\badr[15]_INST_0_i_142_n_0 ),
        .I3(\badr[15]_INST_0_i_228_n_0 ),
        .I4(\badr[15]_INST_0_i_229_n_0 ),
        .I5(\badr[15]_INST_0_i_230_n_0 ),
        .O(\badr[15]_INST_0_i_121_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_122 
       (.I0(\ctl1/stat [1]),
        .I1(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_122_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFDDD0000)) 
    \badr[15]_INST_0_i_123 
       (.I0(\badr[15]_INST_0_i_231_n_0 ),
        .I1(\badr[15]_INST_0_i_232_n_0 ),
        .I2(ctl_fetch1_fl_i_15_n_0),
        .I3(\badr[15]_INST_0_i_233_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I5(\badr[15]_INST_0_i_234_n_0 ),
        .O(\badr[15]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'h0000040054545454)) 
    \badr[15]_INST_0_i_140 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [1]),
        .I3(\bcmd[1]_INST_0_i_8_n_0 ),
        .I4(\badr[15]_INST_0_i_236_n_0 ),
        .I5(\badr[15]_INST_0_i_237_n_0 ),
        .O(\badr[15]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8A8A8AA)) 
    \badr[15]_INST_0_i_141 
       (.I0(\badr[15]_INST_0_i_238_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I2(\badr[15]_INST_0_i_239_n_0 ),
        .I3(\badr[15]_INST_0_i_240_n_0 ),
        .I4(\badr[15]_INST_0_i_241_n_0 ),
        .I5(\badr[15]_INST_0_i_242_n_0 ),
        .O(\badr[15]_INST_0_i_141_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_142 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [14]),
        .O(\badr[15]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAABAAAAAA)) 
    \badr[15]_INST_0_i_143 
       (.I0(\badr[15]_INST_0_i_243_n_0 ),
        .I1(\badr[15]_INST_0_i_244_n_0 ),
        .I2(\badr[15]_INST_0_i_245_n_0 ),
        .I3(\bdatw[9]_INST_0_i_20_n_0 ),
        .I4(\fch/ir1 [0]),
        .I5(\pc0[15]_i_3_n_0 ),
        .O(\badr[15]_INST_0_i_143_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_144 
       (.I0(\ctl1/stat [0]),
        .I1(\ctl1/stat [1]),
        .O(\badr[15]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'hFFBAFFBAFFFFFFBA)) 
    \badr[15]_INST_0_i_145 
       (.I0(\badr[15]_INST_0_i_246_n_0 ),
        .I1(\badr[15]_INST_0_i_247_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I3(\badr[15]_INST_0_i_248_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I5(\badr[15]_INST_0_i_249_n_0 ),
        .O(\badr[15]_INST_0_i_145_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \badr[15]_INST_0_i_146 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .I2(\bcmd[0]_INST_0_i_16_n_0 ),
        .I3(\fadr[15]_INST_0_i_21_n_0 ),
        .I4(\badr[15]_INST_0_i_215_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_15_n_0 ),
        .O(\badr[15]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'h04FFFFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_147 
       (.I0(\badr[15]_INST_0_i_250_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [14]),
        .O(\badr[15]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'h54FF545454FF54FF)) 
    \badr[15]_INST_0_i_148 
       (.I0(\badr[15]_INST_0_i_251_n_0 ),
        .I1(\badr[15]_INST_0_i_252_n_0 ),
        .I2(\badr[15]_INST_0_i_253_n_0 ),
        .I3(\badr[15]_INST_0_i_254_n_0 ),
        .I4(\badr[15]_INST_0_i_255_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_29_n_0 ),
        .O(\badr[15]_INST_0_i_148_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_28_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_159 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [15]),
        .O(\badr[15]_INST_0_i_159_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAFBAAAAAAAA)) 
    \badr[15]_INST_0_i_16 
       (.I0(\badr[15]_INST_0_i_62_n_0 ),
        .I1(\badr[15]_INST_0_i_63_n_0 ),
        .I2(\badr[15]_INST_0_i_64_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\badr[15]_INST_0_i_65_n_0 ),
        .I5(\bdatw[8]_INST_0_i_19_n_0 ),
        .O(ctl_sela0_rn[2]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_160 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [15]),
        .O(\badr[15]_INST_0_i_160_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_163 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\badr[15]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_164 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [15]),
        .O(\badr[15]_INST_0_i_164_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \badr[15]_INST_0_i_165 
       (.I0(\fch/ir0 [11]),
        .I1(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I2(\fch/ir0 [2]),
        .I3(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I4(\badr[15]_INST_0_i_256_n_0 ),
        .I5(\badr[15]_INST_0_i_257_n_0 ),
        .O(\badr[15]_INST_0_i_165_n_0 ));
  LUT4 #(
    .INIT(16'hFE7E)) 
    \badr[15]_INST_0_i_166 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [3]),
        .O(\badr[15]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8AAA802A822AA)) 
    \badr[15]_INST_0_i_167 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [3]),
        .O(\badr[15]_INST_0_i_167_n_0 ));
  LUT6 #(
    .INIT(64'hFBBBFBBBBBBBFBBB)) 
    \badr[15]_INST_0_i_168 
       (.I0(\badr[15]_INST_0_i_258_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\badr[15]_INST_0_i_259_n_0 ),
        .I3(\fch/ir0 [5]),
        .I4(\stat[1]_i_20_n_0 ),
        .I5(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_168_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AACCCAAA)) 
    \badr[15]_INST_0_i_169 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [8]),
        .I5(\stat[1]_i_24_n_0 ),
        .O(\badr[15]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAAAFE)) 
    \badr[15]_INST_0_i_17 
       (.I0(ctl_sela0),
        .I1(\badr[15]_INST_0_i_67_n_0 ),
        .I2(\badr[15]_INST_0_i_68_n_0 ),
        .I3(\badr[15]_INST_0_i_69_n_0 ),
        .I4(\badr[15]_INST_0_i_70_n_0 ),
        .I5(\ctl0/stat [2]),
        .O(\badr[15]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF404040)) 
    \badr[15]_INST_0_i_170 
       (.I0(\badr[15]_INST_0_i_260_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\badr[15]_INST_0_i_261_n_0 ),
        .I4(\stat[0]_i_26_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\badr[15]_INST_0_i_170_n_0 ));
  LUT6 #(
    .INIT(64'hFF02000000000000)) 
    \badr[15]_INST_0_i_171 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .I3(\badr[15]_INST_0_i_262_n_0 ),
        .I4(crdy),
        .I5(\fch/ir0 [5]),
        .O(\badr[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'h003AFF00000A0000)) 
    \badr[15]_INST_0_i_172 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [2]),
        .O(\badr[15]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \badr[15]_INST_0_i_173 
       (.I0(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I1(\stat[1]_i_24_n_0 ),
        .I2(\fch/ir0 [4]),
        .I3(\ccmd[2]_INST_0_i_5_n_0 ),
        .I4(\pc0[15]_i_3_n_0 ),
        .I5(\fadr[15]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_173_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010000)) 
    \badr[15]_INST_0_i_174 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I4(\badr[15]_INST_0_i_263_n_0 ),
        .I5(\badr[15]_INST_0_i_264_n_0 ),
        .O(\badr[15]_INST_0_i_174_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDDDFDDDD)) 
    \badr[15]_INST_0_i_175 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [9]),
        .I4(crdy),
        .I5(\fch/ir0 [8]),
        .O(\badr[15]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFDDDDF5FFD5D5)) 
    \badr[15]_INST_0_i_176 
       (.I0(\fch/ir0 [8]),
        .I1(\badr[15]_INST_0_i_265_n_0 ),
        .I2(\ctl0/stat [0]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\ccmd[4]_INST_0_i_17_n_0 ),
        .O(\badr[15]_INST_0_i_176_n_0 ));
  LUT5 #(
    .INIT(32'hCDCDCDCF)) 
    \badr[15]_INST_0_i_177 
       (.I0(\badr[15]_INST_0_i_266_n_0 ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [11]),
        .I4(crdy),
        .O(\badr[15]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'h2323333323233330)) 
    \badr[15]_INST_0_i_178 
       (.I0(\badr[15]_INST_0_i_267_n_0 ),
        .I1(\badr[15]_INST_0_i_268_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [9]),
        .I5(\badr[15]_INST_0_i_269_n_0 ),
        .O(\badr[15]_INST_0_i_178_n_0 ));
  LUT6 #(
    .INIT(64'h00040000FFFFFFFF)) 
    \badr[15]_INST_0_i_179 
       (.I0(\ccmd[2]_INST_0_i_5_n_0 ),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(\fch/ir0 [14]),
        .I3(\badr[15]_INST_0_i_270_n_0 ),
        .I4(\badr[15]_INST_0_i_271_n_0 ),
        .I5(\ctl0/stat [0]),
        .O(\badr[15]_INST_0_i_179_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_18 
       (.I0(\badr[15]_INST_0_i_28_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .O(\badr[15]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h84B44474FFFFFFFF)) 
    \badr[15]_INST_0_i_180 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [12]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\ccmd[2]_INST_0_i_15_n_0 ),
        .O(\badr[15]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'hDFFF5D33DFFF5D03)) 
    \badr[15]_INST_0_i_181 
       (.I0(crdy),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [3]),
        .I5(\pc0[15]_i_3_n_0 ),
        .O(\badr[15]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_182 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [12]),
        .I2(\ccmd[2]_INST_0_i_5_n_0 ),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [9]),
        .O(\badr[15]_INST_0_i_182_n_0 ));
  LUT6 #(
    .INIT(64'h470077D5FFFF77F7)) 
    \badr[15]_INST_0_i_183 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(crdy),
        .O(\badr[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'h000000000F0F0035)) 
    \badr[15]_INST_0_i_184 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [15]),
        .I5(\ctl0/stat [0]),
        .O(\badr[15]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \badr[15]_INST_0_i_185 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [3]),
        .I3(\badr[15]_INST_0_i_272_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [2]),
        .O(\badr[15]_INST_0_i_185_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_186 
       (.I0(\fch/ir0 [11]),
        .I1(\ctl0/stat [1]),
        .O(\badr[15]_INST_0_i_186_n_0 ));
  LUT4 #(
    .INIT(16'hFF10)) 
    \badr[15]_INST_0_i_187 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [13]),
        .I2(\ccmd[0]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_273_n_0 ),
        .O(\badr[15]_INST_0_i_187_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055FFF7FF)) 
    \badr[15]_INST_0_i_188 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [8]),
        .I2(crdy),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [9]),
        .I5(\ctl0/stat [0]),
        .O(\badr[15]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'h22222222222222A2)) 
    \badr[15]_INST_0_i_189 
       (.I0(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(\badr[15]_INST_0_i_274_n_0 ),
        .I3(\bdatw[15]_INST_0_i_154_n_0 ),
        .I4(\badr[15]_INST_0_i_275_n_0 ),
        .I5(\badr[15]_INST_0_i_276_n_0 ),
        .O(\badr[15]_INST_0_i_189_n_0 ));
  LUT5 #(
    .INIT(32'hDFDFDFFF)) 
    \badr[15]_INST_0_i_190 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [12]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir0 [14]),
        .O(\badr[15]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF000EFFFFFFFF)) 
    \badr[15]_INST_0_i_191 
       (.I0(\badr[15]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_68_n_0 ),
        .I2(\badr[15]_INST_0_i_69_n_0 ),
        .I3(\badr[15]_INST_0_i_70_n_0 ),
        .I4(\ctl0/stat [2]),
        .I5(ctl_sela0),
        .O(\badr[15]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'h00000000007F7F7F)) 
    \badr[15]_INST_0_i_192 
       (.I0(\badr[15]_INST_0_i_277_n_0 ),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(crdy),
        .I3(\badr[15]_INST_0_i_278_n_0 ),
        .I4(\stat[0]_i_26_n_0 ),
        .I5(\badr[15]_INST_0_i_279_n_0 ),
        .O(\badr[15]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'h7000000050000000)) 
    \badr[15]_INST_0_i_193 
       (.I0(\badr[15]_INST_0_i_280_n_0 ),
        .I1(\badr[15]_INST_0_i_281_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [11]),
        .I4(\badrx[15]_INST_0_i_4_n_0 ),
        .I5(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_193_n_0 ));
  LUT6 #(
    .INIT(64'h08AA080808080808)) 
    \badr[15]_INST_0_i_194 
       (.I0(\fch/ir0 [3]),
        .I1(\badr[15]_INST_0_i_282_n_0 ),
        .I2(\badr[15]_INST_0_i_283_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(crdy),
        .I5(\badr[15]_INST_0_i_262_n_0 ),
        .O(\badr[15]_INST_0_i_194_n_0 ));
  LUT6 #(
    .INIT(64'h00000000002A0000)) 
    \badr[15]_INST_0_i_195 
       (.I0(\badr[15]_INST_0_i_284_n_0 ),
        .I1(\badr[15]_INST_0_i_285_n_0 ),
        .I2(\ccmd[4]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [11]),
        .I5(\badr[15]_INST_0_i_286_n_0 ),
        .O(\badr[15]_INST_0_i_195_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFEFF)) 
    \badr[15]_INST_0_i_196 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [0]),
        .I4(\pc0[15]_i_3_n_0 ),
        .O(\badr[15]_INST_0_i_196_n_0 ));
  LUT5 #(
    .INIT(32'hBF0F0F0F)) 
    \badr[15]_INST_0_i_197 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [12]),
        .O(\badr[15]_INST_0_i_197_n_0 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \badr[15]_INST_0_i_198 
       (.I0(\fadr[15]_INST_0_i_14_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [10]),
        .I5(\rgf_selc0_rn_wb[0]_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_198_n_0 ));
  LUT6 #(
    .INIT(64'hDDDD0DDDFFFFFFFF)) 
    \badr[15]_INST_0_i_199 
       (.I0(\badr[15]_INST_0_i_257_n_0 ),
        .I1(\badr[15]_INST_0_i_256_n_0 ),
        .I2(\stat[0]_i_8__1_n_0 ),
        .I3(\badr[15]_INST_0_i_287_n_0 ),
        .I4(\fch/ir0 [6]),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_199_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF1FF)) 
    \badr[15]_INST_0_i_200 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [15]),
        .I3(\ctl0/stat [0]),
        .I4(\ctl0/stat [1]),
        .O(\badr[15]_INST_0_i_200_n_0 ));
  LUT6 #(
    .INIT(64'h8088808080808080)) 
    \badr[15]_INST_0_i_201 
       (.I0(\fch/ir0 [1]),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I3(\badr[15]_INST_0_i_256_n_0 ),
        .I4(\stat[2]_i_10_n_0 ),
        .I5(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_201_n_0 ));
  LUT3 #(
    .INIT(8'h8E)) 
    \badr[15]_INST_0_i_202 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [0]),
        .O(\badr[15]_INST_0_i_202_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \badr[15]_INST_0_i_203 
       (.I0(\ccmd[2]_INST_0_i_5_n_0 ),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [14]),
        .O(\badr[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'h202AAAAAAAAAAAAA)) 
    \badr[15]_INST_0_i_204 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [8]),
        .O(\badr[15]_INST_0_i_204_n_0 ));
  LUT6 #(
    .INIT(64'h5FFFFFFF7F7F7F7F)) 
    \badr[15]_INST_0_i_205 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(crdy),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [8]),
        .O(\badr[15]_INST_0_i_205_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F700F200)) 
    \badr[15]_INST_0_i_206 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [11]),
        .I4(\badr[15]_INST_0_i_288_n_0 ),
        .I5(\badr[15]_INST_0_i_289_n_0 ),
        .O(\badr[15]_INST_0_i_206_n_0 ));
  LUT4 #(
    .INIT(16'h1011)) 
    \badr[15]_INST_0_i_207 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\badr[15]_INST_0_i_290_n_0 ),
        .I3(crdy),
        .O(\badr[15]_INST_0_i_207_n_0 ));
  LUT6 #(
    .INIT(64'h5D5D0C0CFF5D0C0C)) 
    \badr[15]_INST_0_i_208 
       (.I0(\badr[15]_INST_0_i_291_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I2(\badr[15]_INST_0_i_292_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\stat[2]_i_10_n_0 ),
        .I5(\badr[15]_INST_0_i_293_n_0 ),
        .O(\badr[15]_INST_0_i_208_n_0 ));
  LUT6 #(
    .INIT(64'hDF00DFDFDFDFDFDF)) 
    \badr[15]_INST_0_i_210 
       (.I0(\badr[15]_INST_0_i_294_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\bcmd[0]_INST_0_i_23_n_0 ),
        .I3(\badr[15]_INST_0_i_295_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I5(\fch/ir1 [2]),
        .O(\badr[15]_INST_0_i_210_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \badr[15]_INST_0_i_211 
       (.I0(\rgf_selc1_rn_wb[0]_i_24_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\badr[15]_INST_0_i_296_n_0 ),
        .I3(\badr[15]_INST_0_i_297_n_0 ),
        .I4(\bdatw[9]_INST_0_i_65_n_0 ),
        .I5(\badr[15]_INST_0_i_298_n_0 ),
        .O(\badr[15]_INST_0_i_211_n_0 ));
  LUT4 #(
    .INIT(16'h7F77)) 
    \badr[15]_INST_0_i_212 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_212_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_213 
       (.I0(\fch/ir1 [10]),
        .I1(\ctl1/stat [1]),
        .O(\badr[15]_INST_0_i_213_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_214 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_214_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_215 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [4]),
        .O(\badr[15]_INST_0_i_215_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEA00C0)) 
    \badr[15]_INST_0_i_216 
       (.I0(\badr[15]_INST_0_i_299_n_0 ),
        .I1(\badr[15]_INST_0_i_300_n_0 ),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_216_n_0 ));
  LUT6 #(
    .INIT(64'hAAEE00E0BBFF0BFF)) 
    \badr[15]_INST_0_i_217 
       (.I0(\badr[15]_INST_0_i_301_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [2]),
        .I4(\fadr[15]_INST_0_i_21_n_0 ),
        .I5(\fch/ir1 [5]),
        .O(\badr[15]_INST_0_i_217_n_0 ));
  LUT6 #(
    .INIT(64'hEE1EFE5FFFFFFFFF)) 
    \badr[15]_INST_0_i_218 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [2]),
        .I5(\badr[15]_INST_0_i_302_n_0 ),
        .O(\badr[15]_INST_0_i_218_n_0 ));
  LUT6 #(
    .INIT(64'h0400FFFF04000400)) 
    \badr[15]_INST_0_i_219 
       (.I0(\badr[15]_INST_0_i_303_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [2]),
        .I4(\badr[15]_INST_0_i_304_n_0 ),
        .I5(\fch/ir1 [5]),
        .O(\badr[15]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'h0000EF4000000000)) 
    \badr[15]_INST_0_i_220 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_220_n_0 ));
  LUT6 #(
    .INIT(64'h3303332030001300)) 
    \badr[15]_INST_0_i_221 
       (.I0(\fch/ir1 [6]),
        .I1(\fadr[15]_INST_0_i_21_n_0 ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [2]),
        .O(\badr[15]_INST_0_i_221_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDFFFDFFFD5F5)) 
    \badr[15]_INST_0_i_222 
       (.I0(\bcmd[0]_INST_0_i_23_n_0 ),
        .I1(\badr[15]_INST_0_i_305_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\ctl1/stat [0]),
        .I5(\badr[15]_INST_0_i_306_n_0 ),
        .O(\badr[15]_INST_0_i_222_n_0 ));
  LUT6 #(
    .INIT(64'h00F011F1FFFF11F1)) 
    \badr[15]_INST_0_i_223 
       (.I0(\badr[15]_INST_0_i_307_n_0 ),
        .I1(\badr[15]_INST_0_i_308_n_0 ),
        .I2(\badr[15]_INST_0_i_309_n_0 ),
        .I3(\badr[15]_INST_0_i_310_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_10_n_0 ),
        .I5(\badr[15]_INST_0_i_311_n_0 ),
        .O(\badr[15]_INST_0_i_223_n_0 ));
  LUT6 #(
    .INIT(64'h000000800000F030)) 
    \badr[15]_INST_0_i_224 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [13]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [12]),
        .O(\badr[15]_INST_0_i_224_n_0 ));
  LUT6 #(
    .INIT(64'h55555555DDD0DDDD)) 
    \badr[15]_INST_0_i_225 
       (.I0(\badr[15]_INST_0_i_312_n_0 ),
        .I1(\fch/ir1 [13]),
        .I2(\bdatw[15]_INST_0_i_208_n_0 ),
        .I3(\stat[2]_i_13_n_0 ),
        .I4(\fch_irq_lev[1]_i_5_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_225_n_0 ));
  LUT5 #(
    .INIT(32'h3131A2B2)) 
    \badr[15]_INST_0_i_226 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [0]),
        .I3(\pc0[15]_i_3_n_0 ),
        .I4(\fch/ir1 [1]),
        .O(\badr[15]_INST_0_i_226_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF5555F0F04540)) 
    \badr[15]_INST_0_i_227 
       (.I0(\fch/ir1 [14]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [6]),
        .I4(\fch/ir1 [15]),
        .I5(\ctl1/stat [0]),
        .O(\badr[15]_INST_0_i_227_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2AAAFFFFFFFF)) 
    \badr[15]_INST_0_i_228 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [12]),
        .O(\badr[15]_INST_0_i_228_n_0 ));
  LUT6 #(
    .INIT(64'hF232E2BAE2BAE2BA)) 
    \badr[15]_INST_0_i_229 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_229_n_0 ));
  LUT6 #(
    .INIT(64'h0202020202FF0202)) 
    \badr[15]_INST_0_i_230 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [13]),
        .I3(\badr[15]_INST_0_i_313_n_0 ),
        .I4(\fch_irq_lev[1]_i_5_n_0 ),
        .I5(\stat[2]_i_13_n_0 ),
        .O(\badr[15]_INST_0_i_230_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01005555)) 
    \badr[15]_INST_0_i_231 
       (.I0(\badr[15]_INST_0_i_314_n_0 ),
        .I1(\badr[15]_INST_0_i_315_n_0 ),
        .I2(\badr[15]_INST_0_i_316_n_0 ),
        .I3(\badr[15]_INST_0_i_317_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I5(\badr[15]_INST_0_i_318_n_0 ),
        .O(\badr[15]_INST_0_i_231_n_0 ));
  LUT6 #(
    .INIT(64'h003F000200FF0002)) 
    \badr[15]_INST_0_i_232 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [13]),
        .O(\badr[15]_INST_0_i_232_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[15]_INST_0_i_233 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [13]),
        .O(\badr[15]_INST_0_i_233_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \badr[15]_INST_0_i_234 
       (.I0(\badr[15]_INST_0_i_319_n_0 ),
        .I1(\badr[15]_INST_0_i_320_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I3(\fch_irq_lev[1]_i_4_n_0 ),
        .I4(\badr[15]_INST_0_i_321_n_0 ),
        .I5(\badr[15]_INST_0_i_252_n_0 ),
        .O(\badr[15]_INST_0_i_234_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00F2FFFFFFFF)) 
    \badr[15]_INST_0_i_235 
       (.I0(\badr[15]_INST_0_i_120_n_0 ),
        .I1(\badr[15]_INST_0_i_121_n_0 ),
        .I2(\badr[15]_INST_0_i_122_n_0 ),
        .I3(\badr[15]_INST_0_i_123_n_0 ),
        .I4(\ctl1/stat [2]),
        .I5(ctl_sela1),
        .O(\badr[15]_INST_0_i_235_n_0 ));
  LUT6 #(
    .INIT(64'hBBB0BBBBFFFFFFFF)) 
    \badr[15]_INST_0_i_236 
       (.I0(\fch/ir1 [6]),
        .I1(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I2(\bcmd[0]_INST_0_i_7_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [0]),
        .O(\badr[15]_INST_0_i_236_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    \badr[15]_INST_0_i_237 
       (.I0(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\bdatw[9]_INST_0_i_65_n_0 ),
        .I3(\badr[15]_INST_0_i_297_n_0 ),
        .I4(\badr[15]_INST_0_i_296_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_237_n_0 ));
  LUT5 #(
    .INIT(32'hEABFBFEA)) 
    \badr[15]_INST_0_i_238 
       (.I0(\fch/ir1 [13]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_238_n_0 ));
  LUT6 #(
    .INIT(64'h0000000D000D000D)) 
    \badr[15]_INST_0_i_239 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\badr[15]_INST_0_i_322_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\badr[15]_INST_0_i_323_n_0 ),
        .I4(\badr[15]_INST_0_i_299_n_0 ),
        .I5(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_239_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2000AAAAA0A0)) 
    \badr[15]_INST_0_i_240 
       (.I0(\fch/ir1 [10]),
        .I1(\badr[15]_INST_0_i_324_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I3(\fch/ir1 [7]),
        .I4(\badr[15]_INST_0_i_325_n_0 ),
        .I5(\badr[15]_INST_0_i_326_n_0 ),
        .O(\badr[15]_INST_0_i_240_n_0 ));
  LUT6 #(
    .INIT(64'h45404444FFFFFFFF)) 
    \badr[15]_INST_0_i_241 
       (.I0(\badr[15]_INST_0_i_327_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_241_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2B8E2F0)) 
    \badr[15]_INST_0_i_242 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [6]),
        .I5(\fadr[15]_INST_0_i_21_n_0 ),
        .O(\badr[15]_INST_0_i_242_n_0 ));
  LUT6 #(
    .INIT(64'hC000C5C5C000C505)) 
    \badr[15]_INST_0_i_243 
       (.I0(\stat[0]_i_22_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [15]),
        .I3(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_243_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[15]_INST_0_i_244 
       (.I0(\bcmd[0]_INST_0_i_16_n_0 ),
        .I1(\fadr[15]_INST_0_i_21_n_0 ),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [5]),
        .O(\badr[15]_INST_0_i_244_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_245 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [13]),
        .O(\badr[15]_INST_0_i_245_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \badr[15]_INST_0_i_246 
       (.I0(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\badr[15]_INST_0_i_296_n_0 ),
        .I3(\badr[15]_INST_0_i_297_n_0 ),
        .I4(\bdatw[9]_INST_0_i_65_n_0 ),
        .I5(\badr[15]_INST_0_i_298_n_0 ),
        .O(\badr[15]_INST_0_i_246_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFDFCFFFDFFFF)) 
    \badr[15]_INST_0_i_247 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [15]),
        .I2(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [2]),
        .O(\badr[15]_INST_0_i_247_n_0 ));
  LUT6 #(
    .INIT(64'hF200000000000000)) 
    \badr[15]_INST_0_i_248 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [14]),
        .I2(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I3(\badr[15]_INST_0_i_144_n_0 ),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_248_n_0 ));
  LUT6 #(
    .INIT(64'hBBB0BBBBFFFFFFFF)) 
    \badr[15]_INST_0_i_249 
       (.I0(\fch/ir1 [6]),
        .I1(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I2(\bcmd[0]_INST_0_i_7_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [1]),
        .O(\badr[15]_INST_0_i_249_n_0 ));
  LUT6 #(
    .INIT(64'hFF24DB00FF708F00)) 
    \badr[15]_INST_0_i_250 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_250_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEA00C0)) 
    \badr[15]_INST_0_i_251 
       (.I0(\badr[15]_INST_0_i_299_n_0 ),
        .I1(\badr[15]_INST_0_i_300_n_0 ),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_251_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[15]_INST_0_i_252 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_252_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFE0E0F0FFEFEF)) 
    \badr[15]_INST_0_i_253 
       (.I0(\badr[15]_INST_0_i_328_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [4]),
        .O(\badr[15]_INST_0_i_253_n_0 ));
  LUT6 #(
    .INIT(64'hC0E0FFFFC0E0C0E0)) 
    \badr[15]_INST_0_i_254 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_302_n_0 ),
        .I3(\bcmd[0]_INST_0_i_7_n_0 ),
        .I4(\stat[0]_i_30__0_n_0 ),
        .I5(\badr[15]_INST_0_i_329_n_0 ),
        .O(\badr[15]_INST_0_i_254_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF7BBFFF7FFB)) 
    \badr[15]_INST_0_i_255 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_255_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \badr[15]_INST_0_i_256 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [3]),
        .O(\badr[15]_INST_0_i_256_n_0 ));
  LUT5 #(
    .INIT(32'h80000000)) 
    \badr[15]_INST_0_i_257 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_257_n_0 ));
  LUT6 #(
    .INIT(64'h4040404044400040)) 
    \badr[15]_INST_0_i_258 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_258_n_0 ));
  LUT4 #(
    .INIT(16'h4044)) 
    \badr[15]_INST_0_i_259 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(crdy),
        .I3(\fch/ir0 [8]),
        .O(\badr[15]_INST_0_i_259_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \badr[15]_INST_0_i_260 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [2]),
        .O(\badr[15]_INST_0_i_260_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_261 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_261_n_0 ));
  LUT5 #(
    .INIT(32'h44040404)) 
    \badr[15]_INST_0_i_262 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_262_n_0 ));
  LUT6 #(
    .INIT(64'h2A022A022A020000)) 
    \badr[15]_INST_0_i_263 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .I4(crdy),
        .I5(\ctl0/stat [0]),
        .O(\badr[15]_INST_0_i_263_n_0 ));
  LUT6 #(
    .INIT(64'h0440444400440444)) 
    \badr[15]_INST_0_i_264 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [11]),
        .O(\badr[15]_INST_0_i_264_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \badr[15]_INST_0_i_265 
       (.I0(\fch/ir0 [6]),
        .I1(\ctl0/stat [0]),
        .I2(\fch/ir0 [9]),
        .O(\badr[15]_INST_0_i_265_n_0 ));
  LUT6 #(
    .INIT(64'h4545C5554155C555)) 
    \badr[15]_INST_0_i_266 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_266_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFD6FFFFF7EE)) 
    \badr[15]_INST_0_i_267 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_267_n_0 ));
  LUT6 #(
    .INIT(64'h0040FFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_268 
       (.I0(\ctl0/stat [0]),
        .I1(crdy),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\badr[15]_INST_0_i_268_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_269 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_269_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF0D0000)) 
    \badr[15]_INST_0_i_27 
       (.I0(\badr[15]_INST_0_i_87_n_0 ),
        .I1(\badr[15]_INST_0_i_88_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .I3(\badr[15]_INST_0_i_89_n_0 ),
        .I4(\bdatw[8]_INST_0_i_19_n_0 ),
        .I5(\badr[15]_INST_0_i_90_n_0 ),
        .O(ctl_sela0_rn[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_270 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [15]),
        .O(\badr[15]_INST_0_i_270_n_0 ));
  LUT4 #(
    .INIT(16'h2B22)) 
    \badr[15]_INST_0_i_271 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [2]),
        .O(\badr[15]_INST_0_i_271_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_272 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_272_n_0 ));
  LUT6 #(
    .INIT(64'h03000F000F020F02)) 
    \badr[15]_INST_0_i_273 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\fch/ir0 [12]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [14]),
        .O(\badr[15]_INST_0_i_273_n_0 ));
  LUT6 #(
    .INIT(64'hFFFCFDDCFFFFFFFC)) 
    \badr[15]_INST_0_i_274 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [6]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_274_n_0 ));
  LUT6 #(
    .INIT(64'h1000100010000000)) 
    \badr[15]_INST_0_i_275 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [5]),
        .O(\badr[15]_INST_0_i_275_n_0 ));
  LUT4 #(
    .INIT(16'h4004)) 
    \badr[15]_INST_0_i_276 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_276_n_0 ));
  LUT6 #(
    .INIT(64'h3272767210501050)) 
    \badr[15]_INST_0_i_277 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [0]),
        .O(\badr[15]_INST_0_i_277_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_278 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_278_n_0 ));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    \badr[15]_INST_0_i_279 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [3]),
        .O(\badr[15]_INST_0_i_279_n_0 ));
  LUT6 #(
    .INIT(64'h5454545544444444)) 
    \badr[15]_INST_0_i_28 
       (.I0(\ctl0/stat [2]),
        .I1(\badr[15]_INST_0_i_91_n_0 ),
        .I2(\badr[15]_INST_0_i_92_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\badr[15]_INST_0_i_93_n_0 ),
        .I5(\ccmd[4]_INST_0_i_8_n_0 ),
        .O(\badr[15]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFBBF7FFFFB)) 
    \badr[15]_INST_0_i_280 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [3]),
        .O(\badr[15]_INST_0_i_280_n_0 ));
  LUT5 #(
    .INIT(32'hCFCFFFF1)) 
    \badr[15]_INST_0_i_281 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [5]),
        .O(\badr[15]_INST_0_i_281_n_0 ));
  LUT5 #(
    .INIT(32'h08000808)) 
    \badr[15]_INST_0_i_282 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(crdy),
        .I4(\fch/ir0 [8]),
        .O(\badr[15]_INST_0_i_282_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[15]_INST_0_i_283 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .O(\badr[15]_INST_0_i_283_n_0 ));
  LUT5 #(
    .INIT(32'hEF2FFF0F)) 
    \badr[15]_INST_0_i_284 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [8]),
        .O(\badr[15]_INST_0_i_284_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \badr[15]_INST_0_i_285 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [0]),
        .O(\badr[15]_INST_0_i_285_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000407F)) 
    \badr[15]_INST_0_i_286 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [8]),
        .O(\badr[15]_INST_0_i_286_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \badr[15]_INST_0_i_287 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .O(\badr[15]_INST_0_i_287_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \badr[15]_INST_0_i_288 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [1]),
        .O(\badr[15]_INST_0_i_288_n_0 ));
  LUT6 #(
    .INIT(64'hF3F50070C0A00070)) 
    \badr[15]_INST_0_i_289 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [1]),
        .O(\badr[15]_INST_0_i_289_n_0 ));
  LUT6 #(
    .INIT(64'hF800FD0FFAF0FFFF)) 
    \badr[15]_INST_0_i_290 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [1]),
        .O(\badr[15]_INST_0_i_290_n_0 ));
  LUT6 #(
    .INIT(64'hFDF7FFFFFE7EFFFF)) 
    \badr[15]_INST_0_i_291 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [7]),
        .O(\badr[15]_INST_0_i_291_n_0 ));
  LUT5 #(
    .INIT(32'h00F0FBFB)) 
    \badr[15]_INST_0_i_292 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(crdy),
        .I4(\fch/ir0 [4]),
        .O(\badr[15]_INST_0_i_292_n_0 ));
  LUT5 #(
    .INIT(32'h0FFFFFFB)) 
    \badr[15]_INST_0_i_293 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [3]),
        .O(\badr[15]_INST_0_i_293_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_294 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_294_n_0 ));
  LUT6 #(
    .INIT(64'hFFBF00000000FFFF)) 
    \badr[15]_INST_0_i_295 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_295_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_296 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_296_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_297 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_297_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \badr[15]_INST_0_i_298 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [13]),
        .O(\badr[15]_INST_0_i_298_n_0 ));
  LUT5 #(
    .INIT(32'h44040404)) 
    \badr[15]_INST_0_i_299 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_299_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [15]),
        .I5(\rgf/ivec/iv [15]),
        .O(\badr[15]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_300 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_300_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF8CFFFF)) 
    \badr[15]_INST_0_i_301 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_301_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[15]_INST_0_i_302 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_302_n_0 ));
  LUT4 #(
    .INIT(16'hFE7E)) 
    \badr[15]_INST_0_i_303 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_303_n_0 ));
  LUT4 #(
    .INIT(16'hAABA)) 
    \badr[15]_INST_0_i_304 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .O(\badr[15]_INST_0_i_304_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFBFEFFFFF67E)) 
    \badr[15]_INST_0_i_305 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [7]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_305_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[15]_INST_0_i_306 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_306_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5CCC)) 
    \badr[15]_INST_0_i_307 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [10]),
        .O(\badr[15]_INST_0_i_307_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0D00000E00000)) 
    \badr[15]_INST_0_i_308 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_308_n_0 ));
  LUT4 #(
    .INIT(16'hF80F)) 
    \badr[15]_INST_0_i_309 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_309_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \badr[15]_INST_0_i_310 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [11]),
        .O(\badr[15]_INST_0_i_310_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \badr[15]_INST_0_i_311 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .O(\badr[15]_INST_0_i_311_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \badr[15]_INST_0_i_312 
       (.I0(\fch/ir1 [14]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [15]),
        .O(\badr[15]_INST_0_i_312_n_0 ));
  LUT5 #(
    .INIT(32'hDF0FFFDF)) 
    \badr[15]_INST_0_i_313 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [0]),
        .O(\badr[15]_INST_0_i_313_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F2FFF0FFF0FFF)) 
    \badr[15]_INST_0_i_314 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [10]),
        .O(\badr[15]_INST_0_i_314_n_0 ));
  LUT6 #(
    .INIT(64'h1110000000000000)) 
    \badr[15]_INST_0_i_315 
       (.I0(\fch/ir1 [3]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [4]),
        .O(\badr[15]_INST_0_i_315_n_0 ));
  LUT5 #(
    .INIT(32'h1111D311)) 
    \badr[15]_INST_0_i_316 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [7]),
        .I4(\ctl1/stat [0]),
        .O(\badr[15]_INST_0_i_316_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDFFFDFFF0C)) 
    \badr[15]_INST_0_i_317 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [4]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [6]),
        .O(\badr[15]_INST_0_i_317_n_0 ));
  LUT6 #(
    .INIT(64'hF7F7FFF7F7F7FFFF)) 
    \badr[15]_INST_0_i_318 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [15]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [14]),
        .I5(\rgf/sreg/sr [7]),
        .O(\badr[15]_INST_0_i_318_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_319 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [4]),
        .O(\badr[15]_INST_0_i_319_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_320 
       (.I0(\ctl1/stat [1]),
        .I1(\fch/ir1 [1]),
        .O(\badr[15]_INST_0_i_320_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_321 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_321_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF80A0F0FFDFFF)) 
    \badr[15]_INST_0_i_322 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_322_n_0 ));
  LUT6 #(
    .INIT(64'h8080800000008000)) 
    \badr[15]_INST_0_i_323 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_323_n_0 ));
  LUT5 #(
    .INIT(32'hFFFC0FFD)) 
    \badr[15]_INST_0_i_324 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_324_n_0 ));
  LUT5 #(
    .INIT(32'h0000AA8A)) 
    \badr[15]_INST_0_i_325 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_325_n_0 ));
  LUT6 #(
    .INIT(64'hFDF7FFFFFE7EFFFF)) 
    \badr[15]_INST_0_i_326 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [0]),
        .I5(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_326_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_327 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_327_n_0 ));
  LUT4 #(
    .INIT(16'hD0DF)) 
    \badr[15]_INST_0_i_328 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .O(\badr[15]_INST_0_i_328_n_0 ));
  LUT6 #(
    .INIT(64'hFF04FFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_329 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [10]),
        .O(\badr[15]_INST_0_i_329_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_35 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .O(\rgf/a0bus_sel_cr [5]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[15]_INST_0_i_36 
       (.CI(\badr[11]_INST_0_i_29_n_0 ),
        .CO({\badr[15]_INST_0_i_36_n_1 ,\badr[15]_INST_0_i_36_n_2 ,\badr[15]_INST_0_i_36_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rgf/sptr/sp [14:12]}),
        .O(\rgf/sptr/data3 [15:12]),
        .S({\badr[15]_INST_0_i_110_n_0 ,\badr[15]_INST_0_i_111_n_0 ,\badr[15]_INST_0_i_112_n_0 ,\badr[15]_INST_0_i_113_n_0 }));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_37 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .O(\rgf/a0bus_sel_cr [2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_38 
       (.I0(\badr[15]_INST_0_i_28_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .O(\rgf/a0bus_sel_cr [1]));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[15]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_52_n_0 ),
        .I1(ctl_sela1_rn),
        .O(\badr[15]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h4544454545444544)) 
    \badr[15]_INST_0_i_40 
       (.I0(\ctl1/stat [2]),
        .I1(\badr[15]_INST_0_i_114_n_0 ),
        .I2(\badr[15]_INST_0_i_115_n_0 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\badr[15]_INST_0_i_117_n_0 ),
        .I5(\badr[15]_INST_0_i_118_n_0 ),
        .O(\badr[15]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAFFAE)) 
    \badr[15]_INST_0_i_41 
       (.I0(ctl_sela1),
        .I1(\badr[15]_INST_0_i_120_n_0 ),
        .I2(\badr[15]_INST_0_i_121_n_0 ),
        .I3(\badr[15]_INST_0_i_122_n_0 ),
        .I4(\badr[15]_INST_0_i_123_n_0 ),
        .I5(\ctl1/stat [2]),
        .O(\badr[15]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_42 
       (.I0(\badr[15]_INST_0_i_52_n_0 ),
        .I1(ctl_sela1_rn),
        .O(\badr[15]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFABAAAA)) 
    \badr[15]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_140_n_0 ),
        .I1(\badr[15]_INST_0_i_141_n_0 ),
        .I2(\badr[15]_INST_0_i_142_n_0 ),
        .I3(\badr[15]_INST_0_i_143_n_0 ),
        .I4(\badr[15]_INST_0_i_144_n_0 ),
        .I5(\ctl1/stat [2]),
        .O(ctl_sela1_rn));
  LUT6 #(
    .INIT(64'h4544454445444545)) 
    \badr[15]_INST_0_i_52 
       (.I0(\ctl1/stat [2]),
        .I1(\badr[15]_INST_0_i_145_n_0 ),
        .I2(\badr[15]_INST_0_i_115_n_0 ),
        .I3(\badr[15]_INST_0_i_146_n_0 ),
        .I4(\badr[15]_INST_0_i_147_n_0 ),
        .I5(\badr[15]_INST_0_i_148_n_0 ),
        .O(\badr[15]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_59 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(\rgf/a1bus_sel_cr [5]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[15]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/sreg/sr [15]),
        .O(\badr[15]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_60 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(\rgf/a1bus_sel_cr [2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_61 
       (.I0(\badr[15]_INST_0_i_52_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .O(\rgf/a1bus_sel_cr [1]));
  LUT6 #(
    .INIT(64'h4000400040005050)) 
    \badr[15]_INST_0_i_62 
       (.I0(\ctl0/stat [2]),
        .I1(\badr[15]_INST_0_i_165_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\fadr[15]_INST_0_i_15_n_0 ),
        .I5(\fadr[15]_INST_0_i_14_n_0 ),
        .O(\badr[15]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF7577)) 
    \badr[15]_INST_0_i_63 
       (.I0(\stat[2]_i_10_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\badr[15]_INST_0_i_166_n_0 ),
        .I3(\fch/ir0 [2]),
        .I4(\badr[15]_INST_0_i_167_n_0 ),
        .O(\badr[15]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEE0EEE0)) 
    \badr[15]_INST_0_i_64 
       (.I0(\badr[15]_INST_0_i_168_n_0 ),
        .I1(\badr[15]_INST_0_i_169_n_0 ),
        .I2(\badr[15]_INST_0_i_170_n_0 ),
        .I3(\badr[15]_INST_0_i_171_n_0 ),
        .I4(\stat[0]_i_29__0_n_0 ),
        .I5(\badr[15]_INST_0_i_172_n_0 ),
        .O(\badr[15]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hC400FFFFC400C000)) 
    \badr[15]_INST_0_i_65 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [15]),
        .I2(\bcmd[2]_INST_0_i_7_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [11]),
        .I5(\badr[15]_INST_0_i_173_n_0 ),
        .O(\badr[15]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \badr[15]_INST_0_i_66 
       (.I0(\stat[2]_i_6_n_0 ),
        .I1(\badr[15]_INST_0_i_174_n_0 ),
        .I2(\badr[15]_INST_0_i_175_n_0 ),
        .I3(\badr[15]_INST_0_i_176_n_0 ),
        .I4(\badr[15]_INST_0_i_177_n_0 ),
        .I5(\badr[15]_INST_0_i_178_n_0 ),
        .O(ctl_sela0));
  LUT6 #(
    .INIT(64'h555555557F7F7F77)) 
    \badr[15]_INST_0_i_67 
       (.I0(\ccmd[0]_INST_0_i_15_n_0 ),
        .I1(\badr[15]_INST_0_i_179_n_0 ),
        .I2(\badr[15]_INST_0_i_180_n_0 ),
        .I3(\badr[15]_INST_0_i_181_n_0 ),
        .I4(\badr[15]_INST_0_i_182_n_0 ),
        .I5(\fch/ir0 [13]),
        .O(\badr[15]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFEA0000)) 
    \badr[15]_INST_0_i_68 
       (.I0(\bdatw[8]_INST_0_i_41_n_0 ),
        .I1(\ctl0/stat [0]),
        .I2(\bdatw[8]_INST_0_i_43_n_0 ),
        .I3(\badr[15]_INST_0_i_183_n_0 ),
        .I4(\fch/ir0 [13]),
        .I5(\badr[15]_INST_0_i_184_n_0 ),
        .O(\badr[15]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \badr[15]_INST_0_i_69 
       (.I0(\fch/ir0 [12]),
        .I1(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I2(\ccmd[1]_INST_0_i_21_n_0 ),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [13]),
        .I5(\badr[15]_INST_0_i_185_n_0 ),
        .O(\badr[15]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h88888888A8AAA8A8)) 
    \badr[15]_INST_0_i_70 
       (.I0(\badr[15]_INST_0_i_186_n_0 ),
        .I1(\badr[15]_INST_0_i_187_n_0 ),
        .I2(\badr[15]_INST_0_i_188_n_0 ),
        .I3(\badr[15]_INST_0_i_189_n_0 ),
        .I4(\fch/ir0 [14]),
        .I5(\badr[15]_INST_0_i_190_n_0 ),
        .O(\badr[15]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hEABFBFEA)) 
    \badr[15]_INST_0_i_87 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [12]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir0 [11]),
        .I4(\rgf/sreg/sr [5]),
        .O(\badr[15]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF1)) 
    \badr[15]_INST_0_i_88 
       (.I0(\fch/ir0 [11]),
        .I1(\badr[15]_INST_0_i_192_n_0 ),
        .I2(\badr[15]_INST_0_i_193_n_0 ),
        .I3(\badr[15]_INST_0_i_194_n_0 ),
        .I4(\badr[15]_INST_0_i_195_n_0 ),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\badr[15]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0404FF04)) 
    \badr[15]_INST_0_i_89 
       (.I0(\badr[15]_INST_0_i_196_n_0 ),
        .I1(\stat[1]_i_18_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\badr[15]_INST_0_i_197_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .O(\badr[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [15]),
        .I5(\rgf/ivec/iv [15]),
        .O(\badr[15]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEE00E0)) 
    \badr[15]_INST_0_i_90 
       (.I0(\badr[15]_INST_0_i_198_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(\fch/ir0 [0]),
        .I3(\badr[15]_INST_0_i_199_n_0 ),
        .I4(\ccmd[2]_INST_0_i_2_n_0 ),
        .I5(\ctl0/stat [2]),
        .O(\badr[15]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F002F222F2F)) 
    \badr[15]_INST_0_i_91 
       (.I0(\rgf_selc0_rn_wb[0]_i_5_n_0 ),
        .I1(\fadr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_200_n_0 ),
        .I3(\badr[15]_INST_0_i_201_n_0 ),
        .I4(\badr[15]_INST_0_i_202_n_0 ),
        .I5(\fadr[15]_INST_0_i_15_n_0 ),
        .O(\badr[15]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h444F444444444444)) 
    \badr[15]_INST_0_i_92 
       (.I0(\badr[15]_INST_0_i_197_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [11]),
        .I4(\bcmd[0]_INST_0_i_25_n_0 ),
        .I5(\badr[15]_INST_0_i_203_n_0 ),
        .O(\badr[15]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF8)) 
    \badr[15]_INST_0_i_93 
       (.I0(\badr[15]_INST_0_i_204_n_0 ),
        .I1(\badr[15]_INST_0_i_205_n_0 ),
        .I2(\badr[15]_INST_0_i_206_n_0 ),
        .I3(\stat[0]_i_7__1_n_0 ),
        .I4(\badr[15]_INST_0_i_207_n_0 ),
        .I5(\badr[15]_INST_0_i_208_n_0 ),
        .O(\badr[15]_INST_0_i_93_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[1]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[1]),
        .I3(a1bus_0[1]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[1]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[1]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [1]),
        .O(\badr[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [1]),
        .I5(\rgf/ivec/iv [1]),
        .O(\badr[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [1]),
        .O(\badr[1]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [1]),
        .O(\badr[1]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\badr[1]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\badr[1]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [1]),
        .O(\badr[1]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [1]),
        .O(\badr[1]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\badr[1]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\badr[1]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[1]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [1]),
        .O(\badr[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [1]),
        .I5(\rgf/ivec/iv [1]),
        .O(\badr[1]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[2]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[2]),
        .I3(a1bus_0[2]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[2]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[2]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [2]),
        .O(\badr[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [2]),
        .I5(\rgf/ivec/iv [2]),
        .O(\badr[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [2]),
        .O(\badr[2]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [2]),
        .O(\badr[2]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\badr[2]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [2]),
        .O(\badr[2]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [2]),
        .O(\badr[2]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [2]),
        .O(\badr[2]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\badr[2]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [2]),
        .O(\badr[2]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[2]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [2]),
        .O(\badr[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [2]),
        .I5(\rgf/ivec/iv [2]),
        .O(\badr[2]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[3]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[3]),
        .I3(a1bus_0[3]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[3]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[3]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [3]),
        .O(\badr[3]_INST_0_i_12_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[3]_INST_0_i_29 
       (.CI(\<const0> ),
        .CO({\badr[3]_INST_0_i_29_n_0 ,\badr[3]_INST_0_i_29_n_1 ,\badr[3]_INST_0_i_29_n_2 ,\badr[3]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf/sptr/sp [3:1],\<const0> }),
        .O({\rgf/sptr/data3 [3:1],\NLW_badr[3]_INST_0_i_29_O_UNCONNECTED [0]}),
        .S({\badr[3]_INST_0_i_48_n_0 ,\badr[3]_INST_0_i_49_n_0 ,\badr[3]_INST_0_i_50_n_0 ,\rgf/sptr/sp [0]}));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [3]),
        .I5(\rgf/ivec/iv [3]),
        .O(\badr[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [3]),
        .O(\badr[3]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [3]),
        .O(\badr[3]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\badr[3]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\badr[3]_INST_0_i_47_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_48 
       (.I0(\rgf/sptr/sp [3]),
        .O(\badr[3]_INST_0_i_48_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_49 
       (.I0(\rgf/sptr/sp [2]),
        .O(\badr[3]_INST_0_i_49_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[3]_INST_0_i_50 
       (.I0(\rgf/sptr/sp [1]),
        .O(\badr[3]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [3]),
        .O(\badr[3]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [3]),
        .O(\badr[3]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\badr[3]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_54 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\badr[3]_INST_0_i_54_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[3]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [3]),
        .O(\badr[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [3]),
        .I5(\rgf/ivec/iv [3]),
        .O(\badr[3]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[4]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[4]),
        .I3(a1bus_0[4]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[4]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[4]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [4]),
        .O(\badr[4]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [4]),
        .I5(\rgf/ivec/iv [4]),
        .O(\badr[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [4]),
        .O(\badr[4]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [4]),
        .O(\badr[4]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\badr[4]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [4]),
        .O(\badr[4]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [4]),
        .O(\badr[4]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [4]),
        .O(\badr[4]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\badr[4]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [4]),
        .O(\badr[4]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[4]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [4]),
        .O(\badr[4]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [4]),
        .I5(\rgf/ivec/iv [4]),
        .O(\badr[4]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[5]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[5]),
        .I3(a1bus_0[5]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[5]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[5]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [5]),
        .O(\badr[5]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [5]),
        .I5(\rgf/ivec/iv [5]),
        .O(\badr[5]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [5]),
        .O(\badr[5]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [5]),
        .O(\badr[5]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\badr[5]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [5]),
        .O(\badr[5]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [5]),
        .O(\badr[5]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [5]),
        .O(\badr[5]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\badr[5]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [5]),
        .O(\badr[5]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[5]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [5]),
        .O(\badr[5]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [5]),
        .I5(\rgf/ivec/iv [5]),
        .O(\badr[5]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[6]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[6]),
        .I3(a1bus_0[6]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[6]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[6]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\badr[6]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [6]),
        .I5(\rgf/ivec/iv [6]),
        .O(\badr[6]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [6]),
        .O(\badr[6]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [6]),
        .O(\badr[6]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [6]),
        .O(\badr[6]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [6]),
        .O(\badr[6]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [6]),
        .O(\badr[6]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [6]),
        .O(\badr[6]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [6]),
        .O(\badr[6]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [6]),
        .O(\badr[6]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[6]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\badr[6]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [6]),
        .I5(\rgf/ivec/iv [6]),
        .O(\badr[6]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[7]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[7]),
        .I3(a1bus_0[7]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[7]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[7]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [7]),
        .O(\badr[7]_INST_0_i_12_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[7]_INST_0_i_29 
       (.CI(\badr[3]_INST_0_i_29_n_0 ),
        .CO({\badr[7]_INST_0_i_29_n_0 ,\badr[7]_INST_0_i_29_n_1 ,\badr[7]_INST_0_i_29_n_2 ,\badr[7]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [7:4]),
        .O(\rgf/sptr/data3 [7:4]),
        .S({\badr[7]_INST_0_i_48_n_0 ,\badr[7]_INST_0_i_49_n_0 ,\badr[7]_INST_0_i_50_n_0 ,\badr[7]_INST_0_i_51_n_0 }));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [7]),
        .I5(\rgf/ivec/iv [7]),
        .O(\badr[7]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [7]),
        .O(\badr[7]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [7]),
        .O(\badr[7]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [7]),
        .O(\badr[7]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [7]),
        .O(\badr[7]_INST_0_i_47_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_48 
       (.I0(\rgf/sptr/sp [7]),
        .O(\badr[7]_INST_0_i_48_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_49 
       (.I0(\rgf/sptr/sp [6]),
        .O(\badr[7]_INST_0_i_49_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_50 
       (.I0(\rgf/sptr/sp [5]),
        .O(\badr[7]_INST_0_i_50_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \badr[7]_INST_0_i_51 
       (.I0(\rgf/sptr/sp [4]),
        .O(\badr[7]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [7]),
        .O(\badr[7]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [7]),
        .O(\badr[7]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_54 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [7]),
        .O(\badr[7]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_55 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [7]),
        .O(\badr[7]_INST_0_i_55_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[7]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [7]),
        .O(\badr[7]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [7]),
        .I5(\rgf/ivec/iv [7]),
        .O(\badr[7]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[8]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[8]),
        .I3(a1bus_0[8]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[8]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[8]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\badr[8]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [8]),
        .I5(\rgf/ivec/iv [8]),
        .O(\badr[8]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [8]),
        .O(\badr[8]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [8]),
        .O(\badr[8]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [8]),
        .O(\badr[8]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [8]),
        .O(\badr[8]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [8]),
        .O(\badr[8]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [8]),
        .O(\badr[8]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [8]),
        .O(\badr[8]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [8]),
        .O(\badr[8]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[8]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\badr[8]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [8]),
        .I5(\rgf/ivec/iv [8]),
        .O(\badr[8]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hE0E0EE00)) 
    \badr[9]_INST_0 
       (.I0(bcmd[0]),
        .I1(bcmd[1]),
        .I2(a0bus_0[9]),
        .I3(a1bus_0[9]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(badr[9]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[9]_INST_0_i_12 
       (.I0(\badr[15]_INST_0_i_40_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/sreg/sr [9]),
        .O(\badr[9]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_3 
       (.I0(\badr[15]_INST_0_i_15_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_17_n_0 ),
        .I3(\badr[15]_INST_0_i_18_n_0 ),
        .I4(\rgf/treg/tr [9]),
        .I5(\rgf/ivec/iv [9]),
        .O(\badr[9]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [9]),
        .O(\badr[9]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [9]),
        .O(\badr[9]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [9]),
        .O(\badr[9]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [9]),
        .O(\badr[9]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr21 [9]),
        .O(\badr[9]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr22 [9]),
        .O(\badr[9]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr25 [9]),
        .O(\badr[9]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [9]),
        .O(\badr[9]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[9]_INST_0_i_6 
       (.I0(ctl_sela0_rn[2]),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(\badr[15]_INST_0_i_17_n_0 ),
        .I4(\rgf/sreg/sr [9]),
        .O(\badr[9]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_9 
       (.I0(\badr[15]_INST_0_i_39_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_41_n_0 ),
        .I3(\badr[15]_INST_0_i_42_n_0 ),
        .I4(\rgf/treg/tr [9]),
        .I5(\rgf/ivec/iv [9]),
        .O(\badr[9]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[0]_INST_0 
       (.I0(\rgf/treg/tr [0]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[10]_INST_0 
       (.I0(\rgf/treg/tr [10]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[11]_INST_0 
       (.I0(\rgf/treg/tr [11]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[11]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[12]_INST_0 
       (.I0(\rgf/treg/tr [12]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[12]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[13]_INST_0 
       (.I0(\rgf/treg/tr [13]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[14]_INST_0 
       (.I0(\rgf/treg/tr [14]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[14]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[15]_INST_0 
       (.I0(\rgf/treg/tr [15]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[15]));
  MUXF7 \badrx[15]_INST_0_i_1 
       (.I0(\badrx[15]_INST_0_i_2_n_0 ),
        .I1(\badrx[15]_INST_0_i_3_n_0 ),
        .O(\badrx[15]_INST_0_i_1_n_0 ),
        .S(\bcmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFFFFFFFFFFFFF)) 
    \badrx[15]_INST_0_i_2 
       (.I0(\bcmd[2]_INST_0_i_4_n_0 ),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [9]),
        .O(\badrx[15]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBF)) 
    \badrx[15]_INST_0_i_3 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\badrx[15]_INST_0_i_4_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\ctl0/stat [0]),
        .I5(\badrx[15]_INST_0_i_5_n_0 ),
        .O(\badrx[15]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badrx[15]_INST_0_i_4 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .O(\badrx[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    \badrx[15]_INST_0_i_5 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\ctl0/stat [2]),
        .I4(\ctl0/stat [1]),
        .I5(\fch/ir0 [15]),
        .O(\badrx[15]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[1]_INST_0 
       (.I0(\rgf/treg/tr [1]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[2]_INST_0 
       (.I0(\rgf/treg/tr [2]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[3]_INST_0 
       (.I0(\rgf/treg/tr [3]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[4]_INST_0 
       (.I0(\rgf/treg/tr [4]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[5]_INST_0 
       (.I0(\rgf/treg/tr [5]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[6]_INST_0 
       (.I0(\rgf/treg/tr [6]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[6]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[7]_INST_0 
       (.I0(\rgf/treg/tr [7]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[7]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[8]_INST_0 
       (.I0(\rgf/treg/tr [8]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[8]));
  LUT2 #(
    .INIT(4'h2)) 
    \badrx[9]_INST_0 
       (.I0(\rgf/treg/tr [9]),
        .I1(\badrx[15]_INST_0_i_1_n_0 ),
        .O(badrx[9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn00/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn00/grn1 ),
        .O(\rgf/p_2_in [9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn01/grn1 ),
        .O(\bank02/grn01/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn02/grn1 ),
        .O(\bank02/grn02/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn03/grn1 ),
        .O(\bank02/grn03/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn04/grn1 ),
        .O(\bank02/grn04/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn05/grn1 ),
        .O(\bank02/grn05/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn06/grn1 ),
        .O(\bank02/grn06/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn07/grn1 ),
        .O(\bank02/grn07/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn20/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn20/grn1 ),
        .O(\bank02/grn20/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn21/grn1 ),
        .O(\bank02/grn21/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn22/grn1 ),
        .O(\bank02/grn22/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn23/grn1 ),
        .O(\bank02/grn23/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn24/grn1 ),
        .O(\bank02/grn24/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn25/grn1 ),
        .O(\bank02/grn25/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn26/grn1 ),
        .O(\bank02/grn26/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank02/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn27/grn1 ),
        .O(\bank02/grn27/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn00/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn00/grn1 ),
        .O(\bank13/grn00/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn01/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn01/grn1 ),
        .O(\bank13/grn01/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn02/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn02/grn1 ),
        .O(\bank13/grn02/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn03/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn03/grn1 ),
        .O(\bank13/grn03/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn04/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn04/grn1 ),
        .O(\bank13/grn04/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn05/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn05/grn1 ),
        .O(\bank13/grn05/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn06/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn06/grn1 ),
        .O(\bank13/grn06/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn07/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn07/grn1 ),
        .O(\bank13/grn07/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn20/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn20/grn1 ),
        .O(\bank13/grn20/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn21/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn21/grn1 ),
        .O(\bank13/grn21/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn22/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn22/grn1 ),
        .O(\bank13/grn22/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn23/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn23/grn1 ),
        .O(\bank13/grn23/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn24/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn24/grn1 ),
        .O(\bank13/grn24/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn25/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn25/grn1 ),
        .O(\bank13/grn25/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn26/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn26/grn1 ),
        .O(\bank13/grn26/grn[9]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[10]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[11]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[12]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[13]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[14]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[15]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[7]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[8]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \bank13/grn27/grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn27/grn1 ),
        .O(\bank13/grn27/grn[9]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[0]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(bbus_o[0]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[0]_INST_0_i_1 
       (.I0(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[0]_INST_0_i_4_n_0 ),
        .I3(\rgf/b0bus_b02 [0]),
        .I4(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I5(\rgf/b0bus_out/bbus_o[0]_INST_0_i_7_n_0 ),
        .O(\bbus_o[0]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[0]_INST_0_i_15 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\rgf/sreg/sr [0]),
        .O(\bbus_o[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0FF0FFD2)) 
    \bbus_o[0]_INST_0_i_2 
       (.I0(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I1(\fch/ir0 [1]),
        .I2(\bdatw[15]_INST_0_i_22_n_0 ),
        .I3(\bdatw[15]_INST_0_i_19_n_0 ),
        .I4(\fch/ir0 [0]),
        .I5(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bbus_o[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[0]_INST_0_i_23 
       (.I0(\bdatw[15]_INST_0_i_80_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/bank13/gr20 [0]),
        .O(\bbus_o[0]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[0]_INST_0_i_24 
       (.I0(\bdatw[15]_INST_0_i_81_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [0]),
        .O(\bbus_o[0]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[0]_INST_0_i_3 
       (.I0(\fch/eir [0]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[0]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bbus_o[0]_INST_0_i_8 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [2]),
        .O(\bbus_o[0]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[10]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[10]_INST_0_i_1_n_0 ),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[11]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[11]_INST_0_i_1_n_0 ),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[12]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[12]_INST_0_i_1_n_0 ),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[13]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[13]_INST_0_i_1_n_0 ),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[14]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[14]_INST_0_i_1_n_0 ),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[15]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_1_n_0 ),
        .O(bbus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[1]_INST_0 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(bbus_o[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \bbus_o[1]_INST_0_i_1 
       (.I0(\bbus_o[1]_INST_0_i_2_n_0 ),
        .I1(\rgf/b0bus_out/bbus_o[1]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_b02 [1]),
        .I3(\rgf/b0bus_out/bbus_o[1]_INST_0_i_5_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[1]_INST_0_i_6_n_0 ),
        .I5(\bbus_o[1]_INST_0_i_7_n_0 ),
        .O(\bbus_o[1]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[1]_INST_0_i_14 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\rgf/sreg/sr [1]),
        .O(\bbus_o[1]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[1]_INST_0_i_2 
       (.I0(\fch/eir [1]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[1]_INST_0_i_22 
       (.I0(\bdatw[15]_INST_0_i_80_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/bank13/gr20 [1]),
        .O(\bbus_o[1]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[1]_INST_0_i_23 
       (.I0(\bdatw[15]_INST_0_i_81_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\bbus_o[1]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEABFBFEFEABFB)) 
    \bbus_o[1]_INST_0_i_7 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\fadr[15]_INST_0_i_14_n_0 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [0]),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [1]),
        .O(\bbus_o[1]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[2]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(bbus_o[2]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[2]_INST_0_i_1 
       (.I0(\bbus_o[2]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[2]_INST_0_i_4_n_0 ),
        .I3(\rgf/b0bus_b02 [2]),
        .I4(\rgf/b0bus_out/bbus_o[2]_INST_0_i_6_n_0 ),
        .I5(\rgf/b0bus_out/bbus_o[2]_INST_0_i_7_n_0 ),
        .O(\bbus_o[2]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[2]_INST_0_i_15 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\rgf/sreg/sr [2]),
        .O(\bbus_o[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hABABAEFEFBFBAEFE)) 
    \bbus_o[2]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_8_n_0 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [1]),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [2]),
        .O(\bbus_o[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[2]_INST_0_i_23 
       (.I0(\bdatw[15]_INST_0_i_80_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/bank13/gr20 [2]),
        .O(\bbus_o[2]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[2]_INST_0_i_24 
       (.I0(\bdatw[15]_INST_0_i_81_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [2]),
        .O(\bbus_o[2]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[2]_INST_0_i_3 
       (.I0(\fch/eir [2]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[2]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \bbus_o[2]_INST_0_i_8 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [0]),
        .O(\bbus_o[2]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[3]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(bbus_o[3]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[3]_INST_0_i_1 
       (.I0(\bbus_o[3]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[3]_INST_0_i_4_n_0 ),
        .I3(\rgf/b0bus_b02 [3]),
        .I4(\rgf/b0bus_out/bbus_o[3]_INST_0_i_6_n_0 ),
        .I5(\rgf/b0bus_out/bbus_o[3]_INST_0_i_7_n_0 ),
        .O(\bbus_o[3]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[3]_INST_0_i_15 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\rgf/sreg/sr [3]),
        .O(\bbus_o[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAFFFBAFAFFFFBA)) 
    \bbus_o[3]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\fch/ir0 [2]),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_8_n_0 ),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [3]),
        .O(\bbus_o[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[3]_INST_0_i_23 
       (.I0(\bdatw[15]_INST_0_i_80_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/bank13/gr20 [3]),
        .O(\bbus_o[3]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[3]_INST_0_i_24 
       (.I0(\bdatw[15]_INST_0_i_81_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\bbus_o[3]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[3]_INST_0_i_3 
       (.I0(\fch/eir [3]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[3]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bbus_o[3]_INST_0_i_8 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [2]),
        .O(\bbus_o[3]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[4]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(bbus_o[4]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[4]_INST_0_i_1 
       (.I0(\bbus_o[4]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[4]_INST_0_i_4_n_0 ),
        .I3(\rgf/b0bus_b02 [4]),
        .I4(\rgf/b0bus_out/bbus_o[4]_INST_0_i_6_n_0 ),
        .I5(\rgf/b0bus_out/bbus_o[4]_INST_0_i_7_n_0 ),
        .O(\bbus_o[4]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bbus_o[4]_INST_0_i_15 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_77_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(\rgf/sreg/sr [4]),
        .O(\bbus_o[4]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hABABEEFEFBFBEEFE)) 
    \bbus_o[4]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_8_n_0 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [3]),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [4]),
        .O(\bbus_o[4]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \bbus_o[4]_INST_0_i_21 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[8]_INST_0_i_5_n_0 ),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\rgf/b0bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \bbus_o[4]_INST_0_i_22 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[8]_INST_0_i_5_n_0 ),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\rgf/b0bus_sel_cr [2]));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \bbus_o[4]_INST_0_i_23 
       (.I0(ctl_selb0_rn[1]),
        .I1(\bdatw[15]_INST_0_i_76_n_0 ),
        .I2(ctl_selb0_rn[0]),
        .I3(\bdatw[8]_INST_0_i_5_n_0 ),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\rgf/b0bus_sel_cr [1]));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \bbus_o[4]_INST_0_i_26 
       (.I0(\bdatw[15]_INST_0_i_80_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/bank13/gr20 [4]),
        .O(\bbus_o[4]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \bbus_o[4]_INST_0_i_28 
       (.I0(\bdatw[15]_INST_0_i_81_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [4]),
        .O(\bbus_o[4]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[4]_INST_0_i_3 
       (.I0(\fch/eir [4]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[4]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bbus_o[4]_INST_0_i_8 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [3]),
        .O(\bbus_o[4]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(bbus_o[5]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bbus_o[5]_INST_0_i_1 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[5]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [5]),
        .I4(\rgf/bank02/p_0_in2_in [5]),
        .I5(\rgf/b0bus_out/bbus_o[5]_INST_0_i_7_n_0 ),
        .O(\bbus_o[5]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[5]_INST_0_i_18 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [5]),
        .O(\bbus_o[5]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h5454510104045101)) 
    \bbus_o[5]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_8_n_0 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [4]),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [5]),
        .O(\bbus_o[5]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0_i_3 
       (.I0(\fch/eir [5]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[5]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \bbus_o[5]_INST_0_i_8 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [3]),
        .O(\bbus_o[5]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[6]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[6]_INST_0_i_1_n_0 ),
        .O(bbus_o[6]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bbus_o[6]_INST_0_i_1 
       (.I0(\bbus_o[6]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[6]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[6]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [6]),
        .I4(\rgf/bank02/p_0_in2_in [6]),
        .I5(\rgf/b0bus_out/bbus_o[6]_INST_0_i_7_n_0 ),
        .O(\bbus_o[6]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[6]_INST_0_i_18 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [6]),
        .O(\bbus_o[6]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h5454510104045101)) 
    \bbus_o[6]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bbus_o[6]_INST_0_i_8_n_0 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [5]),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [6]),
        .O(\bbus_o[6]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[6]_INST_0_i_3 
       (.I0(\fch/eir [6]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[6]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \bbus_o[6]_INST_0_i_8 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [3]),
        .O(\bbus_o[6]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[7]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_1_n_0 ),
        .O(bbus_o[7]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[7]_INST_0_i_1 
       (.I0(\bbus_o[7]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [7]),
        .I4(\rgf/bank02/p_0_in2_in [7]),
        .I5(\rgf/b0bus_out/bbus_o[7]_INST_0_i_7_n_0 ),
        .O(\bbus_o[7]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[7]_INST_0_i_18 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [7]),
        .O(\bbus_o[7]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hABABEEFEBBBBEEFE)) 
    \bbus_o[7]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_8_n_0 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [6]),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [7]),
        .O(\bbus_o[7]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[7]_INST_0_i_3 
       (.I0(\fch/eir [7]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bbus_o[7]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \bbus_o[7]_INST_0_i_8 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [2]),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .O(\bbus_o[7]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[8]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[8]_INST_0_i_1_n_0 ),
        .O(bbus_o[8]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[9]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bdatw[9]_INST_0_i_1_n_0 ),
        .O(bbus_o[9]));
  MUXF7 \bcmd[0]_INST_0 
       (.I0(\bcmd[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_2_n_0 ),
        .O(bcmd[0]),
        .S(\bcmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0200020002000203)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\bcmd[0]_INST_0_i_4_n_0 ),
        .I2(\bcmd[0]_INST_0_i_5_n_0 ),
        .I3(\fch/ir1 [12]),
        .I4(\bcmd[0]_INST_0_i_6_n_0 ),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h4000000004400440)) 
    \bcmd[0]_INST_0_i_10 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [6]),
        .O(\bcmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF35FF)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(\bcmd[0]_INST_0_i_18_n_0 ),
        .I1(\bcmd[0]_INST_0_i_19_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\bcmd[0]_INST_0_i_20_n_0 ),
        .I4(\bcmd[0]_INST_0_i_21_n_0 ),
        .I5(\bcmd[0]_INST_0_i_22_n_0 ),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h4545555445455555)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [1]),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7F0FF50)) 
    \bcmd[0]_INST_0_i_13 
       (.I0(\bcmd[0]_INST_0_i_23_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(\bcmd[0]_INST_0_i_24_n_0 ),
        .O(\bcmd[0]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[0]_INST_0_i_14 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [3]),
        .O(\bcmd[0]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_15 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [0]),
        .O(\bcmd[0]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_16 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .O(\bcmd[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h757DFD7DFD7DFD7D)) 
    \bcmd[0]_INST_0_i_17 
       (.I0(\bcmd[1]_INST_0_i_3_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [7]),
        .O(\bcmd[0]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bcmd[0]_INST_0_i_18 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_6_n_0 ),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [5]),
        .O(\bcmd[0]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[0]_INST_0_i_19 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .O(\bcmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF4F)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(\bcmd[0]_INST_0_i_8_n_0 ),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\bcmd[0]_INST_0_i_10_n_0 ),
        .I4(\bcmd[0]_INST_0_i_11_n_0 ),
        .I5(\bcmd[0]_INST_0_i_12_n_0 ),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_20 
       (.I0(\fch/ir0 [15]),
        .I1(\ctl0/stat [1]),
        .I2(\ctl0/stat [2]),
        .O(\bcmd[0]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h02A2A2A2)) 
    \bcmd[0]_INST_0_i_21 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [3]),
        .O(\bcmd[0]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \bcmd[0]_INST_0_i_22 
       (.I0(\fch/ir0 [5]),
        .I1(\bcmd[0]_INST_0_i_25_n_0 ),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\bdatw[10]_INST_0_i_15_n_0 ),
        .I4(\fch/ir0 [4]),
        .I5(\ctl0/stat [0]),
        .O(\bcmd[0]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[0]_INST_0_i_23 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [10]),
        .O(\bcmd[0]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[0]_INST_0_i_24 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .O(\bcmd[0]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[0]_INST_0_i_25 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [3]),
        .O(\bcmd[0]_INST_0_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_26 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [7]),
        .O(\bcmd[0]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF28)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [11]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [6]),
        .I5(\bcmd[0]_INST_0_i_13_n_0 ),
        .O(\bcmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(\fch/ir1 [5]),
        .I1(\bcmd[0]_INST_0_i_14_n_0 ),
        .I2(\fch/ir1 [4]),
        .I3(\ctl1/stat [0]),
        .I4(\bcmd[0]_INST_0_i_15_n_0 ),
        .I5(\bcmd[0]_INST_0_i_16_n_0 ),
        .O(\bcmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF13121313)) 
    \bcmd[0]_INST_0_i_5 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .I5(\bcmd[0]_INST_0_i_17_n_0 ),
        .O(\bcmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [2]),
        .O(\bcmd[0]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .O(\bcmd[0]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [6]),
        .O(\bcmd[0]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[0]_INST_0_i_9 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\ctl0/stat [0]),
        .O(\bcmd[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0400040004FF0400)) 
    \bcmd[1]_INST_0 
       (.I0(\ctl0/stat [2]),
        .I1(\bcmd[1]_INST_0_i_1_n_0 ),
        .I2(\bcmd[1]_INST_0_i_2_n_0 ),
        .I3(\bcmd[2]_INST_0_i_1_n_0 ),
        .I4(\bcmd[1]_INST_0_i_3_n_0 ),
        .I5(\bcmd[1]_INST_0_i_4_n_0 ),
        .O(bcmd[1]));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [15]),
        .O(\bcmd[1]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00001819)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [12]),
        .I2(\ctl1/stat [0]),
        .I3(\pc0[15]_i_3_n_0 ),
        .I4(\bcmd[1]_INST_0_i_16_n_0 ),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(crdy),
        .O(\bcmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000200F00000000)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .I4(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEFFFFFE)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\bcmd[1]_INST_0_i_17_n_0 ),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFFFFFFFF7E)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [9]),
        .O(\bcmd[1]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [3]),
        .O(\bcmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEFFEFF)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(\bcmd[1]_INST_0_i_18_n_0 ),
        .I1(\bcmd[0]_INST_0_i_7_n_0 ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [3]),
        .I5(\bcmd[1]_INST_0_i_19_n_0 ),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h67FFFFFF67FFFF67)) 
    \bcmd[1]_INST_0_i_17 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [2]),
        .O(\bcmd[1]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0FFFFFFE)) 
    \bcmd[1]_INST_0_i_18 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [8]),
        .O(\bcmd[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFFFFFFFF7E)) 
    \bcmd[1]_INST_0_i_19 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [11]),
        .O(\bcmd[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF9FFF)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [9]),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\fch/ir0 [6]),
        .I4(\bcmd[1]_INST_0_i_6_n_0 ),
        .I5(\bcmd[1]_INST_0_i_7_n_0 ),
        .O(\bcmd[1]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(\ctl1/stat [1]),
        .I1(\fch/ir1 [15]),
        .I2(\ctl1/stat [2]),
        .O(\bcmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF9FFF)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(\fch/ir1 [9]),
        .I1(\ctl1/stat [0]),
        .I2(\bcmd[1]_INST_0_i_8_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\bcmd[1]_INST_0_i_9_n_0 ),
        .I5(\bcmd[1]_INST_0_i_10_n_0 ),
        .O(\bcmd[1]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h3033233333333333)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\bcmd[1]_INST_0_i_12_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [8]),
        .O(\bcmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001819)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [12]),
        .I2(\ctl0/stat [0]),
        .I3(\pc0[15]_i_3_n_0 ),
        .I4(\bcmd[1]_INST_0_i_13_n_0 ),
        .I5(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [12]),
        .O(\bcmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h7FF50FFF0FFFFFFF)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(\fch/ir1 [7]),
        .I1(\bcmd[1]_INST_0_i_15_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [10]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  MUXF7 \bcmd[2]_INST_0 
       (.I0(\bcmd[2]_INST_0_i_2_n_0 ),
        .I1(\bcmd[2]_INST_0_i_3_n_0 ),
        .O(bcmd[2]),
        .S(\bcmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF2F33333333)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(\mem/bctl/ctl/p_0_in [5]),
        .I1(\mem/bctl/ctl/p_0_in [4]),
        .I2(fch_memacc1),
        .I3(\fch/ir0_id ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(\mem/bctl/fch_term_fl ),
        .O(\bcmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(\ctl1/stat [0]),
        .I1(\bcmd[2]_INST_0_i_4_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\bcmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000020002000000)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\ctl0/stat [0]),
        .I2(\ctl0/stat [1]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [11]),
        .O(\bcmd[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \bcmd[2]_INST_0_i_4 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\ctl1/stat [1]),
        .I5(\ctl1/stat [2]),
        .O(\bcmd[2]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[2]_INST_0_i_5 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [10]),
        .O(\bcmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \bcmd[2]_INST_0_i_6 
       (.I0(\bcmd[2]_INST_0_i_7_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [14]),
        .I3(\ctl0/stat [2]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [7]),
        .O(\bcmd[2]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[2]_INST_0_i_7 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [12]),
        .O(\bcmd[2]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[0]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[8]_INST_0_i_3_n_0 ),
        .O(bdatw[0]));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[10]_INST_0 
       (.I0(\bdatw[10]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[10]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[10]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[10]));
  LUT5 #(
    .INIT(32'h00000051)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(\bdatw[10]_INST_0_i_4_n_0 ),
        .I1(\fch/eir [10]),
        .I2(\bdatw[10]_INST_0_i_5_n_0 ),
        .I3(\rgf/b0bus_out/bdatw[10]_INST_0_i_6_n_0 ),
        .I4(\rgf/b0bus_out/bdatw[10]_INST_0_i_7_n_0 ),
        .O(\bdatw[10]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[10]_INST_0_i_14 
       (.I0(\bdatw[10]_INST_0_i_33_n_0 ),
        .I1(\bdatw[10]_INST_0_i_34_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[10]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_37_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[10]_INST_0_i_38_n_0 ),
        .O(\bdatw[10]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[10]_INST_0_i_15 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [2]),
        .O(\bdatw[10]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(\bdatw[10]_INST_0_i_8_n_0 ),
        .I1(\bdatw[10]_INST_0_i_9_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[10]_INST_0_i_10_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_11_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_12_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[10]_INST_0_i_13_n_0 ),
        .O(\bdatw[10]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bdatw[10]_INST_0_i_21 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(ctl_selb0_rn[0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_77_n_0 ),
        .O(\rgf/b0bus_sel_cr [0]));
  LUT5 #(
    .INIT(32'h00000040)) 
    \bdatw[10]_INST_0_i_22 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [0]),
        .I4(\bdatw[15]_INST_0_i_40_n_0 ),
        .O(\bdatw[10]_INST_0_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\bdatw[10]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[10]_INST_0_i_32 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [10]),
        .O(\bdatw[10]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h221DEE1DFFFFFFFF)) 
    \bdatw[10]_INST_0_i_33 
       (.I0(\bdatw[10]_INST_0_i_53_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(\fch/ir1 [2]),
        .I3(ctl_selb1_0),
        .I4(\fch/ir1 [1]),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bdatw[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[10]_INST_0_i_34 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [2]),
        .O(\bdatw[10]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h1044101110111011)) 
    \bdatw[10]_INST_0_i_4 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bdatw[15]_INST_0_i_22_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\bdatw[15]_INST_0_i_19_n_0 ),
        .I4(\bdatw[15]_INST_0_i_20_n_0 ),
        .I5(\bdatw[10]_INST_0_i_15_n_0 ),
        .O(\bdatw[10]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \bdatw[10]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_22_n_0 ),
        .I1(\bdatw[15]_INST_0_i_19_n_0 ),
        .I2(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bdatw[10]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \bdatw[10]_INST_0_i_53 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [2]),
        .O(\bdatw[10]_INST_0_i_53_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[10]_INST_0_i_67 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\rgf/sreg/sr [2]),
        .O(\bdatw[10]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_72 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr03 [2]),
        .O(\bdatw[10]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_73 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr04 [2]),
        .O(\bdatw[10]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[10]_INST_0_i_74 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr07 [2]),
        .O(\bdatw[10]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_75 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr06 [2]),
        .O(\bdatw[10]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_76 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr23 [2]),
        .O(\bdatw[10]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_77 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr24 [2]),
        .O(\bdatw[10]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[10]_INST_0_i_78 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr27 [2]),
        .O(\bdatw[10]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[10]_INST_0_i_79 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [2]),
        .O(\bdatw[10]_INST_0_i_79_n_0 ));
  LUT5 #(
    .INIT(32'hD7D7F7D7)) 
    \bdatw[10]_INST_0_i_8 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[10]_INST_0_i_22_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(\fch/ir1 [9]),
        .O(\bdatw[10]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[10]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [10]),
        .O(\bdatw[10]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[11]_INST_0 
       (.I0(\bdatw[11]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[11]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[11]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[11]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(\bdatw[11]_INST_0_i_4_n_0 ),
        .I1(\bdatw[11]_INST_0_i_5_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[11]_INST_0_i_6_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [11]),
        .I4(\rgf/bank02/p_0_in2_in [11]),
        .I5(\rgf/b0bus_out/bdatw[11]_INST_0_i_9_n_0 ),
        .O(\bdatw[11]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8AAA200002222000)) 
    \bdatw[11]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(\bdatw[11]_INST_0_i_27_n_0 ),
        .I3(\bdatw[11]_INST_0_i_28_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\fch/ir1 [10]),
        .O(\bdatw[11]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[11]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [11]),
        .O(\bdatw[11]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[11]_INST_0_i_16 
       (.I0(\bdatw[11]_INST_0_i_39_n_0 ),
        .I1(\bdatw[11]_INST_0_i_40_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[11]_INST_0_i_41_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_42_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[11]_INST_0_i_44_n_0 ),
        .O(\bdatw[11]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(\bdatw[11]_INST_0_i_10_n_0 ),
        .I1(\bdatw[11]_INST_0_i_11_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[11]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_14_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[11]_INST_0_i_15_n_0 ),
        .O(\bdatw[11]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_26 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [11]),
        .O(\bdatw[11]_INST_0_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_27 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [1]),
        .O(\bdatw[11]_INST_0_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_28 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [2]),
        .O(\bdatw[11]_INST_0_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[11]_INST_0_i_3 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\bdatw[11]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[11]_INST_0_i_38 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [11]),
        .O(\bdatw[11]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0F70AF70FFFFFFFF)) 
    \bdatw[11]_INST_0_i_39 
       (.I0(\bdatw[15]_INST_0_i_40_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\bdatw[11]_INST_0_i_57_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\fch/ir1 [2]),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bdatw[11]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h1011104410111011)) 
    \bdatw[11]_INST_0_i_4 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bdatw[15]_INST_0_i_22_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\bdatw[15]_INST_0_i_19_n_0 ),
        .I4(\fadr[15]_INST_0_i_10_n_0 ),
        .I5(\bdatw[15]_INST_0_i_20_n_0 ),
        .O(\bdatw[11]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[11]_INST_0_i_40 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [3]),
        .O(\bdatw[11]_INST_0_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_5 
       (.I0(\fch/eir [11]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bdatw[11]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \bdatw[11]_INST_0_i_57 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [2]),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .O(\bdatw[11]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[11]_INST_0_i_71 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\rgf/sreg/sr [3]),
        .O(\bdatw[11]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_72 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr03 [3]),
        .O(\bdatw[11]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_73 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr04 [3]),
        .O(\bdatw[11]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[11]_INST_0_i_74 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr07 [3]),
        .O(\bdatw[11]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_75 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr06 [3]),
        .O(\bdatw[11]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_76 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr23 [3]),
        .O(\bdatw[11]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_77 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr24 [3]),
        .O(\bdatw[11]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[11]_INST_0_i_78 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr27 [3]),
        .O(\bdatw[11]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[11]_INST_0_i_79 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\bdatw[11]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[12]_INST_0 
       (.I0(\bdatw[12]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[12]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[12]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[12]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(\bdatw[12]_INST_0_i_4_n_0 ),
        .I1(\bdatw[12]_INST_0_i_5_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[12]_INST_0_i_6_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [12]),
        .I4(\rgf/bank02/p_0_in2_in [12]),
        .I5(\rgf/b0bus_out/bdatw[12]_INST_0_i_9_n_0 ),
        .O(\bdatw[12]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDF5575FFDF)) 
    \bdatw[12]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[14]_INST_0_i_29_n_0 ),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [1]),
        .I4(ctl_selb1_0),
        .I5(\bdatw[14]_INST_0_i_30_n_0 ),
        .O(\bdatw[12]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[12]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [12]),
        .O(\bdatw[12]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[12]_INST_0_i_16 
       (.I0(\bdatw[12]_INST_0_i_38_n_0 ),
        .I1(\bdatw[12]_INST_0_i_39_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[12]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_42_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[12]_INST_0_i_43_n_0 ),
        .O(\bdatw[12]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \bdatw[12]_INST_0_i_17 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [3]),
        .O(\bdatw[12]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(\bdatw[12]_INST_0_i_10_n_0 ),
        .I1(\bdatw[12]_INST_0_i_11_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[12]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[12]_INST_0_i_15_n_0 ),
        .O(\bdatw[12]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_27 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [12]),
        .O(\bdatw[12]_INST_0_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\bdatw[12]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[12]_INST_0_i_37 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [12]),
        .O(\bdatw[12]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h5027FA27FFFFFFFF)) 
    \bdatw[12]_INST_0_i_38 
       (.I0(\bdatw[15]_INST_0_i_40_n_0 ),
        .I1(\fch/ir1 [4]),
        .I2(\bdatw[12]_INST_0_i_56_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\fch/ir1 [3]),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bdatw[12]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[12]_INST_0_i_39 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [4]),
        .O(\bdatw[12]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h0000308B)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(\fch/ir0 [10]),
        .I1(\bdatw[15]_INST_0_i_19_n_0 ),
        .I2(\bdatw[12]_INST_0_i_17_n_0 ),
        .I3(\bdatw[15]_INST_0_i_22_n_0 ),
        .I4(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bdatw[12]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[12]_INST_0_i_5 
       (.I0(\fch/eir [12]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bdatw[12]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[12]_INST_0_i_56 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [2]),
        .O(\bdatw[12]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[12]_INST_0_i_70 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\rgf/sreg/sr [4]),
        .O(\bdatw[12]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_71 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr03 [4]),
        .O(\bdatw[12]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_72 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr04 [4]),
        .O(\bdatw[12]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[12]_INST_0_i_73 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr07 [4]),
        .O(\bdatw[12]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_74 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr06 [4]),
        .O(\bdatw[12]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_75 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr23 [4]),
        .O(\bdatw[12]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_76 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr24 [4]),
        .O(\bdatw[12]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[12]_INST_0_i_77 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr27 [4]),
        .O(\bdatw[12]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_78 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [4]),
        .O(\bdatw[12]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFEFEFFFEFF)) 
    \bdatw[12]_INST_0_i_79 
       (.I0(\bdatw[12]_INST_0_i_80_n_0 ),
        .I1(\bdatw[12]_INST_0_i_81_n_0 ),
        .I2(\bdatw[12]_INST_0_i_82_n_0 ),
        .I3(\ctl1/stat [0]),
        .I4(\bdatw[12]_INST_0_i_83_n_0 ),
        .I5(\stat[2]_i_5__0_n_0 ),
        .O(\bdatw[12]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h1151115511111155)) 
    \bdatw[12]_INST_0_i_80 
       (.I0(\bcmd[2]_INST_0_i_4_n_0 ),
        .I1(\bcmd[1]_INST_0_i_3_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(\bdatw[15]_INST_0_i_208_n_0 ),
        .O(\bdatw[12]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    \bdatw[12]_INST_0_i_81 
       (.I0(\bdatw[12]_INST_0_i_84_n_0 ),
        .I1(\bdatw[12]_INST_0_i_85_n_0 ),
        .I2(\bdatw[12]_INST_0_i_86_n_0 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\bdatw[15]_INST_0_i_219_n_0 ),
        .I5(\bdatw[12]_INST_0_i_87_n_0 ),
        .O(\bdatw[12]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFBFBFFFBAAAAAAAA)) 
    \bdatw[12]_INST_0_i_82 
       (.I0(\fch/ir1 [15]),
        .I1(\bdatw[12]_INST_0_i_88_n_0 ),
        .I2(\bdatw[15]_INST_0_i_215_n_0 ),
        .I3(\stat[1]_i_5__0_n_0 ),
        .I4(\bdatw[12]_INST_0_i_89_n_0 ),
        .I5(\ctl1/stat [0]),
        .O(\bdatw[12]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h0000000DDDDD000D)) 
    \bdatw[12]_INST_0_i_83 
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(\bdatw[12]_INST_0_i_90_n_0 ),
        .I2(\bdatw[12]_INST_0_i_91_n_0 ),
        .I3(\bdatw[12]_INST_0_i_92_n_0 ),
        .I4(\fch/ir1 [12]),
        .I5(\bdatw[15]_INST_0_i_210_n_0 ),
        .O(\bdatw[12]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAAAAAEFAAEF)) 
    \bdatw[12]_INST_0_i_84 
       (.I0(\ctl1/stat [0]),
        .I1(\bdatw[15]_INST_0_i_274_n_0 ),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [11]),
        .I4(\bdatw[15]_INST_0_i_275_n_0 ),
        .I5(\bdatw[15]_INST_0_i_285_n_0 ),
        .O(\bdatw[12]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h000E0000000E000E)) 
    \bdatw[12]_INST_0_i_85 
       (.I0(\bdatw[12]_INST_0_i_93_n_0 ),
        .I1(\bdatw[15]_INST_0_i_273_n_0 ),
        .I2(\bdatw[15]_INST_0_i_205_n_0 ),
        .I3(\bdatw[15]_INST_0_i_286_n_0 ),
        .I4(\bdatw[15]_INST_0_i_275_n_0 ),
        .I5(\bdatw[15]_INST_0_i_285_n_0 ),
        .O(\bdatw[12]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \bdatw[12]_INST_0_i_86 
       (.I0(\badr[15]_INST_0_i_296_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [5]),
        .I3(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_14_n_0 ),
        .O(\bdatw[12]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \bdatw[12]_INST_0_i_87 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [8]),
        .O(\bdatw[12]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF088C0002)) 
    \bdatw[12]_INST_0_i_88 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [1]),
        .I4(\stat[2]_i_5__0_n_0 ),
        .I5(\fch/ir1 [7]),
        .O(\bdatw[12]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \bdatw[12]_INST_0_i_89 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [10]),
        .I4(\bdatw[12]_INST_0_i_94_n_0 ),
        .I5(ctl_fetch1_fl_i_17_n_0),
        .O(\bdatw[12]_INST_0_i_89_n_0 ));
  MUXF7 \bdatw[12]_INST_0_i_90 
       (.I0(\bdatw[15]_INST_0_i_211_n_0 ),
        .I1(\bdatw[12]_INST_0_i_95_n_0 ),
        .O(\bdatw[12]_INST_0_i_90_n_0 ),
        .S(\fch/ir1 [11]));
  LUT5 #(
    .INIT(32'h30B003B0)) 
    \bdatw[12]_INST_0_i_91 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [13]),
        .I4(\rgf/sreg/sr [6]),
        .O(\bdatw[12]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h00000002AAAA0002)) 
    \bdatw[12]_INST_0_i_92 
       (.I0(\bdatw[12]_INST_0_i_96_n_0 ),
        .I1(\bcmd[0]_INST_0_i_7_n_0 ),
        .I2(\badr[15]_INST_0_i_214_n_0 ),
        .I3(\bdatw[15]_INST_0_i_208_n_0 ),
        .I4(\fch/ir1 [14]),
        .I5(\rgf/sreg/sr [5]),
        .O(\bdatw[12]_INST_0_i_92_n_0 ));
  LUT4 #(
    .INIT(16'h6FFF)) 
    \bdatw[12]_INST_0_i_93 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .O(\bdatw[12]_INST_0_i_93_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[12]_INST_0_i_94 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .O(\bdatw[12]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h0000A800AAAAAAAA)) 
    \bdatw[12]_INST_0_i_95 
       (.I0(\bdatw[15]_INST_0_i_214_n_0 ),
        .I1(\bdatw[12]_INST_0_i_97_n_0 ),
        .I2(\bdatw[12]_INST_0_i_98_n_0 ),
        .I3(\fch/ir1 [9]),
        .I4(\bdatw[15]_INST_0_i_280_n_0 ),
        .I5(\bdatw[15]_INST_0_i_212_n_0 ),
        .O(\bdatw[12]_INST_0_i_95_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[12]_INST_0_i_96 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [11]),
        .O(\bdatw[12]_INST_0_i_96_n_0 ));
  LUT5 #(
    .INIT(32'h88800880)) 
    \bdatw[12]_INST_0_i_97 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [5]),
        .O(\bdatw[12]_INST_0_i_97_n_0 ));
  LUT4 #(
    .INIT(16'h3BBB)) 
    \bdatw[12]_INST_0_i_98 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .O(\bdatw[12]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[13]_INST_0 
       (.I0(\bdatw[13]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[13]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[13]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[13]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(\bdatw[13]_INST_0_i_4_n_0 ),
        .I1(\bdatw[13]_INST_0_i_5_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[13]_INST_0_i_6_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [13]),
        .I4(\rgf/bank02/p_0_in2_in [13]),
        .I5(\rgf/b0bus_out/bdatw[13]_INST_0_i_9_n_0 ),
        .O(\bdatw[13]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h7555DFFFFDDDDFFF)) 
    \bdatw[13]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(\bdatw[13]_INST_0_i_28_n_0 ),
        .I3(\bdatw[15]_INST_0_i_42_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\fch/ir1 [10]),
        .O(\bdatw[13]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[13]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [13]),
        .O(\bdatw[13]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_16 
       (.I0(\bdatw[13]_INST_0_i_39_n_0 ),
        .I1(\bdatw[13]_INST_0_i_40_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[13]_INST_0_i_41_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_42_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_43_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[13]_INST_0_i_44_n_0 ),
        .O(\bdatw[13]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \bdatw[13]_INST_0_i_17 
       (.I0(\bdatw[15]_INST_0_i_19_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [2]),
        .O(\bdatw[13]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13]_INST_0_i_10_n_0 ),
        .I1(\bdatw[13]_INST_0_i_11_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[13]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_14_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[13]_INST_0_i_15_n_0 ),
        .O(\bdatw[13]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[13]_INST_0_i_27 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [13]),
        .O(\bdatw[13]_INST_0_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_28 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .O(\bdatw[13]_INST_0_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hA3)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\bdatw[13]_INST_0_i_16_n_0 ),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(\bdatw[13]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[13]_INST_0_i_38 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [13]),
        .O(\bdatw[13]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hAA0080AA220080AA)) 
    \bdatw[13]_INST_0_i_39 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(\fch/ir1 [5]),
        .I3(\bdatw[13]_INST_0_i_57_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\fch/ir1 [4]),
        .O(\bdatw[13]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h41414041)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(\bdatw[8]_INST_0_i_5_n_0 ),
        .I1(\bdatw[13]_INST_0_i_17_n_0 ),
        .I2(\bdatw[15]_INST_0_i_22_n_0 ),
        .I3(\bdatw[15]_INST_0_i_19_n_0 ),
        .I4(\fch/ir0 [10]),
        .O(\bdatw[13]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[13]_INST_0_i_40 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [5]),
        .O(\bdatw[13]_INST_0_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_5 
       (.I0(\fch/eir [13]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bdatw[13]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \bdatw[13]_INST_0_i_57 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [0]),
        .O(\bdatw[13]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[13]_INST_0_i_67 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [5]),
        .O(\bdatw[13]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[14]_INST_0 
       (.I0(\bdatw[14]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[14]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[14]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[14]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(\bdatw[14]_INST_0_i_4_n_0 ),
        .I1(\bdatw[14]_INST_0_i_5_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[14]_INST_0_i_6_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [14]),
        .I4(\rgf/bank02/p_0_in2_in [14]),
        .I5(\rgf/b0bus_out/bdatw[14]_INST_0_i_9_n_0 ),
        .O(\bdatw[14]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000200088882888)) 
    \bdatw[14]_INST_0_i_10 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(ctl_selb1_0),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [2]),
        .I4(\bdatw[14]_INST_0_i_29_n_0 ),
        .I5(\bdatw[14]_INST_0_i_30_n_0 ),
        .O(\bdatw[14]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[14]_INST_0_i_11 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [14]),
        .O(\bdatw[14]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_16 
       (.I0(\bdatw[14]_INST_0_i_41_n_0 ),
        .I1(\bdatw[14]_INST_0_i_42_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[14]_INST_0_i_43_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_44_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_45_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[14]_INST_0_i_46_n_0 ),
        .O(\bdatw[14]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[14]_INST_0_i_17 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .O(\bdatw[14]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_18 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [2]),
        .O(\bdatw[14]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(\bdatw[14]_INST_0_i_10_n_0 ),
        .I1(\bdatw[14]_INST_0_i_11_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[14]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[14]_INST_0_i_15_n_0 ),
        .O(\bdatw[14]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[14]_INST_0_i_28 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [14]),
        .O(\bdatw[14]_INST_0_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \bdatw[14]_INST_0_i_29 
       (.I0(\bdatw[15]_INST_0_i_40_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [3]),
        .O(\bdatw[14]_INST_0_i_29_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[14]_INST_0_i_16_n_0 ),
        .O(\bdatw[14]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_30 
       (.I0(\bdatw[15]_INST_0_i_40_n_0 ),
        .I1(\fch/ir1 [10]),
        .O(\bdatw[14]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h000000000030AACF)) 
    \bdatw[14]_INST_0_i_4 
       (.I0(\fch/ir0 [10]),
        .I1(\bdatw[14]_INST_0_i_17_n_0 ),
        .I2(\bdatw[14]_INST_0_i_18_n_0 ),
        .I3(\bdatw[15]_INST_0_i_19_n_0 ),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bdatw[14]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[14]_INST_0_i_40 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [14]),
        .O(\bdatw[14]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h2222A8880022A888)) 
    \bdatw[14]_INST_0_i_41 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[14]_INST_0_i_59_n_0 ),
        .I2(\fch/ir1 [6]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\fch/ir1 [5]),
        .O(\bdatw[14]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[14]_INST_0_i_42 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [6]),
        .O(\bdatw[14]_INST_0_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_5 
       (.I0(\fch/eir [14]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bdatw[14]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \bdatw[14]_INST_0_i_59 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [1]),
        .I4(\bdatw[15]_INST_0_i_40_n_0 ),
        .O(\bdatw[14]_INST_0_i_59_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[14]_INST_0_i_69 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\bdatw[14]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[15]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[15]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[15]_INST_0_i_4_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[15]));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(\bdatw[15]_INST_0_i_6_n_0 ),
        .I1(\bdatw[15]_INST_0_i_7_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[15]_INST_0_i_8_n_0 ),
        .I3(\rgf/bank02/p_1_in3_in [15]),
        .I4(\rgf/bank02/p_0_in2_in [15]),
        .I5(\rgf/b0bus_out/bdatw[15]_INST_0_i_11_n_0 ),
        .O(\bdatw[15]_INST_0_i_1_n_0 ));
  MUXF7 \bdatw[15]_INST_0_i_102 
       (.I0(\bdatw[15]_INST_0_i_203_n_0 ),
        .I1(\bdatw[15]_INST_0_i_204_n_0 ),
        .O(\bdatw[15]_INST_0_i_102_n_0 ),
        .S(\bdatw[15]_INST_0_i_202_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \bdatw[15]_INST_0_i_103 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_103_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF004F)) 
    \bdatw[15]_INST_0_i_104 
       (.I0(\bdatw[15]_INST_0_i_205_n_0 ),
        .I1(\bdatw[15]_INST_0_i_206_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\bdatw[15]_INST_0_i_207_n_0 ),
        .I4(\ctl1/stat [0]),
        .O(\bdatw[15]_INST_0_i_104_n_0 ));
  LUT6 #(
    .INIT(64'hFF40FF00FFFFFF00)) 
    \bdatw[15]_INST_0_i_105 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .I2(\sr[15]_i_8_n_0 ),
        .I3(\badr[15]_INST_0_i_116_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(\bdatw[15]_INST_0_i_208_n_0 ),
        .O(\bdatw[15]_INST_0_i_105_n_0 ));
  MUXF7 \bdatw[15]_INST_0_i_106 
       (.I0(\bdatw[15]_INST_0_i_209_n_0 ),
        .I1(\bdatw[15]_INST_0_i_210_n_0 ),
        .O(\bdatw[15]_INST_0_i_106_n_0 ),
        .S(\fch/ir1 [12]));
  LUT6 #(
    .INIT(64'hEE2E2222FFFFFFFF)) 
    \bdatw[15]_INST_0_i_107 
       (.I0(\bdatw[15]_INST_0_i_211_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\bdatw[15]_INST_0_i_212_n_0 ),
        .I3(\bdatw[15]_INST_0_i_213_n_0 ),
        .I4(\bdatw[15]_INST_0_i_214_n_0 ),
        .I5(\bcmd[1]_INST_0_i_8_n_0 ),
        .O(\bdatw[15]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000BAFE)) 
    \bdatw[15]_INST_0_i_108 
       (.I0(\fch/ir1 [7]),
        .I1(\stat[2]_i_5__0_n_0 ),
        .I2(\bdatw[9]_INST_0_i_65_n_0 ),
        .I3(\bdatw[15]_INST_0_i_208_n_0 ),
        .I4(\bdatw[15]_INST_0_i_215_n_0 ),
        .I5(\bdatw[15]_INST_0_i_216_n_0 ),
        .O(\bdatw[15]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hF0F02020F0002020)) 
    \bdatw[15]_INST_0_i_109 
       (.I0(\bdatw[15]_INST_0_i_217_n_0 ),
        .I1(\bdatw[15]_INST_0_i_218_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\bdatw[15]_INST_0_i_219_n_0 ),
        .I4(\ctl1/stat [0]),
        .I5(\bdatw[15]_INST_0_i_220_n_0 ),
        .O(ctl_selb1_rn[1]));
  LUT6 #(
    .INIT(64'h00000000FFFE0000)) 
    \bdatw[15]_INST_0_i_110 
       (.I0(\bdatw[15]_INST_0_i_221_n_0 ),
        .I1(\bdatw[15]_INST_0_i_222_n_0 ),
        .I2(\ctl1/stat [0]),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bcmd[1]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_224_n_0 ),
        .O(ctl_selb1_rn[0]));
  LUT6 #(
    .INIT(64'h1011FFFF10111011)) 
    \bdatw[15]_INST_0_i_111 
       (.I0(\bdatw[15]_INST_0_i_225_n_0 ),
        .I1(\bdatw[15]_INST_0_i_226_n_0 ),
        .I2(\bdatw[15]_INST_0_i_227_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\bdatw[15]_INST_0_i_228_n_0 ),
        .I5(\bdatw[15]_INST_0_i_229_n_0 ),
        .O(ctl_selb1_rn[2]));
  LUT3 #(
    .INIT(8'hFE)) 
    \bdatw[15]_INST_0_i_112 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(ctl_selb1_0),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .O(\bdatw[15]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'hBABABABABABABAAA)) 
    \bdatw[15]_INST_0_i_116 
       (.I0(ctl_selb1_rn[1]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\bdatw[15]_INST_0_i_116_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDFDFFF)) 
    \bdatw[15]_INST_0_i_117 
       (.I0(ctl_selb1_rn[1]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\bdatw[15]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'h7555DFFFFDDDDFFF)) 
    \bdatw[15]_INST_0_i_12 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(\bdatw[15]_INST_0_i_41_n_0 ),
        .I3(\bdatw[15]_INST_0_i_42_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\fch/ir1 [10]),
        .O(\bdatw[15]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_123 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .O(\bdatw[15]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \bdatw[15]_INST_0_i_127 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\rgf/b1bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \bdatw[15]_INST_0_i_128 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\rgf/b1bus_sel_cr [2]));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \bdatw[15]_INST_0_i_129 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[2]),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\rgf/b1bus_sel_cr [1]));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[15]_INST_0_i_13 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [15]),
        .O(\bdatw[15]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFF7FFFF)) 
    \bdatw[15]_INST_0_i_142 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [0]),
        .O(\bdatw[15]_INST_0_i_142_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[15]_INST_0_i_152 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [7]),
        .O(\bdatw[15]_INST_0_i_152_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FFFF0080)) 
    \bdatw[15]_INST_0_i_153 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [11]),
        .O(\bdatw[15]_INST_0_i_153_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[15]_INST_0_i_154 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .O(\bdatw[15]_INST_0_i_154_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_155 
       (.I0(crdy),
        .I1(\fch/ir0 [8]),
        .O(\bdatw[15]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'h1555155515555555)) 
    \bdatw[15]_INST_0_i_156 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [7]),
        .O(\bdatw[15]_INST_0_i_156_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[15]_INST_0_i_157 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .O(\bdatw[15]_INST_0_i_157_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_158 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [7]),
        .O(\bdatw[15]_INST_0_i_158_n_0 ));
  LUT5 #(
    .INIT(32'h359EFFFF)) 
    \bdatw[15]_INST_0_i_159 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [9]),
        .O(\bdatw[15]_INST_0_i_159_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \bdatw[15]_INST_0_i_160 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .O(\bdatw[15]_INST_0_i_160_n_0 ));
  LUT5 #(
    .INIT(32'h3088FFFF)) 
    \bdatw[15]_INST_0_i_161 
       (.I0(crdy),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [11]),
        .O(\bdatw[15]_INST_0_i_161_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[15]_INST_0_i_162 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [13]),
        .O(\bdatw[15]_INST_0_i_162_n_0 ));
  LUT6 #(
    .INIT(64'h0C000800CF0C8808)) 
    \bdatw[15]_INST_0_i_163 
       (.I0(crdy),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [3]),
        .O(\bdatw[15]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF3003FFFFB4B4)) 
    \bdatw[15]_INST_0_i_164 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [11]),
        .I3(\rgf/sreg/sr [6]),
        .I4(\rgf_selc0_wb[1]_i_36_n_0 ),
        .I5(\fch/ir0 [13]),
        .O(\bdatw[15]_INST_0_i_164_n_0 ));
  LUT5 #(
    .INIT(32'hD5FDFFFF)) 
    \bdatw[15]_INST_0_i_165 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .I4(crdy),
        .O(\bdatw[15]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2A010200)) 
    \bdatw[15]_INST_0_i_166 
       (.I0(\stat[2]_i_6_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [0]),
        .I5(\fch/ir0 [7]),
        .O(\bdatw[15]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hFFFCFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_167 
       (.I0(\fch/ir0 [5]),
        .I1(\bdatw[15]_INST_0_i_253_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\bdatw[15]_INST_0_i_254_n_0 ),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [11]),
        .O(\bdatw[15]_INST_0_i_167_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFF7EFFFF7E)) 
    \bdatw[15]_INST_0_i_168 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [4]),
        .O(\bdatw[15]_INST_0_i_168_n_0 ));
  LUT5 #(
    .INIT(32'hA65656A6)) 
    \bdatw[15]_INST_0_i_169 
       (.I0(\fch/ir0 [11]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir0 [14]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\rgf/sreg/sr [7]),
        .O(\bdatw[15]_INST_0_i_169_n_0 ));
  LUT5 #(
    .INIT(32'h0090FFFF)) 
    \bdatw[15]_INST_0_i_170 
       (.I0(\fch/ir0 [11]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [12]),
        .O(\bdatw[15]_INST_0_i_170_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    \bdatw[15]_INST_0_i_171 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(crdy),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [6]),
        .O(\bdatw[15]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'hFCDDFFDDFCFFCCFF)) 
    \bdatw[15]_INST_0_i_172 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [9]),
        .I2(crdy),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [7]),
        .O(\bdatw[15]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'h00001000FFFFFFFF)) 
    \bdatw[15]_INST_0_i_173 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [5]),
        .I4(\ccmd[4]_INST_0_i_16_n_0 ),
        .I5(\fch/ir0 [9]),
        .O(\bdatw[15]_INST_0_i_173_n_0 ));
  LUT5 #(
    .INIT(32'h5FDDDDDD)) 
    \bdatw[15]_INST_0_i_174 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .I2(\bdatw[15]_INST_0_i_255_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .O(\bdatw[15]_INST_0_i_174_n_0 ));
  LUT5 #(
    .INIT(32'hAA2AAA88)) 
    \bdatw[15]_INST_0_i_175 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [8]),
        .O(\bdatw[15]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA8AAA8AAAAAA)) 
    \bdatw[15]_INST_0_i_176 
       (.I0(\bdatw[15]_INST_0_i_156_n_0 ),
        .I1(\stat[0]_i_32_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [10]),
        .I5(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\bdatw[15]_INST_0_i_176_n_0 ));
  LUT6 #(
    .INIT(64'hFFBA000000000000)) 
    \bdatw[15]_INST_0_i_177 
       (.I0(\bdatw[15]_INST_0_i_186_n_0 ),
        .I1(\bdatw[15]_INST_0_i_256_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\bdatw[15]_INST_0_i_185_n_0 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\fch/ir0 [1]),
        .O(\bdatw[15]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \bdatw[15]_INST_0_i_178 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [7]),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [6]),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\bdatw[15]_INST_0_i_178_n_0 ));
  LUT5 #(
    .INIT(32'h04440004)) 
    \bdatw[15]_INST_0_i_179 
       (.I0(\fadr[15]_INST_0_i_15_n_0 ),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [0]),
        .O(\bdatw[15]_INST_0_i_179_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(\bdatw[15]_INST_0_i_60_n_0 ),
        .I1(\bdatw[15]_INST_0_i_61_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[15]_INST_0_i_62_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_63_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_64_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[15]_INST_0_i_65_n_0 ),
        .O(\bdatw[15]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAABBBBBAAAB)) 
    \bdatw[15]_INST_0_i_180 
       (.I0(\ctl0/stat [0]),
        .I1(\fadr[15]_INST_0_i_15_n_0 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fadr[15]_INST_0_i_14_n_0 ),
        .I4(crdy),
        .I5(\bdatw[15]_INST_0_i_257_n_0 ),
        .O(\bdatw[15]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \bdatw[15]_INST_0_i_181 
       (.I0(\fch/ir0 [7]),
        .I1(\stat[2]_i_10_n_0 ),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [5]),
        .O(\bdatw[15]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'h000000000B0B080B)) 
    \bdatw[15]_INST_0_i_182 
       (.I0(\bdatw[15]_INST_0_i_258_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\bdatw[15]_INST_0_i_259_n_0 ),
        .I3(crdy),
        .I4(\bdatw[15]_INST_0_i_260_n_0 ),
        .I5(\bdatw[15]_INST_0_i_185_n_0 ),
        .O(\bdatw[15]_INST_0_i_182_n_0 ));
  LUT6 #(
    .INIT(64'h00E0E0E0FFFFFFFF)) 
    \bdatw[15]_INST_0_i_183 
       (.I0(\fadr[15]_INST_0_i_15_n_0 ),
        .I1(\bdatw[15]_INST_0_i_257_n_0 ),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [0]),
        .I4(\bdatw[15]_INST_0_i_178_n_0 ),
        .I5(\bcmd[0]_INST_0_i_20_n_0 ),
        .O(\bdatw[15]_INST_0_i_183_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \bdatw[15]_INST_0_i_184 
       (.I0(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I1(\fch/ir0 [2]),
        .I2(\bcmd[1]_INST_0_i_1_n_0 ),
        .I3(\bdatw[15]_INST_0_i_261_n_0 ),
        .I4(\bcmd[0]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_262_n_0 ),
        .O(\bdatw[15]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'h88A8A8888888A8A8)) 
    \bdatw[15]_INST_0_i_185 
       (.I0(\fch/ir0 [6]),
        .I1(\bdatw[15]_INST_0_i_263_n_0 ),
        .I2(\badr[15]_INST_0_i_257_n_0 ),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [4]),
        .O(\bdatw[15]_INST_0_i_185_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888A8A8A8)) 
    \bdatw[15]_INST_0_i_186 
       (.I0(\bdatw[15]_INST_0_i_264_n_0 ),
        .I1(\bdatw[15]_INST_0_i_265_n_0 ),
        .I2(\ccmd[4]_INST_0_i_13_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [8]),
        .O(\bdatw[15]_INST_0_i_186_n_0 ));
  LUT6 #(
    .INIT(64'hFD00550075005500)) 
    \bdatw[15]_INST_0_i_187 
       (.I0(\bdatw[15]_INST_0_i_258_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I5(crdy),
        .O(\bdatw[15]_INST_0_i_187_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \bdatw[15]_INST_0_i_188 
       (.I0(\bcmd[1]_INST_0_i_5_n_0 ),
        .I1(\ctl0/stat [0]),
        .I2(\ctl0/stat [1]),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [2]),
        .O(\bdatw[15]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDFDDDF)) 
    \bdatw[15]_INST_0_i_189 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(\bdatw[15]_INST_0_i_183_n_0 ),
        .I2(\bdatw[15]_INST_0_i_266_n_0 ),
        .I3(\bdatw[15]_INST_0_i_267_n_0 ),
        .I4(\fadr[15]_INST_0_i_15_n_0 ),
        .I5(\ctl0/stat [0]),
        .O(\bdatw[15]_INST_0_i_189_n_0 ));
  LUT6 #(
    .INIT(64'h45FFFFFF0000FFFF)) 
    \bdatw[15]_INST_0_i_19 
       (.I0(\bdatw[15]_INST_0_i_66_n_0 ),
        .I1(\bdatw[15]_INST_0_i_67_n_0 ),
        .I2(\bdatw[15]_INST_0_i_68_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\bcmd[0]_INST_0_i_20_n_0 ),
        .I5(\bdatw[15]_INST_0_i_69_n_0 ),
        .O(\bdatw[15]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBBABAAAAAAAA)) 
    \bdatw[15]_INST_0_i_190 
       (.I0(\ctl0/stat [0]),
        .I1(\bdatw[15]_INST_0_i_268_n_0 ),
        .I2(\bdatw[15]_INST_0_i_175_n_0 ),
        .I3(\bdatw[15]_INST_0_i_269_n_0 ),
        .I4(\bdatw[15]_INST_0_i_72_n_0 ),
        .I5(\stat[2]_i_6_n_0 ),
        .O(\bdatw[15]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2AA0AAAAAAAA)) 
    \bdatw[15]_INST_0_i_191 
       (.I0(\ctl0/stat [0]),
        .I1(\stat[2]_i_6_n_0 ),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [13]),
        .I4(\bdatw[15]_INST_0_i_270_n_0 ),
        .I5(\bdatw[15]_INST_0_i_166_n_0 ),
        .O(\bdatw[15]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888A8AAAA)) 
    \bdatw[15]_INST_0_i_192 
       (.I0(\stat[2]_i_6_n_0 ),
        .I1(\bdatw[15]_INST_0_i_72_n_0 ),
        .I2(\bdatw[15]_INST_0_i_172_n_0 ),
        .I3(\bdatw[15]_INST_0_i_271_n_0 ),
        .I4(\bdatw[15]_INST_0_i_175_n_0 ),
        .I5(\bdatw[15]_INST_0_i_268_n_0 ),
        .O(\bdatw[15]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(\bdatw[15]_INST_0_i_12_n_0 ),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[15]_INST_0_i_14_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_15_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_16_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[15]_INST_0_i_17_n_0 ),
        .O(\bdatw[15]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_20 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .O(\bdatw[15]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h1F0F)) 
    \bdatw[15]_INST_0_i_202 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [13]),
        .I3(\rgf/sreg/sr [6]),
        .O(\bdatw[15]_INST_0_i_202_n_0 ));
  LUT5 #(
    .INIT(32'h8BBBB888)) 
    \bdatw[15]_INST_0_i_203 
       (.I0(\bdatw[15]_INST_0_i_272_n_0 ),
        .I1(\fch/ir1 [14]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [11]),
        .O(\bdatw[15]_INST_0_i_203_n_0 ));
  LUT6 #(
    .INIT(64'hC03F3FC050AF50AF)) 
    \bdatw[15]_INST_0_i_204 
       (.I0(\rgf/sreg/sr [4]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [11]),
        .I4(\rgf/sreg/sr [5]),
        .I5(\fch/ir1 [14]),
        .O(\bdatw[15]_INST_0_i_204_n_0 ));
  LUT6 #(
    .INIT(64'h6666447466764474)) 
    \bdatw[15]_INST_0_i_205 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [7]),
        .O(\bdatw[15]_INST_0_i_205_n_0 ));
  LUT5 #(
    .INIT(32'hBFFFFFBF)) 
    \bdatw[15]_INST_0_i_206 
       (.I0(\bdatw[15]_INST_0_i_273_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [9]),
        .O(\bdatw[15]_INST_0_i_206_n_0 ));
  LUT6 #(
    .INIT(64'h04FF04FF04FF0404)) 
    \bdatw[15]_INST_0_i_207 
       (.I0(\bdatw[15]_INST_0_i_274_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [11]),
        .I3(\bdatw[15]_INST_0_i_275_n_0 ),
        .I4(\fch/ir1 [10]),
        .I5(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .O(\bdatw[15]_INST_0_i_207_n_0 ));
  LUT4 #(
    .INIT(16'hF773)) 
    \bdatw[15]_INST_0_i_208 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [1]),
        .O(\bdatw[15]_INST_0_i_208_n_0 ));
  LUT6 #(
    .INIT(64'h0F00CF35000FCF35)) 
    \bdatw[15]_INST_0_i_209 
       (.I0(\bdatw[15]_INST_0_i_276_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [14]),
        .I5(\rgf/sreg/sr [5]),
        .O(\bdatw[15]_INST_0_i_209_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_21 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [2]),
        .O(\bdatw[15]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01010100)) 
    \bdatw[15]_INST_0_i_210 
       (.I0(\bcmd[0]_INST_0_i_24_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\stat[0]_i_13__0_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\bdatw[15]_INST_0_i_277_n_0 ),
        .O(\bdatw[15]_INST_0_i_210_n_0 ));
  LUT6 #(
    .INIT(64'h33F13FF1FFFFFFFF)) 
    \bdatw[15]_INST_0_i_211 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_211_n_0 ));
  LUT5 #(
    .INIT(32'hFFFAFF3F)) 
    \bdatw[15]_INST_0_i_212 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_212_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022F20000)) 
    \bdatw[15]_INST_0_i_213 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\bdatw[15]_INST_0_i_278_n_0 ),
        .I2(\bdatw[15]_INST_0_i_279_n_0 ),
        .I3(ctl_fetch1_fl_i_12_n_0),
        .I4(\fch/ir1 [9]),
        .I5(\bdatw[15]_INST_0_i_280_n_0 ),
        .O(\bdatw[15]_INST_0_i_213_n_0 ));
  LUT4 #(
    .INIT(16'hBFEE)) 
    \bdatw[15]_INST_0_i_214 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_214_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFF8)) 
    \bdatw[15]_INST_0_i_215 
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [2]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [13]),
        .I4(\bdatw[15]_INST_0_i_281_n_0 ),
        .I5(\badr[15]_INST_0_i_296_n_0 ),
        .O(\bdatw[15]_INST_0_i_215_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA8AAAAAAAA)) 
    \bdatw[15]_INST_0_i_216 
       (.I0(\stat[1]_i_5__0_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [12]),
        .I5(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .O(\bdatw[15]_INST_0_i_216_n_0 ));
  LUT6 #(
    .INIT(64'h10005555FFFFFFFF)) 
    \bdatw[15]_INST_0_i_217 
       (.I0(\bdatw[15]_INST_0_i_282_n_0 ),
        .I1(\bdatw[15]_INST_0_i_283_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(ctl_fetch1_fl_i_11_n_0),
        .I5(\fch/ir1 [11]),
        .O(\bdatw[15]_INST_0_i_217_n_0 ));
  LUT6 #(
    .INIT(64'h55557757FFFFFFFF)) 
    \bdatw[15]_INST_0_i_218 
       (.I0(\bdatw[15]_INST_0_i_284_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\bdatw[15]_INST_0_i_285_n_0 ),
        .I3(\bdatw[15]_INST_0_i_275_n_0 ),
        .I4(\bdatw[15]_INST_0_i_286_n_0 ),
        .I5(\bcmd[1]_INST_0_i_8_n_0 ),
        .O(\bdatw[15]_INST_0_i_218_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \bdatw[15]_INST_0_i_219 
       (.I0(\badr[15]_INST_0_i_296_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [5]),
        .I3(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_208_n_0 ),
        .O(\bdatw[15]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBAFFFAFAF)) 
    \bdatw[15]_INST_0_i_22 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[15]_INST_0_i_71_n_0 ),
        .I2(\stat[2]_i_6_n_0 ),
        .I3(\bdatw[15]_INST_0_i_72_n_0 ),
        .I4(\bdatw[15]_INST_0_i_73_n_0 ),
        .I5(\ctl0/stat [0]),
        .O(\bdatw[15]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \bdatw[15]_INST_0_i_220 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [11]),
        .I3(\bcmd[1]_INST_0_i_8_n_0 ),
        .I4(\fch/ir1 [9]),
        .I5(\bdatw[15]_INST_0_i_287_n_0 ),
        .O(\bdatw[15]_INST_0_i_220_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF088C0000)) 
    \bdatw[15]_INST_0_i_221 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [1]),
        .I4(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I5(\badr[15]_INST_0_i_116_n_0 ),
        .O(\bdatw[15]_INST_0_i_221_n_0 ));
  LUT6 #(
    .INIT(64'h0000000039040004)) 
    \bdatw[15]_INST_0_i_222 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [0]),
        .I5(\bdatw[15]_INST_0_i_288_n_0 ),
        .O(\bdatw[15]_INST_0_i_222_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \bdatw[15]_INST_0_i_223 
       (.I0(\bdatw[15]_INST_0_i_225_n_0 ),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [0]),
        .I5(\bdatw[15]_INST_0_i_289_n_0 ),
        .O(\bdatw[15]_INST_0_i_223_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0B0B0B000B0B0)) 
    \bdatw[15]_INST_0_i_224 
       (.I0(\bdatw[15]_INST_0_i_208_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I2(\ctl1/stat [0]),
        .I3(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I4(\fch/ir1 [0]),
        .I5(\bdatw[15]_INST_0_i_290_n_0 ),
        .O(\bdatw[15]_INST_0_i_224_n_0 ));
  LUT6 #(
    .INIT(64'h00F100F1000000F1)) 
    \bdatw[15]_INST_0_i_225 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\bdatw[15]_INST_0_i_275_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [6]),
        .I5(\bdatw[15]_INST_0_i_274_n_0 ),
        .O(\bdatw[15]_INST_0_i_225_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_226 
       (.I0(\fch/ir1 [15]),
        .I1(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat [2]),
        .I4(\fch/ir1 [2]),
        .I5(\badr[15]_INST_0_i_144_n_0 ),
        .O(\bdatw[15]_INST_0_i_226_n_0 ));
  LUT6 #(
    .INIT(64'h7030FFCC33330FFF)) 
    \bdatw[15]_INST_0_i_227 
       (.I0(\bdatw[15]_INST_0_i_283_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_227_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_228 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [12]),
        .I4(\bdatw[15]_INST_0_i_291_n_0 ),
        .I5(\bcmd[1]_INST_0_i_3_n_0 ),
        .O(\bdatw[15]_INST_0_i_228_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \bdatw[15]_INST_0_i_229 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [9]),
        .O(\bdatw[15]_INST_0_i_229_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_23 
       (.I0(ctl_selb0_rn[1]),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_76_n_0 ),
        .I3(\bdatw[15]_INST_0_i_77_n_0 ),
        .O(\rgf/b0bus_sel_cr [4]));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[15]_INST_0_i_230 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[1]),
        .O(\bdatw[15]_INST_0_i_230_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDFDFFF)) 
    \bdatw[15]_INST_0_i_231 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\bdatw[15]_INST_0_i_231_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAAAAAAAAAAAAA)) 
    \bdatw[15]_INST_0_i_232 
       (.I0(\ctl1/stat [0]),
        .I1(\stat[0]_i_30__0_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\bcmd[1]_INST_0_i_8_n_0 ),
        .I5(\bdatw[15]_INST_0_i_292_n_0 ),
        .O(\bdatw[15]_INST_0_i_232_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_233 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[2]),
        .O(\bdatw[15]_INST_0_i_233_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_238 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .O(\bdatw[15]_INST_0_i_238_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_24 
       (.I0(ctl_selb0_rn[1]),
        .I1(ctl_selb0_rn[0]),
        .I2(\bdatw[15]_INST_0_i_76_n_0 ),
        .I3(\bdatw[15]_INST_0_i_77_n_0 ),
        .O(\rgf/b0bus_sel_cr [3]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_253 
       (.I0(\ctl0/stat [1]),
        .I1(\ctl0/stat [2]),
        .O(\bdatw[15]_INST_0_i_253_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[15]_INST_0_i_254 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .O(\bdatw[15]_INST_0_i_254_n_0 ));
  LUT3 #(
    .INIT(8'h43)) 
    \bdatw[15]_INST_0_i_255 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [4]),
        .O(\bdatw[15]_INST_0_i_255_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF505000F03838)) 
    \bdatw[15]_INST_0_i_256 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(crdy),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [9]),
        .O(\bdatw[15]_INST_0_i_256_n_0 ));
  LUT4 #(
    .INIT(16'hD4FF)) 
    \bdatw[15]_INST_0_i_257 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [2]),
        .O(\bdatw[15]_INST_0_i_257_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0C64)) 
    \bdatw[15]_INST_0_i_258 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .O(\bdatw[15]_INST_0_i_258_n_0 ));
  LUT6 #(
    .INIT(64'h2000200030000000)) 
    \bdatw[15]_INST_0_i_259 
       (.I0(crdy),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [11]),
        .I4(\ccmd[4]_INST_0_i_17_n_0 ),
        .I5(\fch/ir0 [8]),
        .O(\bdatw[15]_INST_0_i_259_n_0 ));
  LUT6 #(
    .INIT(64'h0FFFC4D53FFFC4D5)) 
    \bdatw[15]_INST_0_i_260 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [7]),
        .O(\bdatw[15]_INST_0_i_260_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_261 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [6]),
        .O(\bdatw[15]_INST_0_i_261_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_262 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [11]),
        .O(\bdatw[15]_INST_0_i_262_n_0 ));
  LUT6 #(
    .INIT(64'h000000E000000000)) 
    \bdatw[15]_INST_0_i_263 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(crdy),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\bdatw[15]_INST_0_i_263_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_264 
       (.I0(crdy),
        .I1(\fch/ir0 [11]),
        .O(\bdatw[15]_INST_0_i_264_n_0 ));
  LUT5 #(
    .INIT(32'hC000B030)) 
    \bdatw[15]_INST_0_i_265 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [9]),
        .O(\bdatw[15]_INST_0_i_265_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA888888888)) 
    \bdatw[15]_INST_0_i_266 
       (.I0(\bcmd[1]_INST_0_i_5_n_0 ),
        .I1(\bdatw[15]_INST_0_i_181_n_0 ),
        .I2(\bdatw[15]_INST_0_i_185_n_0 ),
        .I3(\bdatw[15]_INST_0_i_186_n_0 ),
        .I4(\bdatw[15]_INST_0_i_187_n_0 ),
        .I5(\fch/ir0 [0]),
        .O(\bdatw[15]_INST_0_i_266_n_0 ));
  LUT6 #(
    .INIT(64'h00C0C0CC00000050)) 
    \bdatw[15]_INST_0_i_267 
       (.I0(\pc0[15]_i_3_n_0 ),
        .I1(crdy),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [2]),
        .O(\bdatw[15]_INST_0_i_267_n_0 ));
  LUT6 #(
    .INIT(64'hFF1F0000FFFFFFFF)) 
    \bdatw[15]_INST_0_i_268 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [6]),
        .I3(\rgf_selc0_wb[1]_i_38_n_0 ),
        .I4(\bdatw[15]_INST_0_i_156_n_0 ),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\bdatw[15]_INST_0_i_268_n_0 ));
  LUT6 #(
    .INIT(64'h8AAA8A8A8AAA8AAA)) 
    \bdatw[15]_INST_0_i_269 
       (.I0(\bdatw[15]_INST_0_i_172_n_0 ),
        .I1(\bdatw[15]_INST_0_i_295_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\bdatw[15]_INST_0_i_296_n_0 ),
        .I4(\bdatw[15]_INST_0_i_255_n_0 ),
        .I5(\bdatw[15]_INST_0_i_158_n_0 ),
        .O(\bdatw[15]_INST_0_i_269_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF6FF6)) 
    \bdatw[15]_INST_0_i_270 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .I4(\bdatw[15]_INST_0_i_297_n_0 ),
        .I5(\bdatw[15]_INST_0_i_168_n_0 ),
        .O(\bdatw[15]_INST_0_i_270_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BABB0000)) 
    \bdatw[15]_INST_0_i_271 
       (.I0(\bdatw[15]_INST_0_i_298_n_0 ),
        .I1(\ccmd[4]_INST_0_i_22_n_0 ),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .I5(\bdatw[15]_INST_0_i_295_n_0 ),
        .O(\bdatw[15]_INST_0_i_271_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF9FFFF)) 
    \bdatw[15]_INST_0_i_272 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [5]),
        .I2(\badr[15]_INST_0_i_311_n_0 ),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [11]),
        .I5(\stat[1]_i_19_n_0 ),
        .O(\bdatw[15]_INST_0_i_272_n_0 ));
  LUT5 #(
    .INIT(32'hE2490000)) 
    \bdatw[15]_INST_0_i_273 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [9]),
        .O(\bdatw[15]_INST_0_i_273_n_0 ));
  LUT4 #(
    .INIT(16'h777F)) 
    \bdatw[15]_INST_0_i_274 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [9]),
        .O(\bdatw[15]_INST_0_i_274_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEEE)) 
    \bdatw[15]_INST_0_i_275 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .O(\bdatw[15]_INST_0_i_275_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[15]_INST_0_i_276 
       (.I0(\bdatw[15]_INST_0_i_208_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [8]),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\bdatw[15]_INST_0_i_276_n_0 ));
  LUT6 #(
    .INIT(64'h0A0A050559A9A959)) 
    \bdatw[15]_INST_0_i_277 
       (.I0(\fch/ir1 [11]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [14]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\fch/ir1 [13]),
        .O(\bdatw[15]_INST_0_i_277_n_0 ));
  LUT3 #(
    .INIT(8'h43)) 
    \bdatw[15]_INST_0_i_278 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [4]),
        .O(\bdatw[15]_INST_0_i_278_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_279 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_279_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \bdatw[15]_INST_0_i_280 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_280_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_281 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_281_n_0 ));
  LUT6 #(
    .INIT(64'h31117555755D75F5)) 
    \bdatw[15]_INST_0_i_282 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [10]),
        .O(\bdatw[15]_INST_0_i_282_n_0 ));
  LUT3 #(
    .INIT(8'hC6)) 
    \bdatw[15]_INST_0_i_283 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [5]),
        .O(\bdatw[15]_INST_0_i_283_n_0 ));
  LUT3 #(
    .INIT(8'hCE)) 
    \bdatw[15]_INST_0_i_284 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_284_n_0 ));
  LUT6 #(
    .INIT(64'hABAAAAAAAAAAAAAA)) 
    \bdatw[15]_INST_0_i_285 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [12]),
        .O(\bdatw[15]_INST_0_i_285_n_0 ));
  LUT6 #(
    .INIT(64'h4440000000000000)) 
    \bdatw[15]_INST_0_i_286 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_286_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_287 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_287_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_288 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [7]),
        .I5(\bcmd[1]_INST_0_i_8_n_0 ),
        .O(\bdatw[15]_INST_0_i_288_n_0 ));
  LUT6 #(
    .INIT(64'h8BC8000098D80000)) 
    \bdatw[15]_INST_0_i_289 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [7]),
        .O(\bdatw[15]_INST_0_i_289_n_0 ));
  LUT5 #(
    .INIT(32'hFBFFFFFF)) 
    \bdatw[15]_INST_0_i_290 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\bcmd[1]_INST_0_i_8_n_0 ),
        .I4(\fch/ir1 [11]),
        .O(\bdatw[15]_INST_0_i_290_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_291 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_291_n_0 ));
  LUT5 #(
    .INIT(32'h08800388)) 
    \bdatw[15]_INST_0_i_292 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [4]),
        .O(\bdatw[15]_INST_0_i_292_n_0 ));
  LUT6 #(
    .INIT(64'h44444440FFFFFFFF)) 
    \bdatw[15]_INST_0_i_293 
       (.I0(\bdatw[15]_INST_0_i_224_n_0 ),
        .I1(\bcmd[1]_INST_0_i_3_n_0 ),
        .I2(\bdatw[15]_INST_0_i_223_n_0 ),
        .I3(\bdatw[15]_INST_0_i_232_n_0 ),
        .I4(\bdatw[15]_INST_0_i_221_n_0 ),
        .I5(ctl_selb1_rn[1]),
        .O(\bdatw[15]_INST_0_i_293_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFFF)) 
    \bdatw[15]_INST_0_i_294 
       (.I0(ctl_selb1_rn[1]),
        .I1(\bdatw[15]_INST_0_i_224_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\bdatw[15]_INST_0_i_223_n_0 ),
        .I4(\bdatw[15]_INST_0_i_232_n_0 ),
        .I5(\bdatw[15]_INST_0_i_221_n_0 ),
        .O(\bdatw[15]_INST_0_i_294_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \bdatw[15]_INST_0_i_295 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [4]),
        .O(\bdatw[15]_INST_0_i_295_n_0 ));
  LUT4 #(
    .INIT(16'h3BBB)) 
    \bdatw[15]_INST_0_i_296 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .O(\bdatw[15]_INST_0_i_296_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEFEEEFFFFFEEE)) 
    \bdatw[15]_INST_0_i_297 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\ctl0/stat [1]),
        .I3(\ctl0/stat [2]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [10]),
        .O(\bdatw[15]_INST_0_i_297_n_0 ));
  LUT5 #(
    .INIT(32'h88800880)) 
    \bdatw[15]_INST_0_i_298 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [5]),
        .O(\bdatw[15]_INST_0_i_298_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(bcmd[1]),
        .I1(bcmd[2]),
        .O(\bdatw[15]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_38 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [15]),
        .O(\bdatw[15]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0000010001010101)) 
    \bdatw[15]_INST_0_i_39 
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [1]),
        .I3(\fch/ir1 [15]),
        .I4(\bcmd[1]_INST_0_i_8_n_0 ),
        .I5(\bdatw[15]_INST_0_i_102_n_0 ),
        .O(\bdatw[15]_INST_0_i_39_n_0 ));
  LUT3 #(
    .INIT(8'hA3)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(\bbus_o[7]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_18_n_0 ),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(\bdatw[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0070007000FFFFFF)) 
    \bdatw[15]_INST_0_i_40 
       (.I0(\bdatw[15]_INST_0_i_103_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I2(\bdatw[15]_INST_0_i_104_n_0 ),
        .I3(\bdatw[15]_INST_0_i_105_n_0 ),
        .I4(\bcmd[1]_INST_0_i_3_n_0 ),
        .I5(\bcmd[2]_INST_0_i_4_n_0 ),
        .O(\bdatw[15]_INST_0_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_41 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .O(\bdatw[15]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_42 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [0]),
        .O(\bdatw[15]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A008A)) 
    \bdatw[15]_INST_0_i_43 
       (.I0(\stat[2]_i_5__0_n_0 ),
        .I1(\bdatw[15]_INST_0_i_106_n_0 ),
        .I2(\bdatw[15]_INST_0_i_107_n_0 ),
        .I3(\ctl1/stat [0]),
        .I4(\bdatw[15]_INST_0_i_108_n_0 ),
        .I5(\fch/ir1 [15]),
        .O(ctl_selb1_0));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[15]_INST_0_i_44 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .O(\rgf/b1bus_sel_cr [4]));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_45 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .O(\rgf/b1bus_sel_cr [3]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_5 
       (.I0(bcmd[2]),
        .I1(bcmd[1]),
        .O(\bdatw[15]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[15]_INST_0_i_59 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [15]),
        .O(\bdatw[15]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h0000000030008BBB)) 
    \bdatw[15]_INST_0_i_6 
       (.I0(\fch/ir0 [10]),
        .I1(\bdatw[15]_INST_0_i_19_n_0 ),
        .I2(\bdatw[15]_INST_0_i_20_n_0 ),
        .I3(\bdatw[15]_INST_0_i_21_n_0 ),
        .I4(\bdatw[15]_INST_0_i_22_n_0 ),
        .I5(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bdatw[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAA0080AA220080AA)) 
    \bdatw[15]_INST_0_i_60 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(\fch/ir1 [7]),
        .I3(\bdatw[15]_INST_0_i_142_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[15]_INST_0_i_61 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [7]),
        .O(\bdatw[15]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \bdatw[15]_INST_0_i_66 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [10]),
        .O(\bdatw[15]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hBBFBFFFFAAAAAAAA)) 
    \bdatw[15]_INST_0_i_67 
       (.I0(\ctl0/stat [0]),
        .I1(\bdatw[15]_INST_0_i_153_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\bdatw[15]_INST_0_i_154_n_0 ),
        .I4(\bdatw[15]_INST_0_i_155_n_0 ),
        .I5(\bdatw[15]_INST_0_i_156_n_0 ),
        .O(\bdatw[15]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4040FF40)) 
    \bdatw[15]_INST_0_i_68 
       (.I0(\bdatw[15]_INST_0_i_157_n_0 ),
        .I1(\bdatw[15]_INST_0_i_158_n_0 ),
        .I2(\bdatw[15]_INST_0_i_159_n_0 ),
        .I3(\ccmd[4]_INST_0_i_17_n_0 ),
        .I4(\bdatw[15]_INST_0_i_160_n_0 ),
        .I5(\bdatw[15]_INST_0_i_161_n_0 ),
        .O(\bdatw[15]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFFFDFFFDFD)) 
    \bdatw[15]_INST_0_i_69 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_5_n_0 ),
        .I2(\bdatw[15]_INST_0_i_162_n_0 ),
        .I3(\bdatw[15]_INST_0_i_163_n_0 ),
        .I4(\fadr[15]_INST_0_i_14_n_0 ),
        .I5(\pc0[15]_i_3_n_0 ),
        .O(\bdatw[15]_INST_0_i_69_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(\fch/eir [15]),
        .I1(\bdatw[10]_INST_0_i_5_n_0 ),
        .O(\bdatw[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBBA)) 
    \bdatw[15]_INST_0_i_70 
       (.I0(\fch/ir0 [15]),
        .I1(\bdatw[15]_INST_0_i_164_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [14]),
        .I5(\bdatw[15]_INST_0_i_165_n_0 ),
        .O(\bdatw[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0200000200000002)) 
    \bdatw[15]_INST_0_i_71 
       (.I0(\bdatw[15]_INST_0_i_166_n_0 ),
        .I1(\bdatw[15]_INST_0_i_167_n_0 ),
        .I2(\bdatw[15]_INST_0_i_168_n_0 ),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [14]),
        .I5(\stat[2]_i_6_n_0 ),
        .O(\bdatw[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1F1F1FFFFFFF1)) 
    \bdatw[15]_INST_0_i_72 
       (.I0(\bdatw[15]_INST_0_i_169_n_0 ),
        .I1(\fch/ir0 [13]),
        .I2(\bdatw[15]_INST_0_i_170_n_0 ),
        .I3(\ccmd[4]_INST_0_i_13_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I5(\bdatw[15]_INST_0_i_171_n_0 ),
        .O(\bdatw[15]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7500FFFF)) 
    \bdatw[15]_INST_0_i_73 
       (.I0(\bdatw[15]_INST_0_i_172_n_0 ),
        .I1(\bdatw[15]_INST_0_i_173_n_0 ),
        .I2(\bdatw[15]_INST_0_i_174_n_0 ),
        .I3(\bdatw[15]_INST_0_i_175_n_0 ),
        .I4(\bcmd[0]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_176_n_0 ),
        .O(\bdatw[15]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCC8C8C000C8C8)) 
    \bdatw[15]_INST_0_i_74 
       (.I0(\bdatw[15]_INST_0_i_177_n_0 ),
        .I1(\bcmd[0]_INST_0_i_20_n_0 ),
        .I2(\bdatw[15]_INST_0_i_178_n_0 ),
        .I3(\fch/ir0 [1]),
        .I4(\ctl0/stat [0]),
        .I5(\bdatw[15]_INST_0_i_179_n_0 ),
        .O(ctl_selb0_rn[1]));
  LUT6 #(
    .INIT(64'h00000000EAEEEAEA)) 
    \bdatw[15]_INST_0_i_75 
       (.I0(\bdatw[15]_INST_0_i_180_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\bdatw[15]_INST_0_i_181_n_0 ),
        .I3(\bdatw[15]_INST_0_i_182_n_0 ),
        .I4(\fch/ir0 [0]),
        .I5(\bdatw[15]_INST_0_i_183_n_0 ),
        .O(ctl_selb0_rn[0]));
  LUT6 #(
    .INIT(64'h4444444455555554)) 
    \bdatw[15]_INST_0_i_76 
       (.I0(\ctl0/stat [2]),
        .I1(\bdatw[15]_INST_0_i_184_n_0 ),
        .I2(\bdatw[15]_INST_0_i_185_n_0 ),
        .I3(\bdatw[15]_INST_0_i_186_n_0 ),
        .I4(\bdatw[15]_INST_0_i_187_n_0 ),
        .I5(\bdatw[15]_INST_0_i_188_n_0 ),
        .O(\bdatw[15]_INST_0_i_76_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \bdatw[15]_INST_0_i_77 
       (.I0(\bdatw[15]_INST_0_i_22_n_0 ),
        .I1(\bdatw[15]_INST_0_i_19_n_0 ),
        .I2(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bdatw[15]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    \bdatw[15]_INST_0_i_80 
       (.I0(\bdatw[15]_INST_0_i_76_n_0 ),
        .I1(\bdatw[8]_INST_0_i_5_n_0 ),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\bdatw[15]_INST_0_i_190_n_0 ),
        .I4(\bdatw[15]_INST_0_i_191_n_0 ),
        .I5(\bdatw[15]_INST_0_i_70_n_0 ),
        .O(\bdatw[15]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBBAFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_81 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[15]_INST_0_i_71_n_0 ),
        .I2(\bdatw[15]_INST_0_i_192_n_0 ),
        .I3(\ctl0/stat [0]),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bdatw[15]_INST_0_i_81_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[1]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[9]_INST_0_i_3_n_0 ),
        .O(bdatw[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[2]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[10]_INST_0_i_3_n_0 ),
        .O(bdatw[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[3]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[11]_INST_0_i_3_n_0 ),
        .O(bdatw[3]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[4]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[12]_INST_0_i_3_n_0 ),
        .O(bdatw[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[5]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[13]_INST_0_i_3_n_0 ),
        .O(bdatw[5]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[6]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[14]_INST_0_i_3_n_0 ),
        .O(bdatw[6]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[7]_INST_0 
       (.I0(bcmd[1]),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(bdatw[7]));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[8]_INST_0 
       (.I0(\bdatw[8]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[8]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[8]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[8]));
  LUT6 #(
    .INIT(64'h000000000000DD0D)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(\bdatw[8]_INST_0_i_4_n_0 ),
        .I1(\bdatw[8]_INST_0_i_5_n_0 ),
        .I2(\fch/eir [8]),
        .I3(\bdatw[10]_INST_0_i_5_n_0 ),
        .I4(\rgf/b0bus_out/bdatw[8]_INST_0_i_6_n_0 ),
        .I5(\rgf/b0bus_out/bdatw[8]_INST_0_i_7_n_0 ),
        .O(\bdatw[8]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[8]_INST_0_i_14 
       (.I0(\bdatw[8]_INST_0_i_35_n_0 ),
        .I1(\bdatw[8]_INST_0_i_36_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[8]_INST_0_i_37_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_38_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[8]_INST_0_i_40_n_0 ),
        .O(\bdatw[8]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[8]_INST_0_i_15 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [2]),
        .O(\bdatw[8]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hC03F3FC050AF50AF)) 
    \bdatw[8]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [4]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(\rgf/sreg/sr [5]),
        .I5(\fch/ir0 [14]),
        .O(\bdatw[8]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h04FF)) 
    \bdatw[8]_INST_0_i_17 
       (.I0(\fch/ir0 [14]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [13]),
        .O(\bdatw[8]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFEFEFF)) 
    \bdatw[8]_INST_0_i_18 
       (.I0(\bdatw[8]_INST_0_i_41_n_0 ),
        .I1(\bdatw[8]_INST_0_i_42_n_0 ),
        .I2(\bdatw[8]_INST_0_i_43_n_0 ),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [5]),
        .I5(\bdatw[8]_INST_0_i_44_n_0 ),
        .O(\bdatw[8]_INST_0_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bdatw[8]_INST_0_i_19 
       (.I0(\ctl0/stat [0]),
        .I1(\ctl0/stat [1]),
        .I2(\ctl0/stat [2]),
        .O(\bdatw[8]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_8_n_0 ),
        .I1(\bdatw[8]_INST_0_i_9_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[8]_INST_0_i_10_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_11_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_12_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[8]_INST_0_i_13_n_0 ),
        .O(\bdatw[8]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\bdatw[8]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[8]_INST_0_i_34 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\bdatw[8]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFF0233FDFFFFFFFF)) 
    \bdatw[8]_INST_0_i_35 
       (.I0(\bdatw[8]_INST_0_i_59_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [1]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bdatw[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[8]_INST_0_i_36 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [0]),
        .O(\bdatw[8]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455A55555)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_22_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .I4(\bdatw[8]_INST_0_i_15_n_0 ),
        .I5(\bdatw[15]_INST_0_i_19_n_0 ),
        .O(\bdatw[8]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \bdatw[8]_INST_0_i_41 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [12]),
        .O(\bdatw[8]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[8]_INST_0_i_42 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [7]),
        .O(\bdatw[8]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \bdatw[8]_INST_0_i_43 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [6]),
        .O(\bdatw[8]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h5F5D555F555D5F5F)) 
    \bdatw[8]_INST_0_i_44 
       (.I0(\fch/ir0 [13]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [11]),
        .I5(\rgf/sreg/sr [7]),
        .O(\bdatw[8]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hF800F8F8FFFFFFFF)) 
    \bdatw[8]_INST_0_i_5 
       (.I0(\bdatw[8]_INST_0_i_16_n_0 ),
        .I1(\bdatw[8]_INST_0_i_17_n_0 ),
        .I2(\bdatw[8]_INST_0_i_18_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\fch/ir0 [15]),
        .I5(\bdatw[8]_INST_0_i_19_n_0 ),
        .O(\bdatw[8]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[8]_INST_0_i_59 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [3]),
        .O(\bdatw[8]_INST_0_i_59_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[8]_INST_0_i_73 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\rgf/sreg/sr [0]),
        .O(\bdatw[8]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_78 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr03 [0]),
        .O(\bdatw[8]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_79 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr04 [0]),
        .O(\bdatw[8]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'h75DF75DFFFDF75DF)) 
    \bdatw[8]_INST_0_i_8 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[14]_INST_0_i_29_n_0 ),
        .I2(\bdatw[9]_INST_0_i_20_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\bdatw[15]_INST_0_i_40_n_0 ),
        .I5(\fch/ir1 [7]),
        .O(\bdatw[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[8]_INST_0_i_80 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr07 [0]),
        .O(\bdatw[8]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_81 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr06 [0]),
        .O(\bdatw[8]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_82 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr23 [0]),
        .O(\bdatw[8]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_83 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr24 [0]),
        .O(\bdatw[8]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[8]_INST_0_i_84 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr27 [0]),
        .O(\bdatw[8]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[8]_INST_0_i_85 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [0]),
        .O(\bdatw[8]_INST_0_i_85_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [8]),
        .O(\bdatw[8]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \bdatw[9]_INST_0 
       (.I0(\bdatw[9]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\bdatw[9]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_3_n_0 ),
        .I4(\bdatw[9]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[9]));
  LUT5 #(
    .INIT(32'h00000051)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(\bdatw[9]_INST_0_i_4_n_0 ),
        .I1(\fch/eir [9]),
        .I2(\bdatw[10]_INST_0_i_5_n_0 ),
        .I3(\rgf/b0bus_out/bdatw[9]_INST_0_i_5_n_0 ),
        .I4(\rgf/b0bus_out/bdatw[9]_INST_0_i_6_n_0 ),
        .O(\bdatw[9]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \bdatw[9]_INST_0_i_13 
       (.I0(\bdatw[9]_INST_0_i_31_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[9]_INST_0_i_32_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_33_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_34_n_0 ),
        .I4(\rgf/b1bus_out/bdatw[9]_INST_0_i_35_n_0 ),
        .I5(\bdatw[9]_INST_0_i_36_n_0 ),
        .O(\bdatw[9]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \bdatw[9]_INST_0_i_14 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .I2(\bdatw[15]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [0]),
        .O(\bdatw[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(\bdatw[9]_INST_0_i_7_n_0 ),
        .I1(\bdatw[9]_INST_0_i_8_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[9]_INST_0_i_9_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_10_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_11_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[9]_INST_0_i_12_n_0 ),
        .O(\bdatw[9]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[9]_INST_0_i_20 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .O(\bdatw[9]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(\bdatw[9]_INST_0_i_13_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(\bdatw[9]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[9]_INST_0_i_30 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_112_n_0 ),
        .I4(\rgf/sreg/sr [9]),
        .O(\bdatw[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[9]_INST_0_i_31 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [1]),
        .O(\bdatw[9]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h221DEE1DFFFFFFFF)) 
    \bdatw[9]_INST_0_i_36 
       (.I0(\bdatw[9]_INST_0_i_65_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(\fch/ir1 [1]),
        .I3(ctl_selb1_0),
        .I4(\fch/ir1 [0]),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bdatw[9]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h0000F00D)) 
    \bdatw[9]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_19_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\bdatw[15]_INST_0_i_22_n_0 ),
        .I3(\bdatw[9]_INST_0_i_14_n_0 ),
        .I4(\bdatw[8]_INST_0_i_5_n_0 ),
        .O(\bdatw[9]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \bdatw[9]_INST_0_i_64 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\bdatw[15]_INST_0_i_112_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(\rgf/sreg/sr [1]),
        .O(\bdatw[9]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[9]_INST_0_i_65 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [0]),
        .O(\bdatw[9]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h08F7F8F7FFFFFFFF)) 
    \bdatw[9]_INST_0_i_7 
       (.I0(\bdatw[9]_INST_0_i_20_n_0 ),
        .I1(\bdatw[15]_INST_0_i_42_n_0 ),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\fch/ir1 [8]),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bdatw[9]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_70 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr03 [1]),
        .O(\bdatw[9]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_71 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr04 [1]),
        .O(\bdatw[9]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[9]_INST_0_i_72 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr07 [1]),
        .O(\bdatw[9]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_73 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr06 [1]),
        .O(\bdatw[9]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_74 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr23 [1]),
        .O(\bdatw[9]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_75 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_233_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr24 [1]),
        .O(\bdatw[9]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[9]_INST_0_i_76 
       (.I0(ctl_selb1_rn[2]),
        .I1(\bdatw[15]_INST_0_i_39_n_0 ),
        .I2(\bdatw[12]_INST_0_i_79_n_0 ),
        .I3(\bdatw[15]_INST_0_i_117_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr27 [1]),
        .O(\bdatw[9]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[9]_INST_0_i_77 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[12]_INST_0_i_79_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_230_n_0 ),
        .I4(\rgf/bank_sel [3]),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\bdatw[9]_INST_0_i_77_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[9]_INST_0_i_8 
       (.I0(\bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\bdatw[15]_INST_0_i_40_n_0 ),
        .I2(ctl_selb1_0),
        .I3(\fch/eir [9]),
        .O(\bdatw[9]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(ccmd[0]));
  LUT6 #(
    .INIT(64'h00F4FFF4FFF4FFF4)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(\ccmd[0]_INST_0_i_2_n_0 ),
        .I1(\ccmd[0]_INST_0_i_3_n_0 ),
        .I2(\ccmd[0]_INST_0_i_4_n_0 ),
        .I3(\ccmd[0]_INST_0_i_5_n_0 ),
        .I4(\ccmd[0]_INST_0_i_6_n_0 ),
        .I5(\ccmd[0]_INST_0_i_7_n_0 ),
        .O(\ccmd[0]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [0]),
        .O(\ccmd[0]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [14]),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h5FCFA0CF)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [14]),
        .I4(\rgf/sreg/sr [5]),
        .O(\ccmd[0]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7F7C4F7)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(\ccmd[0]_INST_0_i_24_n_0 ),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [9]),
        .I3(\ccmd[0]_INST_0_i_25_n_0 ),
        .I4(\ctl0/stat [1]),
        .I5(\ccmd[0]_INST_0_i_26_n_0 ),
        .O(\ccmd[0]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [11]),
        .O(\ccmd[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4000400000004000)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(\ccmd[4]_INST_0_i_17_n_0 ),
        .I1(\ccmd[0]_INST_0_i_27_n_0 ),
        .I2(\bcmd[0]_INST_0_i_19_n_0 ),
        .I3(\ccmd[0]_INST_0_i_28_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [8]),
        .O(\ccmd[0]_INST_0_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h54)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [6]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hCFFFAAFFFFFFFFAA)) 
    \ccmd[0]_INST_0_i_19 
       (.I0(\ccmd[0]_INST_0_i_29_n_0 ),
        .I1(\ccmd[0]_INST_0_i_22_n_0 ),
        .I2(\ccmd[0]_INST_0_i_30_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAAAAAAAAAAA)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(\ccmd[0]_INST_0_i_8_n_0 ),
        .I1(\ccmd[0]_INST_0_i_9_n_0 ),
        .I2(\ccmd[0]_INST_0_i_10_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\ccmd[0]_INST_0_i_11_n_0 ),
        .I5(\ccmd[0]_INST_0_i_12_n_0 ),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \ccmd[0]_INST_0_i_20 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [3]),
        .O(\ccmd[0]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[0]_INST_0_i_21 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .O(\ccmd[0]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[0]_INST_0_i_22 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [4]),
        .O(\ccmd[0]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[0]_INST_0_i_23 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .O(\ccmd[0]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hC03F1000000C0000)) 
    \ccmd[0]_INST_0_i_24 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\ctl0/stat [1]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [7]),
        .O(\ccmd[0]_INST_0_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hC7)) 
    \ccmd[0]_INST_0_i_25 
       (.I0(\fch/ir0 [12]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [11]),
        .O(\ccmd[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FCAA0000)) 
    \ccmd[0]_INST_0_i_26 
       (.I0(\ccmd[0]_INST_0_i_31_n_0 ),
        .I1(\ccmd[0]_INST_0_i_32_n_0 ),
        .I2(\ccmd[0]_INST_0_i_33_n_0 ),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [14]),
        .I5(\ctl0/stat [1]),
        .O(\ccmd[0]_INST_0_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_27 
       (.I0(\fch/ir0 [10]),
        .I1(\ctl0/stat [1]),
        .O(\ccmd[0]_INST_0_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_28 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [4]),
        .O(\ccmd[0]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_29 
       (.I0(\fch/ir0 [7]),
        .I1(crdy),
        .O(\ccmd[0]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAABBAAEEEBBBEEEE)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [15]),
        .I4(\ccmd[0]_INST_0_i_13_n_0 ),
        .I5(\fch/ir0 [12]),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_30 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [3]),
        .O(\ccmd[0]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h2020202022222A22)) 
    \ccmd[0]_INST_0_i_31 
       (.I0(\ccmd[0]_INST_0_i_34_n_0 ),
        .I1(\ccmd[0]_INST_0_i_35_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [4]),
        .I5(\ccmd[0]_INST_0_i_36_n_0 ),
        .O(\ccmd[0]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h00BB000B00200000)) 
    \ccmd[0]_INST_0_i_32 
       (.I0(crdy),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[0]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000240000)) 
    \ccmd[0]_INST_0_i_33 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [7]),
        .I3(\ccmd[0]_INST_0_i_28_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\ccmd[4]_INST_0_i_16_n_0 ),
        .O(\ccmd[0]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hEFEECFCCEFEECCCC)) 
    \ccmd[0]_INST_0_i_34 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\ccmd[0]_INST_0_i_35_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I4(crdy),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[0]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hA0A2AAAAA0A2A0A2)) 
    \ccmd[0]_INST_0_i_35 
       (.I0(\fch/ir0 [8]),
        .I1(crdy),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\ccmd[0]_INST_0_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0_i_36 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [5]),
        .O(\ccmd[0]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA8A8A888A)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(\ccmd[0]_INST_0_i_8_n_0 ),
        .I1(\ccmd[0]_INST_0_i_14_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\ccmd[0]_INST_0_i_15_n_0 ),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [15]),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h0000FB00)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(\fch/ir0 [7]),
        .I1(\ctl0/stat [1]),
        .I2(\fch/ir0 [2]),
        .I3(\ctl0/stat [0]),
        .I4(\ccmd[0]_INST_0_i_16_n_0 ),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000880000FFFC)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(\ccmd[0]_INST_0_i_17_n_0 ),
        .I1(\ccmd[0]_INST_0_i_18_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [15]),
        .I5(\ctl0/stat [1]),
        .O(\ccmd[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4444444400000F00)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(\ccmd[0]_INST_0_i_19_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\ccmd[0]_INST_0_i_20_n_0 ),
        .I3(\ccmd[0]_INST_0_i_21_n_0 ),
        .I4(\ccmd[0]_INST_0_i_22_n_0 ),
        .I5(\fch/ir0 [10]),
        .O(\ccmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FB00)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(\fch/ir0 [12]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [13]),
        .I4(\ctl0/stat [1]),
        .I5(\fch/ir0 [15]),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\ccmd[0]_INST_0_i_22_n_0 ),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [9]),
        .I5(\ccmd[0]_INST_0_i_23_n_0 ),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[1]_INST_0 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'h000000002222FF0F)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_3_n_0 ),
        .I2(\ccmd[1]_INST_0_i_4_n_0 ),
        .I3(\ccmd[1]_INST_0_i_5_n_0 ),
        .I4(\ccmd[1]_INST_0_i_6_n_0 ),
        .I5(\ctl0/stat [1]),
        .O(\ccmd[1]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FFFFFF01)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [11]),
        .I2(\ccmd[1]_INST_0_i_19_n_0 ),
        .I3(\ccmd[1]_INST_0_i_20_n_0 ),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [13]),
        .O(\ccmd[1]_INST_0_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [2]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [4]),
        .O(\ccmd[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFDFFFF)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [11]),
        .I4(\ccmd[1]_INST_0_i_21_n_0 ),
        .I5(\ccmd[1]_INST_0_i_22_n_0 ),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFF7)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [9]),
        .I3(\ctl0/stat [0]),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000100FFFFFFFF)) 
    \ccmd[1]_INST_0_i_15 
       (.I0(\ccmd[4]_INST_0_i_22_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\ctl0/stat [0]),
        .I3(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I4(\badrx[15]_INST_0_i_4_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0A1FFFFFFFFFFFFF)) 
    \ccmd[1]_INST_0_i_16 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(crdy),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [8]),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\ccmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0010000033330030)) 
    \ccmd[1]_INST_0_i_17 
       (.I0(\fch/ir0 [7]),
        .I1(\ccmd[1]_INST_0_i_23_n_0 ),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [5]),
        .O(\ccmd[1]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h2215F215)) 
    \ccmd[1]_INST_0_i_18 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [7]),
        .I4(crdy),
        .O(\ccmd[1]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[1]_INST_0_i_19 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [1]),
        .O(\ccmd[1]_INST_0_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(\fch/ir0 [14]),
        .I1(\ctl0/stat [2]),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_20 
       (.I0(\ctl0/stat [2]),
        .I1(\ctl0/stat [0]),
        .O(\ccmd[1]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[1]_INST_0_i_21 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [15]),
        .O(\ccmd[1]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_22 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [5]),
        .O(\ccmd[1]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFF7FFF7FFFFF)) 
    \ccmd[1]_INST_0_i_23 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [7]),
        .O(\ccmd[1]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFABABFF00FFFF)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(\ccmd[1]_INST_0_i_7_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\ccmd[1]_INST_0_i_8_n_0 ),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [15]),
        .I5(\fch/ir0 [13]),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF51005555)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(\ccmd[1]_INST_0_i_9_n_0 ),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [15]),
        .I5(\ccmd[1]_INST_0_i_10_n_0 ),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000D0D00)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(\fadr[15]_INST_0_i_14_n_0 ),
        .I1(\ccmd[1]_INST_0_i_11_n_0 ),
        .I2(\ccmd[1]_INST_0_i_12_n_0 ),
        .I3(\fch/ir0 [2]),
        .I4(\ctl0/stat [2]),
        .I5(\ccmd[1]_INST_0_i_13_n_0 ),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [15]),
        .O(\ccmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000FB0000)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(\ccmd[1]_INST_0_i_14_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\ccmd[1]_INST_0_i_15_n_0 ),
        .I4(\ccmd[1]_INST_0_i_16_n_0 ),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\ccmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000400F400040000)) 
    \ccmd[1]_INST_0_i_8 
       (.I0(\stat[0]_i_8__1_n_0 ),
        .I1(crdy),
        .I2(\ctl0/stat [0]),
        .I3(\ccmd[1]_INST_0_i_18_n_0 ),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\ccmd[4]_INST_0_i_14_n_0 ),
        .O(\ccmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [8]),
        .I4(crdy),
        .I5(\ccmd[4]_INST_0_i_20_n_0 ),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0 
       (.I0(\ccmd[2]_INST_0_i_1_n_0 ),
        .I1(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(ccmd[2]));
  LUT6 #(
    .INIT(64'h000000000020FFFF)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(\ccmd[2]_INST_0_i_2_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\ctl0/stat [0]),
        .I3(\ctl0/stat [1]),
        .I4(\ctl0/stat [2]),
        .I5(\ccmd[2]_INST_0_i_3_n_0 ),
        .O(\ccmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hEE04FFFFFFFFFFFF)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(\ctl0/stat [1]),
        .I1(\ccmd[2]_INST_0_i_13_n_0 ),
        .I2(crdy),
        .I3(\ccmd[2]_INST_0_i_14_n_0 ),
        .I4(\ccmd[2]_INST_0_i_15_n_0 ),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\ccmd[2]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA80000AAA8)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(\ccmd[2]_INST_0_i_16_n_0 ),
        .I1(\ccmd[2]_INST_0_i_17_n_0 ),
        .I2(\ccmd[2]_INST_0_i_18_n_0 ),
        .I3(\badr[15]_INST_0_i_202_n_0 ),
        .I4(\bcmd[2]_INST_0_i_7_n_0 ),
        .I5(\ccmd[3]_INST_0_i_8_n_0 ),
        .O(\ccmd[2]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAEAAAAAAAA)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(\rgf_selc0_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\ccmd[0]_INST_0_i_23_n_0 ),
        .I4(\ccmd[2]_INST_0_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFCFFFCCCBFFCBFCC)) 
    \ccmd[2]_INST_0_i_13 
       (.I0(\ccmd[2]_INST_0_i_19_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [6]),
        .O(\ccmd[2]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \ccmd[2]_INST_0_i_14 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .O(\ccmd[2]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[2]_INST_0_i_15 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [15]),
        .O(\ccmd[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hDDCCFDDFDDCCDDDD)) 
    \ccmd[2]_INST_0_i_16 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\ccmd[2]_INST_0_i_20_n_0 ),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [7]),
        .O(\ccmd[2]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \ccmd[2]_INST_0_i_17 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [7]),
        .I2(\ccmd[0]_INST_0_i_22_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [13]),
        .O(\ccmd[2]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFEFFFEFFFFF)) 
    \ccmd[2]_INST_0_i_18 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [8]),
        .I4(\ctl0/stat [0]),
        .I5(crdy),
        .O(\ccmd[2]_INST_0_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hD6)) 
    \ccmd[2]_INST_0_i_19 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .O(\ccmd[2]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(\fadr[15]_INST_0_i_14_n_0 ),
        .I1(\ccmd[2]_INST_0_i_4_n_0 ),
        .I2(\ccmd[2]_INST_0_i_5_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .I5(\ccmd[2]_INST_0_i_6_n_0 ),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \ccmd[2]_INST_0_i_20 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [15]),
        .I2(\bcmd[0]_INST_0_i_26_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(crdy),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\ccmd[2]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(\ccmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\ccmd[2]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [5]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  MUXF7 \ccmd[2]_INST_0_i_7 
       (.I0(\ccmd[2]_INST_0_i_9_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\ccmd[2]_INST_0_i_7_n_0 ),
        .S(\fch/ir0 [11]));
  LUT6 #(
    .INIT(64'h5545555545554545)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(\rgf_selc0_wb[1]_i_5_n_0 ),
        .I1(\ccmd[3]_INST_0_i_8_n_0 ),
        .I2(\stat[2]_i_6_n_0 ),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [12]),
        .I5(\fch/ir0 [13]),
        .O(\ccmd[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0EEEEFFFFEEEE)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(\stat[0]_i_14__1_n_0 ),
        .I1(\ccmd[2]_INST_0_i_11_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\fch/ir0 [15]),
        .I4(\ctl0/stat [1]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\ccmd[2]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(ccmd[3]));
  LUT6 #(
    .INIT(64'h0D0D0D0D0F0F0F00)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(\ccmd[3]_INST_0_i_2_n_0 ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(\ccmd[3]_INST_0_i_4_n_0 ),
        .I3(\ccmd[3]_INST_0_i_5_n_0 ),
        .I4(\fch/ir0 [15]),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [4]),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0100010067660000)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [3]),
        .I2(\ctl0/stat [0]),
        .I3(\ctl0/stat [1]),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [0]),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000022E0000)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(crdy),
        .I1(\ctl0/stat [1]),
        .I2(\ctl0/stat [0]),
        .I3(\ccmd[4]_INST_0_i_13_n_0 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .O(\ccmd[3]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0004540000000000)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [6]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [9]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h04040000040400FF)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I1(\ccmd[4]_INST_0_i_19_n_0 ),
        .I2(\ctl0/stat [0]),
        .I3(\ccmd[1]_INST_0_i_14_n_0 ),
        .I4(\ctl0/stat [1]),
        .I5(\ccmd[3]_INST_0_i_16_n_0 ),
        .O(\ccmd[3]_INST_0_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(crdy),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .O(\ccmd[3]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .O(\ccmd[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF08000000)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\ctl0/stat [1]),
        .I3(\fch/ir0 [10]),
        .I4(\ccmd[3]_INST_0_i_6_n_0 ),
        .I5(\ccmd[3]_INST_0_i_7_n_0 ),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [15]),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00050007000A0000)) 
    \ccmd[3]_INST_0_i_4 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [11]),
        .I2(\ctl0/stat [1]),
        .I3(\ccmd[3]_INST_0_i_8_n_0 ),
        .I4(\fch/ir0 [12]),
        .I5(\fch/ir0 [14]),
        .O(\ccmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFA8AA)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(\ccmd[3]_INST_0_i_9_n_0 ),
        .I1(\ccmd[3]_INST_0_i_10_n_0 ),
        .I2(\ccmd[4]_INST_0_i_12_n_0 ),
        .I3(\ccmd[3]_INST_0_i_11_n_0 ),
        .I4(\fch/ir0 [10]),
        .I5(\ccmd[3]_INST_0_i_12_n_0 ),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hBFAFBAAA)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(\ccmd[3]_INST_0_i_13_n_0 ),
        .I1(\ctl0/stat [0]),
        .I2(\fch/ir0 [9]),
        .I3(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I4(crdy),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000060)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\ccmd[4]_INST_0_i_8_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [9]),
        .I5(\ccmd[3]_INST_0_i_14_n_0 ),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [15]),
        .O(\ccmd[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hEFFBFFFFFFFFFFFF)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(\ccmd[3]_INST_0_i_15_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\ccmd[4]_INST_0_i_8_n_0 ),
        .I5(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(ccmd[4]));
  LUT6 #(
    .INIT(64'h1011101010111011)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(\fch/ir0 [15]),
        .I1(\ctl0/stat [2]),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(\ccmd[4]_INST_0_i_5_n_0 ),
        .O(\ccmd[4]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFE00000000000000)) 
    \ccmd[4]_INST_0_i_10 
       (.I0(\ctl0/stat [1]),
        .I1(crdy),
        .I2(\ccmd[4]_INST_0_i_18_n_0 ),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [11]),
        .I5(\ccmd[4]_INST_0_i_19_n_0 ),
        .O(\ccmd[4]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0110011303330333)) 
    \ccmd[4]_INST_0_i_11 
       (.I0(\fch/ir0 [0]),
        .I1(\ccmd[4]_INST_0_i_20_n_0 ),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [3]),
        .I4(\ctl0/stat [0]),
        .I5(\ctl0/stat [1]),
        .O(\ccmd[4]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFEFEFF)) 
    \ccmd[4]_INST_0_i_12 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [12]),
        .I3(\ctl0/stat [0]),
        .I4(crdy),
        .I5(\ctl0/stat [1]),
        .O(\ccmd[4]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \ccmd[4]_INST_0_i_13 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [12]),
        .O(\ccmd[4]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \ccmd[4]_INST_0_i_14 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .O(\ccmd[4]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFBBBBBBBBBBBBBBB)) 
    \ccmd[4]_INST_0_i_15 
       (.I0(\ccmd[4]_INST_0_i_21_n_0 ),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [9]),
        .I4(\ccmd[4]_INST_0_i_22_n_0 ),
        .I5(\ccmd[4]_INST_0_i_8_n_0 ),
        .O(\ccmd[4]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_16 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .O(\ccmd[4]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_17 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .O(\ccmd[4]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0_i_18 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [7]),
        .O(\ccmd[4]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0_i_19 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[4]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF3D3FFDF)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(\ccmd[4]_INST_0_i_6_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [12]),
        .I3(\ccmd[4]_INST_0_i_7_n_0 ),
        .I4(\ccmd[4]_INST_0_i_8_n_0 ),
        .I5(\ccmd[4]_INST_0_i_9_n_0 ),
        .O(\ccmd[4]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \ccmd[4]_INST_0_i_20 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [2]),
        .O(\ccmd[4]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00000000FDD5)) 
    \ccmd[4]_INST_0_i_21 
       (.I0(crdy),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .I4(\ctl0/stat [0]),
        .I5(\ctl0/stat [1]),
        .O(\ccmd[4]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[4]_INST_0_i_22 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .O(\ccmd[4]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h2A22000000000000)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(\ccmd[4]_INST_0_i_10_n_0 ),
        .I1(\ctl0/stat [1]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [10]),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\ccmd[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(\ccmd[4]_INST_0_i_11_n_0 ),
        .I1(\ccmd[4]_INST_0_i_12_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [4]),
        .O(\ccmd[4]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF03707777)) 
    \ccmd[4]_INST_0_i_5 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(crdy),
        .I2(\ctl0/stat [1]),
        .I3(\fch/ir0 [7]),
        .I4(\ccmd[4]_INST_0_i_14_n_0 ),
        .I5(\ccmd[4]_INST_0_i_15_n_0 ),
        .O(\ccmd[4]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAB)) 
    \ccmd[4]_INST_0_i_6 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\ccmd[4]_INST_0_i_16_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\ctl0/stat [1]),
        .I4(\ctl0/stat [0]),
        .I5(\ccmd[4]_INST_0_i_17_n_0 ),
        .O(\ccmd[4]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFF0000EFFF000000)) 
    \ccmd[4]_INST_0_i_7 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [10]),
        .I2(\ccmd[4]_INST_0_i_17_n_0 ),
        .I3(\ctl0/stat [1]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [9]),
        .O(\ccmd[4]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[4]_INST_0_i_8 
       (.I0(\ctl0/stat [1]),
        .I1(\ctl0/stat [0]),
        .O(\ccmd[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF44FFFFFFFFF)) 
    \ccmd[4]_INST_0_i_9 
       (.I0(crdy),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [15]),
        .I4(\ctl0/stat [2]),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\ccmd[4]_INST_0_i_9_n_0 ));
  FDRE \ctl0/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl0/stat_nx [0]),
        .Q(\ctl0/stat [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \ctl0/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl0/stat_nx [1]),
        .Q(\ctl0/stat [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \ctl0/stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl0/stat_nx [2]),
        .Q(\ctl0/stat [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \ctl1/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl1/stat_nx [0]),
        .Q(\ctl1/stat [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \ctl1/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl1/stat_nx [1]),
        .Q(\ctl1/stat [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \ctl1/stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl1/stat_nx [2]),
        .Q(\ctl1/stat [2]),
        .R(\rgf/treg/p_0_in ));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take0_fl_i_1
       (.I0(\ctl0/stat [1]),
        .I1(\ctl0/stat [0]),
        .I2(\ctl0/stat [2]),
        .I3(\fch/ctl_bcc_take0_fl ),
        .O(ctl_bcc_take0_fl_i_1_n_0));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take1_fl_i_1
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [1]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ctl_bcc_take1_fl ),
        .O(ctl_bcc_take1_fl_i_1_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAA2AAAAAAAA)) 
    ctl_fetch0_fl_i_1
       (.I0(ctl_fetch0_fl_i_2_n_0),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\ctl0/stat [2]),
        .I3(\fch/ir0 [15]),
        .I4(brdy),
        .I5(ctl_fetch0_fl_i_3_n_0),
        .O(ctl_fetch0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_10
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [5]),
        .O(ctl_fetch0_fl_i_10_n_0));
  LUT5 #(
    .INIT(32'hDFFFAAAA)) 
    ctl_fetch0_fl_i_11
       (.I0(\fch/ir0 [1]),
        .I1(\rgf/sreg/sr [10]),
        .I2(crdy),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [2]),
        .O(ctl_fetch0_fl_i_11_n_0));
  LUT3 #(
    .INIT(8'h04)) 
    ctl_fetch0_fl_i_12
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [2]),
        .O(ctl_fetch0_fl_i_12_n_0));
  LUT5 #(
    .INIT(32'hBB2B0000)) 
    ctl_fetch0_fl_i_13
       (.I0(irq_lev[1]),
        .I1(\rgf/sreg/sr [3]),
        .I2(\rgf/sreg/sr [2]),
        .I3(irq_lev[0]),
        .I4(irq),
        .O(ctl_fetch0_fl_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    ctl_fetch0_fl_i_14
       (.I0(\stat[1]_i_23_n_0 ),
        .I1(ctl_fetch0_fl_i_28_n_0),
        .I2(\stat[1]_i_24_n_0 ),
        .I3(\bdatw[15]_INST_0_i_20_n_0 ),
        .I4(\fch/ir0 [7]),
        .I5(\ccmd[0]_INST_0_i_22_n_0 ),
        .O(ctl_fetch0_fl_i_14_n_0));
  LUT6 #(
    .INIT(64'hFAFFFAFFEEEEFEFF)) 
    ctl_fetch0_fl_i_15
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .I2(\ctl0/stat [0]),
        .I3(\bcmd[0]_INST_0_i_19_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .I5(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'hB8FFFFFFB800FFFF)) 
    ctl_fetch0_fl_i_16
       (.I0(ctl_fetch0_fl_i_29_n_0),
        .I1(\fch/ir0 [14]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [13]),
        .I5(\rgf/sreg/sr [6]),
        .O(ctl_fetch0_fl_i_16_n_0));
  LUT6 #(
    .INIT(64'h0C0C08080F0F0800)) 
    ctl_fetch0_fl_i_17
       (.I0(\ctl0/stat [0]),
        .I1(crdy),
        .I2(ctl_fetch0_fl_i_30_n_0),
        .I3(\rgf/sreg/sr [10]),
        .I4(\fch/ir0 [8]),
        .I5(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(ctl_fetch0_fl_i_17_n_0));
  LUT6 #(
    .INIT(64'h0000333001333110)) 
    ctl_fetch0_fl_i_18
       (.I0(\ctl0/stat [1]),
        .I1(ctl_fetch0_fl_i_31_n_0),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [0]),
        .I5(\fch/ir0 [3]),
        .O(ctl_fetch0_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'hEFEFEFEFFFEFEFEF)) 
    ctl_fetch0_fl_i_19
       (.I0(\ccmd[0]_INST_0_i_9_n_0 ),
        .I1(ctl_fetch0_fl_i_32_n_0),
        .I2(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .I3(\ctl0/stat [1]),
        .I4(\ctl0/stat [0]),
        .I5(\ccmd[0]_INST_0_i_11_n_0 ),
        .O(ctl_fetch0_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'hF0F0F4F4FFF0F4F4)) 
    ctl_fetch0_fl_i_2
       (.I0(ctl_fetch0_fl_i_4_n_0),
        .I1(ctl_fetch0_fl_i_5_n_0),
        .I2(ctl_fetch0_fl_i_6_n_0),
        .I3(ctl_fetch0_fl_i_7_n_0),
        .I4(\fch/ir0 [11]),
        .I5(ctl_fetch0_fl_i_8_n_0),
        .O(ctl_fetch0_fl_i_2_n_0));
  LUT6 #(
    .INIT(64'h4040404455555555)) 
    ctl_fetch0_fl_i_20
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\bcmd[0]_INST_0_i_19_n_0 ),
        .I2(\ctl0/stat [1]),
        .I3(\stat[0]_i_8__1_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I5(ctl_fetch0_fl_i_33_n_0),
        .O(ctl_fetch0_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF7FF74)) 
    ctl_fetch0_fl_i_21
       (.I0(\fch/ir0 [12]),
        .I1(\bcmd[0]_INST_0_i_19_n_0 ),
        .I2(\ctl0/stat [1]),
        .I3(\ctl0/stat [2]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [15]),
        .O(ctl_fetch0_fl_i_21_n_0));
  LUT6 #(
    .INIT(64'h77777F7F7777777F)) 
    ctl_fetch0_fl_i_22
       (.I0(\bcmd[0]_INST_0_i_19_n_0 ),
        .I1(crdy),
        .I2(ctl_fetch0_fl_i_34_n_0),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFDDDDDCCC)) 
    ctl_fetch0_fl_i_23
       (.I0(\fch/ir0 [10]),
        .I1(\ctl0/stat [1]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [9]),
        .I4(\ctl0/stat [0]),
        .I5(ctl_fetch0_fl_i_35_n_0),
        .O(ctl_fetch0_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'hFFDFFFFFFDFCFFFF)) 
    ctl_fetch0_fl_i_24
       (.I0(\fch/ir0 [3]),
        .I1(ctl_fetch0_fl_i_36_n_0),
        .I2(\fch/ir0 [6]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [5]),
        .O(ctl_fetch0_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'hABABFFAFAAAAAAAA)) 
    ctl_fetch0_fl_i_25
       (.I0(ctl_fetch0_fl_i_37_n_0),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [10]),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(ctl_fetch0_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAAAFFFF)) 
    ctl_fetch0_fl_i_26
       (.I0(ctl_fetch0_fl_i_38_n_0),
        .I1(\fch/ir0 [8]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [6]),
        .I4(\stat[2]_i_6_n_0 ),
        .I5(ctl_fetch0_fl_i_39_n_0),
        .O(ctl_fetch0_fl_i_26_n_0));
  LUT6 #(
    .INIT(64'h700F0FFFFF0F0FFF)) 
    ctl_fetch0_fl_i_27
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [7]),
        .O(ctl_fetch0_fl_i_27_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_28
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .O(ctl_fetch0_fl_i_28_n_0));
  LUT4 #(
    .INIT(16'h8088)) 
    ctl_fetch0_fl_i_29
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(crdy),
        .I3(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(ctl_fetch0_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'hAAEAAAAAAAAAAAAA)) 
    ctl_fetch0_fl_i_3
       (.I0(ctl_fetch0_fl_i_9_n_0),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [3]),
        .I3(\ctl0/stat [1]),
        .I4(ctl_fetch0_fl_i_10_n_0),
        .I5(\stat[2]_i_10_n_0 ),
        .O(ctl_fetch0_fl_i_3_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    ctl_fetch0_fl_i_30
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .O(ctl_fetch0_fl_i_30_n_0));
  LUT6 #(
    .INIT(64'hECEFA0A0ECECA0A0)) 
    ctl_fetch0_fl_i_31
       (.I0(\ctl0/stat [2]),
        .I1(\fch/ir0 [3]),
        .I2(\ctl0/stat [1]),
        .I3(\rgf/sreg/sr [10]),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [2]),
        .O(ctl_fetch0_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hE0E0E0E0FFE0E0E0)) 
    ctl_fetch0_fl_i_32
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [2]),
        .I2(\ctl0/stat [2]),
        .I3(\fch/ir0 [3]),
        .I4(\rgf/sreg/sr [10]),
        .I5(\ctl0/stat [1]),
        .O(ctl_fetch0_fl_i_32_n_0));
  LUT3 #(
    .INIT(8'h8F)) 
    ctl_fetch0_fl_i_33
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [7]),
        .I2(\ctl0/stat [0]),
        .O(ctl_fetch0_fl_i_33_n_0));
  LUT5 #(
    .INIT(32'h0CACFFAC)) 
    ctl_fetch0_fl_i_34
       (.I0(\fch/ir0 [12]),
        .I1(\ctl0/stat [1]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [9]),
        .O(ctl_fetch0_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'h000000001F1FFF1F)) 
    ctl_fetch0_fl_i_35
       (.I0(\rgf/sreg/sr [11]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\ctl0/stat [0]),
        .I4(\rgf/sreg/sr [10]),
        .I5(ctl_fetch0_fl_i_40_n_0),
        .O(ctl_fetch0_fl_i_35_n_0));
  LUT4 #(
    .INIT(16'h4FFF)) 
    ctl_fetch0_fl_i_36
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_36_n_0));
  LUT6 #(
    .INIT(64'h0909090900000900)) 
    ctl_fetch0_fl_i_37
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [13]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [12]),
        .O(ctl_fetch0_fl_i_37_n_0));
  LUT6 #(
    .INIT(64'h00034444FFFFFFFF)) 
    ctl_fetch0_fl_i_38
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir0 [12]),
        .I5(ctl_fetch0_fl_i_33_n_0),
        .O(ctl_fetch0_fl_i_38_n_0));
  LUT5 #(
    .INIT(32'h040404C4)) 
    ctl_fetch0_fl_i_39
       (.I0(\rgf/sreg/sr [6]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir0 [14]),
        .O(ctl_fetch0_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00AE)) 
    ctl_fetch0_fl_i_4
       (.I0(ctl_fetch0_fl_i_11_n_0),
        .I1(ctl_fetch0_fl_i_12_n_0),
        .I2(ctl_fetch0_fl_i_13_n_0),
        .I3(ctl_fetch0_fl_i_14_n_0),
        .I4(\badrx[15]_INST_0_i_4_n_0 ),
        .I5(ctl_fetch0_fl_i_15_n_0),
        .O(ctl_fetch0_fl_i_4_n_0));
  LUT5 #(
    .INIT(32'h1011FFFF)) 
    ctl_fetch0_fl_i_40
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\rgf/sreg/sr [11]),
        .I4(\fch/ir0 [10]),
        .O(ctl_fetch0_fl_i_40_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0E000000)) 
    ctl_fetch0_fl_i_5
       (.I0(\ccmd[0]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [13]),
        .I2(\ctl0/stat [2]),
        .I3(\ccmd[4]_INST_0_i_8_n_0 ),
        .I4(ctl_fetch0_fl_i_16_n_0),
        .I5(ctl_fetch0_fl_i_17_n_0),
        .O(ctl_fetch0_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'hDDD0FFFFDDD0DDD0)) 
    ctl_fetch0_fl_i_6
       (.I0(ctl_fetch0_fl_i_18_n_0),
        .I1(ctl_fetch0_fl_i_19_n_0),
        .I2(ctl_fetch0_fl_i_20_n_0),
        .I3(ctl_fetch0_fl_i_21_n_0),
        .I4(ctl_fetch0_fl_i_22_n_0),
        .I5(ctl_fetch0_fl_i_23_n_0),
        .O(ctl_fetch0_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF9000)) 
    ctl_fetch0_fl_i_7
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .I2(\bcmd[0]_INST_0_i_19_n_0 ),
        .I3(ctl_fetch0_fl_i_24_n_0),
        .I4(ctl_fetch0_fl_i_25_n_0),
        .I5(ctl_fetch0_fl_i_26_n_0),
        .O(ctl_fetch0_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000090000000000)) 
    ctl_fetch0_fl_i_8
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [13]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir0 [14]),
        .I5(\bdatw[8]_INST_0_i_19_n_0 ),
        .O(ctl_fetch0_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'h00000000002A0155)) 
    ctl_fetch0_fl_i_9
       (.I0(\fch/ir0 [9]),
        .I1(\ctl0/stat [0]),
        .I2(\fch/ir0 [6]),
        .I3(\ctl0/stat [1]),
        .I4(\fch/ir0 [8]),
        .I5(ctl_fetch0_fl_i_27_n_0),
        .O(ctl_fetch0_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'h0455045504550404)) 
    ctl_fetch1_fl_i_1
       (.I0(ctl_fetch1_fl_i_2_n_0),
        .I1(brdy),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .I3(ctl_fetch1_fl_i_3_n_0),
        .I4(ctl_fetch1_fl_i_4_n_0),
        .I5(ctl_fetch1_fl_i_5_n_0),
        .O(ctl_fetch1));
  LUT6 #(
    .INIT(64'hFFFFFFFF444444F4)) 
    ctl_fetch1_fl_i_10
       (.I0(ctl_fetch1_fl_i_18_n_0),
        .I1(ctl_fetch1_fl_i_19_n_0),
        .I2(ctl_fetch1_fl_i_20_n_0),
        .I3(ctl_fetch1_fl_i_21_n_0),
        .I4(\bcmd[0]_INST_0_i_24_n_0 ),
        .I5(ctl_fetch1_fl_i_22_n_0),
        .O(ctl_fetch1_fl_i_10_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_11
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .O(ctl_fetch1_fl_i_11_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch1_fl_i_12
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .O(ctl_fetch1_fl_i_12_n_0));
  LUT6 #(
    .INIT(64'h2AAA55FF55555555)) 
    ctl_fetch1_fl_i_13
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [11]),
        .O(ctl_fetch1_fl_i_13_n_0));
  LUT6 #(
    .INIT(64'h00000000FEF00000)) 
    ctl_fetch1_fl_i_14
       (.I0(\rgf/sreg/sr [10]),
        .I1(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [14]),
        .I5(ctl_fetch1_fl_i_23_n_0),
        .O(ctl_fetch1_fl_i_14_n_0));
  LUT5 #(
    .INIT(32'h7F738F83)) 
    ctl_fetch1_fl_i_15
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\rgf/sreg/sr [5]),
        .O(ctl_fetch1_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'h000A2222A0AA2222)) 
    ctl_fetch1_fl_i_16
       (.I0(\fch/ir1 [13]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir1 [14]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir1 [12]),
        .I5(\rgf_selc1_wb[1]_i_29_n_0 ),
        .O(ctl_fetch1_fl_i_16_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch1_fl_i_17
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [5]),
        .O(ctl_fetch1_fl_i_17_n_0));
  LUT6 #(
    .INIT(64'h01000000FFFFFFFF)) 
    ctl_fetch1_fl_i_18
       (.I0(ctl_fetch1_fl_i_24_n_0),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(ctl_fetch1_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF10)) 
    ctl_fetch1_fl_i_19
       (.I0(\bcmd[0]_INST_0_i_24_n_0 ),
        .I1(ctl_fetch1_fl_i_25_n_0),
        .I2(ctl_fetch1_fl_i_26_n_0),
        .I3(ctl_fetch1_fl_i_27_n_0),
        .I4(ctl_fetch1_fl_i_28_n_0),
        .I5(ctl_fetch1_fl_i_29_n_0),
        .O(ctl_fetch1_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'h00000000AAAAFFAE)) 
    ctl_fetch1_fl_i_2
       (.I0(ctl_fetch1_fl_i_6_n_0),
        .I1(ctl_fetch1_fl_i_7_n_0),
        .I2(ctl_fetch1_fl_i_8_n_0),
        .I3(\fch/ir1 [9]),
        .I4(ctl_fetch1_fl_i_9_n_0),
        .I5(ctl_fetch1_fl_i_10_n_0),
        .O(ctl_fetch1_fl_i_2_n_0));
  LUT6 #(
    .INIT(64'hAAAAFFFFFFEAFFEA)) 
    ctl_fetch1_fl_i_20
       (.I0(\ctl1/stat [1]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .I3(\ctl1/stat [0]),
        .I4(ctl_fetch1_fl_i_30_n_0),
        .I5(\fch/ir1 [10]),
        .O(ctl_fetch1_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000808BB0BB)) 
    ctl_fetch1_fl_i_21
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\ctl1/stat [0]),
        .I3(\ctl1/stat [1]),
        .I4(\fch/ir1 [12]),
        .I5(ctl_fetch1_fl_i_31_n_0),
        .O(ctl_fetch1_fl_i_21_n_0));
  LUT6 #(
    .INIT(64'h111F0000111F111F)) 
    ctl_fetch1_fl_i_22
       (.I0(\bcmd[2]_INST_0_i_4_n_0 ),
        .I1(ctl_fetch1_fl_i_32_n_0),
        .I2(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I3(ctl_fetch1_fl_i_33_n_0),
        .I4(ctl_fetch1_fl_i_34_n_0),
        .I5(ctl_fetch1_fl_i_35_n_0),
        .O(ctl_fetch1_fl_i_22_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    ctl_fetch1_fl_i_23
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [10]),
        .O(ctl_fetch1_fl_i_23_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch1_fl_i_24
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .O(ctl_fetch1_fl_i_24_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch1_fl_i_25
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .O(ctl_fetch1_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hF7FFF7FFFFFFFF75)) 
    ctl_fetch1_fl_i_26
       (.I0(\badr[15]_INST_0_i_302_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [5]),
        .O(ctl_fetch1_fl_i_26_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF11F50000)) 
    ctl_fetch1_fl_i_27
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [10]),
        .I4(\bcmd[1]_INST_0_i_8_n_0 ),
        .I5(ctl_fetch1_fl_i_36_n_0),
        .O(ctl_fetch1_fl_i_27_n_0));
  LUT6 #(
    .INIT(64'h44F400F0FFFF00F0)) 
    ctl_fetch1_fl_i_28
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(ctl_fetch1_fl_i_37_n_0),
        .I3(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I4(\ctl1/stat [0]),
        .I5(\rgf_selc1_wb[0]_i_20_n_0 ),
        .O(ctl_fetch1_fl_i_28_n_0));
  LUT6 #(
    .INIT(64'h5D5D5D5DFFFFFF55)) 
    ctl_fetch1_fl_i_29
       (.I0(\stat[2]_i_5__0_n_0 ),
        .I1(\stat[0]_i_34_n_0 ),
        .I2(\rgf/sreg/sr [4]),
        .I3(ctl_fetch1_fl_i_38_n_0),
        .I4(ctl_fetch1_fl_i_39_n_0),
        .I5(\fch/ir1 [12]),
        .O(ctl_fetch1_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    ctl_fetch1_fl_i_3
       (.I0(\bcmd[2]_INST_0_i_4_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [11]),
        .I4(ctl_fetch1_fl_i_11_n_0),
        .I5(ctl_fetch1_fl_i_12_n_0),
        .O(ctl_fetch1_fl_i_3_n_0));
  LUT6 #(
    .INIT(64'hBB00B000BBF0B0FF)) 
    ctl_fetch1_fl_i_30
       (.I0(\rgf/sreg/sr [10]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .I4(\rgf/sreg/sr [11]),
        .I5(\fch/ir1 [9]),
        .O(ctl_fetch1_fl_i_30_n_0));
  LUT3 #(
    .INIT(8'hDC)) 
    ctl_fetch1_fl_i_31
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [10]),
        .O(ctl_fetch1_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'h0002000300020000)) 
    ctl_fetch1_fl_i_32
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [15]),
        .I3(\ctl1/stat [2]),
        .I4(\ctl1/stat [1]),
        .I5(\bcmd[0]_INST_0_i_24_n_0 ),
        .O(ctl_fetch1_fl_i_32_n_0));
  LUT6 #(
    .INIT(64'hFF020000FF02FF02)) 
    ctl_fetch1_fl_i_33
       (.I0(\fadr[15]_INST_0_i_21_n_0 ),
        .I1(ctl_fetch1_fl_i_40_n_0),
        .I2(\ctl1/stat [1]),
        .I3(\bcmd[0]_INST_0_i_24_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_20_n_0 ),
        .I5(\ctl1/stat [0]),
        .O(ctl_fetch1_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFEEEEEE)) 
    ctl_fetch1_fl_i_34
       (.I0(ctl_fetch1_fl_i_41_n_0),
        .I1(\bcmd[0]_INST_0_i_7_n_0 ),
        .I2(\stat[1]_i_18__0_n_0 ),
        .I3(\ctl1/stat [0]),
        .I4(\ctl1/stat [1]),
        .I5(ctl_fetch1_fl_i_42_n_0),
        .O(ctl_fetch1_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'h0000000000FC37D4)) 
    ctl_fetch1_fl_i_35
       (.I0(\ctl1/stat [1]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [3]),
        .I5(ctl_fetch1_fl_i_43_n_0),
        .O(ctl_fetch1_fl_i_35_n_0));
  LUT6 #(
    .INIT(64'h00000000F20000F2)) 
    ctl_fetch1_fl_i_36
       (.I0(\rgf/sreg/sr [4]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\rgf/sreg/sr [5]),
        .I5(\fch/ir1 [13]),
        .O(ctl_fetch1_fl_i_36_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch1_fl_i_37
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir1 [14]),
        .O(ctl_fetch1_fl_i_37_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_38
       (.I0(\fch/ir1 [13]),
        .I1(\rgf/sreg/sr [6]),
        .O(ctl_fetch1_fl_i_38_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_39
       (.I0(\fch/ir1 [14]),
        .I1(\rgf/sreg/sr [5]),
        .O(ctl_fetch1_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'hAFFBAFFBFFFFAFFB)) 
    ctl_fetch1_fl_i_4
       (.I0(ctl_fetch1_fl_i_13_n_0),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\fch/ir1 [6]),
        .O(ctl_fetch1_fl_i_4_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_40
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .O(ctl_fetch1_fl_i_40_n_0));
  LUT6 #(
    .INIT(64'hBABBBAAAB888B888)) 
    ctl_fetch1_fl_i_41
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [3]),
        .I3(\rgf/sreg/sr [10]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [1]),
        .O(ctl_fetch1_fl_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFF8FFFFFFFF)) 
    ctl_fetch1_fl_i_42
       (.I0(\ctl1/stat [2]),
        .I1(\fch/ir1 [2]),
        .I2(\bdatw[11]_INST_0_i_27_n_0 ),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [15]),
        .I5(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .O(ctl_fetch1_fl_i_42_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    ctl_fetch1_fl_i_43
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [13]),
        .O(ctl_fetch1_fl_i_43_n_0));
  LUT6 #(
    .INIT(64'hDD55D040DD55DD55)) 
    ctl_fetch1_fl_i_5
       (.I0(\bcmd[2]_INST_0_i_4_n_0 ),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [1]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [6]),
        .I5(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .O(ctl_fetch1_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBAAABBBBB)) 
    ctl_fetch1_fl_i_6
       (.I0(\fch/ir1 [11]),
        .I1(ctl_fetch1_fl_i_14_n_0),
        .I2(ctl_fetch1_fl_i_15_n_0),
        .I3(\fch/ir1 [13]),
        .I4(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I5(ctl_fetch1_fl_i_16_n_0),
        .O(ctl_fetch1_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFFF0FFFFF10FF10)) 
    ctl_fetch1_fl_i_7
       (.I0(\fch/ir1 [3]),
        .I1(ctl_fetch0_fl_i_13_n_0),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [2]),
        .I4(\rgf/sreg/sr [10]),
        .I5(\fch/ir1 [1]),
        .O(ctl_fetch1_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFF0FFF8FFF0)) 
    ctl_fetch1_fl_i_8
       (.I0(\rgf/sreg/sr [10]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [4]),
        .I3(ctl_fetch1_fl_i_17_n_0),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [1]),
        .O(ctl_fetch1_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hFF5FFFFFFFFFFF51)) 
    ctl_fetch1_fl_i_9
       (.I0(\rgf_selc1_wb[1]_i_20_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [9]),
        .O(ctl_fetch1_fl_i_9_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_ext_fl_i_1
       (.I0(\fadr[15]_INST_0_i_4_n_0 ),
        .O(ctl_fetch_ext_fl_i_1_n_0));
  LUT3 #(
    .INIT(8'hFB)) 
    \eir_fl[15]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .O(\eir_fl[15]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(irq_vec[0]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(\fch/eir [1]),
        .O(\eir_fl[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(irq_vec[1]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(\fch/eir [2]),
        .O(\eir_fl[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(irq_vec[2]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(\fch/eir [3]),
        .O(\eir_fl[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(irq_vec[3]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(\fch/eir [4]),
        .O(\eir_fl[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(irq_vec[4]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(\fch/eir [5]),
        .O(\eir_fl[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \eir_fl[6]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .O(\eir_fl[6]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_2 
       (.I0(irq_vec[5]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(\fch/eir [6]),
        .O(\eir_fl[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_1
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [15]),
        .I2(eir_inferred_i_17_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[15] ),
        .O(\fch/eir [15]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_10
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [6]),
        .I2(eir_inferred_i_26_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[6] ),
        .O(\fch/eir [6]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_11
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [5]),
        .I2(eir_inferred_i_27_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[5] ),
        .O(\fch/eir [5]));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_12
       (.I0(\fch/rst_n_fl ),
        .I1(eir_inferred_i_28_n_0),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/fch_leir_nir ),
        .I4(\fch/nir [4]),
        .I5(\fch/eir_fl_reg_n_0_[4] ),
        .O(\fch/eir [4]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_13
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [3]),
        .I2(eir_inferred_i_29_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[3] ),
        .O(\fch/eir [3]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_14
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [2]),
        .I2(eir_inferred_i_30_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[2] ),
        .O(\fch/eir [2]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_15
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [1]),
        .I2(eir_inferred_i_31_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[1] ),
        .O(\fch/eir [1]));
  LUT6 #(
    .INIT(64'hB800FF00B8000000)) 
    eir_inferred_i_16
       (.I0(\fch/nir [0]),
        .I1(\fch/fch_leir_nir ),
        .I2(eir_inferred_i_32_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[0] ),
        .O(\fch/eir [0]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_17
       (.I0(fdat[15]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[15] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[15]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_18
       (.I0(fdat[14]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[14] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[14]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_19
       (.I0(fdat[13]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[13] ),
        .I3(fdatx[13]),
        .I4(\fch/fch_leir_hir ),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_2
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [14]),
        .I2(eir_inferred_i_18_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[14] ),
        .O(\fch/eir [14]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_20
       (.I0(fdat[12]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[12] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[12]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_21
       (.I0(fdat[11]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[11] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[11]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_22
       (.I0(fdat[10]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[10] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[10]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_23
       (.I0(fdat[9]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[9] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[9]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_24
       (.I0(fdat[8]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[8] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[8]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_25
       (.I0(fdat[7]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[7] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[7]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_26
       (.I0(fdat[6]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[6] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[6]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_27
       (.I0(fdat[5]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[5] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[5]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00B8B8)) 
    eir_inferred_i_28
       (.I0(fdat[4]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[4] ),
        .I3(fdatx[4]),
        .I4(\fch/fch_leir_hir ),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_29
       (.I0(fdat[3]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[3] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[3]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h8A8A0A8A80800080)) 
    eir_inferred_i_3
       (.I0(\fch/rst_n_fl ),
        .I1(eir_inferred_i_19_n_0),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/fch_leir_nir ),
        .I4(\fch/nir [13]),
        .I5(\fch/eir_fl_reg_n_0_[13] ),
        .O(\fch/eir [13]));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_30
       (.I0(fdat[2]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[2] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[2]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h00000000FFB800B8)) 
    eir_inferred_i_31
       (.I0(fdat[1]),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/eir_fl_reg_n_0_[1] ),
        .I3(\fch/fch_leir_hir ),
        .I4(fdatx[1]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_31_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    eir_inferred_i_32
       (.I0(fdatx[0]),
        .I1(\fch/fch_leir_hir ),
        .I2(fdat[0]),
        .I3(\fch/fch_leir_lir ),
        .I4(\fch/eir_fl_reg_n_0_[0] ),
        .O(eir_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_4
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [12]),
        .I2(eir_inferred_i_20_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[12] ),
        .O(\fch/eir [12]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_5
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [11]),
        .I2(eir_inferred_i_21_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[11] ),
        .O(\fch/eir [11]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_6
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [10]),
        .I2(eir_inferred_i_22_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[10] ),
        .O(\fch/eir [10]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_7
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [9]),
        .I2(eir_inferred_i_23_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[9] ),
        .O(\fch/eir [9]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_8
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [8]),
        .I2(eir_inferred_i_24_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[8] ),
        .O(\fch/eir [8]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_9
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/nir [7]),
        .I2(eir_inferred_i_25_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(\fch/eir_fl_reg_n_0_[7] ),
        .O(\fch/eir [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \fadr[0]_INST_0 
       (.I0(\fch/p_2_in [0]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/pcnt/pc [0]),
        .O(fadr[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[10]_INST_0 
       (.I0(\fch/p_2_in [10]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__1_n_6 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [10]),
        .O(fadr[10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[11]_INST_0 
       (.I0(\fch/p_2_in [11]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__1_n_5 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [11]),
        .O(fadr[11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[12]_INST_0 
       (.I0(\fch/p_2_in [12]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__1_n_4 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [12]),
        .O(fadr[12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[13]_INST_0 
       (.I0(\fch/p_2_in [13]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__2_n_7 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [13]),
        .O(fadr[13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[14]_INST_0 
       (.I0(\fch/p_2_in [14]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__2_n_6 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [14]),
        .O(fadr[14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[15]_INST_0 
       (.I0(\fch/p_2_in [15]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__2_n_5 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [15]),
        .O(fadr[15]));
  LUT5 #(
    .INIT(32'h00000070)) 
    \fadr[15]_INST_0_i_1 
       (.I0(\fadr[15]_INST_0_i_3_n_0 ),
        .I1(\fadr[15]_INST_0_i_4_n_0 ),
        .I2(\fadr[15]_INST_0_i_5_n_0 ),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .O(\fadr[15]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \fadr[15]_INST_0_i_10 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [0]),
        .O(\fadr[15]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \fadr[15]_INST_0_i_11 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [11]),
        .O(\fadr[15]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \fadr[15]_INST_0_i_12 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\ccmd[4]_INST_0_i_8_n_0 ),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [4]),
        .I5(\ccmd[2]_INST_0_i_5_n_0 ),
        .O(\fadr[15]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \fadr[15]_INST_0_i_13 
       (.I0(\fadr[15]_INST_0_i_17_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I2(\fadr[15]_INST_0_i_18_n_0 ),
        .I3(\fch/ir1 [15]),
        .I4(\fadr[15]_INST_0_i_19_n_0 ),
        .I5(\fadr[15]_INST_0_i_20_n_0 ),
        .O(ctl_fetch_ext1));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \fadr[15]_INST_0_i_14 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [3]),
        .O(\fadr[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \fadr[15]_INST_0_i_15 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(\ccmd[2]_INST_0_i_5_n_0 ),
        .I5(\ccmd[2]_INST_0_i_4_n_0 ),
        .O(\fadr[15]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \fadr[15]_INST_0_i_16 
       (.I0(\ctl1/stat [0]),
        .I1(\ctl1/stat [1]),
        .I2(\ctl1/stat [2]),
        .O(ctl_bcc_take1));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \fadr[15]_INST_0_i_17 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\badr[15]_INST_0_i_144_n_0 ),
        .I5(\fadr[15]_INST_0_i_21_n_0 ),
        .O(\fadr[15]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \fadr[15]_INST_0_i_18 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [1]),
        .O(\fadr[15]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \fadr[15]_INST_0_i_19 
       (.I0(\fch/ir1 [2]),
        .I1(\ctl1/stat [2]),
        .O(\fadr[15]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A000000000000)) 
    \fadr[15]_INST_0_i_2 
       (.I0(\fadr[15]_INST_0_i_6_n_0 ),
        .I1(\fch/stat [2]),
        .I2(\fch/stat [0]),
        .I3(\fadr[15]_INST_0_i_7_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fch/stat [1]),
        .O(\fadr[15]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_20 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [3]),
        .O(\fadr[15]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \fadr[15]_INST_0_i_21 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .O(\fadr[15]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \fadr[15]_INST_0_i_3 
       (.I0(\fadr[15]_INST_0_i_8_n_0 ),
        .I1(fch_term),
        .O(\fadr[15]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFDFFFFF)) 
    \fadr[15]_INST_0_i_4 
       (.I0(\fadr[15]_INST_0_i_9_n_0 ),
        .I1(\fadr[15]_INST_0_i_10_n_0 ),
        .I2(\ctl0/stat [2]),
        .I3(\fadr[15]_INST_0_i_11_n_0 ),
        .I4(\fadr[15]_INST_0_i_12_n_0 ),
        .I5(ctl_fetch_ext1),
        .O(\fadr[15]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAAAA8)) 
    \fadr[15]_INST_0_i_5 
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir0 [15]),
        .I2(\fadr[15]_INST_0_i_4_n_0 ),
        .I3(\fadr[15]_INST_0_i_14_n_0 ),
        .I4(\fadr[15]_INST_0_i_15_n_0 ),
        .O(\fadr[15]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00E2)) 
    \fadr[15]_INST_0_i_6 
       (.I0(\fch/fch_issu1_fl ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_issu1 ),
        .I3(\fch/stat [2]),
        .I4(\fch/stat [0]),
        .I5(\fadr[15]_INST_0_i_3_n_0 ),
        .O(\fadr[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004540)) 
    \fadr[15]_INST_0_i_7 
       (.I0(\fch/stat [2]),
        .I1(\fch/fch_issu1 ),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_issu1_fl ),
        .I4(\fadr[15]_INST_0_i_4_n_0 ),
        .I5(\fch/stat [0]),
        .O(\fadr[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF80)) 
    \fadr[15]_INST_0_i_8 
       (.I0(\ctl0/stat [1]),
        .I1(\ctl0/stat [0]),
        .I2(\ctl0/stat [2]),
        .I3(\fch/ctl_bcc_take1_fl ),
        .I4(\fch/ctl_bcc_take0_fl ),
        .I5(ctl_bcc_take1),
        .O(\fadr[15]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fadr[15]_INST_0_i_9 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [13]),
        .O(\fadr[15]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[1]_INST_0 
       (.I0(\fch/p_2_in [1]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry_n_7 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [1]),
        .O(fadr[1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[2]_INST_0 
       (.I0(\fch/p_2_in [2]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry_n_6 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [2]),
        .O(fadr[2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[3]_INST_0 
       (.I0(\fch/p_2_in [3]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry_n_5 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [3]),
        .O(fadr[3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[4]_INST_0 
       (.I0(\fch/p_2_in [4]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry_n_4 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [4]),
        .O(fadr[4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[5]_INST_0 
       (.I0(\fch/p_2_in [5]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__0_n_7 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [5]),
        .O(fadr[5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[6]_INST_0 
       (.I0(\fch/p_2_in [6]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__0_n_6 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [6]),
        .O(fadr[6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[7]_INST_0 
       (.I0(\fch/p_2_in [7]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__0_n_5 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [7]),
        .O(fadr[7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[8]_INST_0 
       (.I0(\fch/p_2_in [8]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__0_n_4 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [8]),
        .O(fadr[8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[9]_INST_0 
       (.I0(\fch/p_2_in [9]),
        .I1(\fadr[15]_INST_0_i_1_n_0 ),
        .I2(\fch/fch_pc_nx4_carry__1_n_7 ),
        .I3(\fadr[15]_INST_0_i_2_n_0 ),
        .I4(\rgf/pcnt/pc [9]),
        .O(fadr[9]));
  FDRE \fch/ctl_bcc_take0_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take0_fl_i_1_n_0),
        .Q(\fch/ctl_bcc_take0_fl ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/ctl_bcc_take1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take1_fl_i_1_n_0),
        .Q(\fch/ctl_bcc_take1_fl ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/ctl_fetch0_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch0),
        .Q(\fch/ctl_fetch0_fl ),
        .R(\<const0> ));
  FDRE \fch/ctl_fetch1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch1),
        .Q(\fch/ctl_fetch1_fl ),
        .R(\<const0> ));
  FDRE \fch/ctl_fetch_ext_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_ext_fl_i_1_n_0),
        .Q(\fch/ctl_fetch_ext_fl ),
        .R(\<const0> ));
  FDRE \fch/eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [0]),
        .Q(\fch/eir_fl_reg_n_0_[0] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [10]),
        .Q(\fch/eir_fl_reg_n_0_[10] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [11]),
        .Q(\fch/eir_fl_reg_n_0_[11] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [12]),
        .Q(\fch/eir_fl_reg_n_0_[12] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [13]),
        .Q(\fch/eir_fl_reg_n_0_[13] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [14]),
        .Q(\fch/eir_fl_reg_n_0_[14] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [15]),
        .Q(\fch/eir_fl_reg_n_0_[15] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[1]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[1] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[2]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[2] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[3]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[3] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[4]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[4] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[5]_i_1_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[5] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[6]_i_2_n_0 ),
        .Q(\fch/eir_fl_reg_n_0_[6] ),
        .R(\eir_fl[6]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [7]),
        .Q(\fch/eir_fl_reg_n_0_[7] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [8]),
        .Q(\fch/eir_fl_reg_n_0_[8] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [9]),
        .Q(\fch/eir_fl_reg_n_0_[9] ),
        .R(\eir_fl[15]_i_1_n_0 ));
  FDRE \fch/fadr_1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fadr[1]),
        .Q(\fch/fadr_1_fl ),
        .R(\<const0> ));
  FDRE \fch/fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[0]_i_1_n_0 ),
        .Q(fch_irq_lev[0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[1]_i_1_n_0 ),
        .Q(fch_irq_lev[1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/fch_irq_req_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(\fch/fch_irq_req_fl ),
        .R(\<const0> ));
  FDRE \fch/fch_issu1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fch_issu1_ir ),
        .Q(\fch/fch_issu1_fl ),
        .R(\<const0> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx2_carry 
       (.CI(\<const0> ),
        .CO({\fch/fch_pc_nx2_carry_n_0 ,\fch/fch_pc_nx2_carry_n_1 ,\fch/fch_pc_nx2_carry_n_2 ,\fch/fch_pc_nx2_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/pcnt/pc [1],\<const0> }),
        .O(\fch/p_2_in [3:0]),
        .S({\rgf/pcnt/pc [3:2],fch_pc_nx2_carry_i_1_n_0,\rgf/pcnt/pc [0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx2_carry__0 
       (.CI(\fch/fch_pc_nx2_carry_n_0 ),
        .CO({\fch/fch_pc_nx2_carry__0_n_0 ,\fch/fch_pc_nx2_carry__0_n_1 ,\fch/fch_pc_nx2_carry__0_n_2 ,\fch/fch_pc_nx2_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in [7:4]),
        .S(\rgf/pcnt/pc [7:4]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx2_carry__1 
       (.CI(\fch/fch_pc_nx2_carry__0_n_0 ),
        .CO({\fch/fch_pc_nx2_carry__1_n_0 ,\fch/fch_pc_nx2_carry__1_n_1 ,\fch/fch_pc_nx2_carry__1_n_2 ,\fch/fch_pc_nx2_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in [11:8]),
        .S(\rgf/pcnt/pc [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx2_carry__2 
       (.CI(\fch/fch_pc_nx2_carry__1_n_0 ),
        .CO({\fch/fch_pc_nx2_carry__2_n_1 ,\fch/fch_pc_nx2_carry__2_n_2 ,\fch/fch_pc_nx2_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in [15:12]),
        .S(\rgf/pcnt/pc [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx4_carry 
       (.CI(\<const0> ),
        .CO({\fch/fch_pc_nx4_carry_n_0 ,\fch/fch_pc_nx4_carry_n_1 ,\fch/fch_pc_nx4_carry_n_2 ,\fch/fch_pc_nx4_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/pcnt/pc [2],\<const0> }),
        .O({\fch/fch_pc_nx4_carry_n_4 ,\fch/fch_pc_nx4_carry_n_5 ,\fch/fch_pc_nx4_carry_n_6 ,\fch/fch_pc_nx4_carry_n_7 }),
        .S({\rgf/pcnt/pc [4:3],fch_pc_nx4_carry_i_1_n_0,\rgf/pcnt/pc [1]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx4_carry__0 
       (.CI(\fch/fch_pc_nx4_carry_n_0 ),
        .CO({\fch/fch_pc_nx4_carry__0_n_0 ,\fch/fch_pc_nx4_carry__0_n_1 ,\fch/fch_pc_nx4_carry__0_n_2 ,\fch/fch_pc_nx4_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fch/fch_pc_nx4_carry__0_n_4 ,\fch/fch_pc_nx4_carry__0_n_5 ,\fch/fch_pc_nx4_carry__0_n_6 ,\fch/fch_pc_nx4_carry__0_n_7 }),
        .S(\rgf/pcnt/pc [8:5]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx4_carry__1 
       (.CI(\fch/fch_pc_nx4_carry__0_n_0 ),
        .CO({\fch/fch_pc_nx4_carry__1_n_0 ,\fch/fch_pc_nx4_carry__1_n_1 ,\fch/fch_pc_nx4_carry__1_n_2 ,\fch/fch_pc_nx4_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fch/fch_pc_nx4_carry__1_n_4 ,\fch/fch_pc_nx4_carry__1_n_5 ,\fch/fch_pc_nx4_carry__1_n_6 ,\fch/fch_pc_nx4_carry__1_n_7 }),
        .S(\rgf/pcnt/pc [12:9]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/fch_pc_nx4_carry__2 
       (.CI(\fch/fch_pc_nx4_carry__1_n_0 ),
        .CO({\fch/fch_pc_nx4_carry__2_n_2 ,\fch/fch_pc_nx4_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fch/fch_pc_nx4_carry__2_n_5 ,\fch/fch_pc_nx4_carry__2_n_6 ,\fch/fch_pc_nx4_carry__2_n_7 }),
        .S({\<const0> ,\rgf/pcnt/pc [15:13]}));
  FDRE \fch/fch_term_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(\fch/fch_term_fl ),
        .R(\<const0> ));
  FDRE \fch/fctl/fch_leir_hir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_leir_hir_t ),
        .Q(\fch/fch_leir_hir ),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \fch/fctl/fch_leir_lir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_leir_lir_t ),
        .Q(\fch/fch_leir_lir ),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \fch/fctl/fch_leir_nir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_leir_nir_t ),
        .Q(\fch/fch_leir_nir ),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \fch/fctl/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/stat_nx [0]),
        .Q(\fch/stat [0]),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \fch/fctl/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/stat_nx [1]),
        .Q(\fch/stat [1]),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \fch/fctl/stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/stat_nx [2]),
        .Q(\fch/stat [2]),
        .R(\stat[2]_i_1__1_n_0 ));
  FDRE \fch/ir0_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [0]),
        .Q(\fch/ir0_fl [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [10]),
        .Q(\fch/ir0_fl [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [11]),
        .Q(\fch/ir0_fl [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [12]),
        .Q(\fch/ir0_fl [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [13]),
        .Q(\fch/ir0_fl [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [14]),
        .Q(\fch/ir0_fl [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [15]),
        .Q(\fch/ir0_fl [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [1]),
        .Q(\fch/ir0_fl [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [2]),
        .Q(\fch/ir0_fl [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [3]),
        .Q(\fch/ir0_fl [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [4]),
        .Q(\fch/ir0_fl [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [5]),
        .Q(\fch/ir0_fl [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [6]),
        .Q(\fch/ir0_fl [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [7]),
        .Q(\fch/ir0_fl [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [8]),
        .Q(\fch/ir0_fl [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [9]),
        .Q(\fch/ir0_fl [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/p_0_in ),
        .Q(\fch/ir0_id_fl [20]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir0_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0_id ),
        .Q(\fch/ir0_id_fl [21]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [0]),
        .Q(\fch/ir1_fl [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [10]),
        .Q(\fch/ir1_fl [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [11]),
        .Q(\fch/ir1_fl [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [12]),
        .Q(\fch/ir1_fl [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [13]),
        .Q(\fch/ir1_fl [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [14]),
        .Q(\fch/ir1_fl [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [15]),
        .Q(\fch/ir1_fl [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [1]),
        .Q(\fch/ir1_fl [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [2]),
        .Q(\fch/ir1_fl [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [3]),
        .Q(\fch/ir1_fl [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [4]),
        .Q(\fch/ir1_fl [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [5]),
        .Q(\fch/ir1_fl [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [6]),
        .Q(\fch/ir1_fl [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [7]),
        .Q(\fch/ir1_fl [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [8]),
        .Q(\fch/ir1_fl [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [9]),
        .Q(\fch/ir1_fl [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_wrbufn1),
        .Q(\fch/ir1_id_fl [20]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/ir1_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_memacc1),
        .Q(\fch/ir1_id_fl [21]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[12] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [12]),
        .Q(\fch/nir_id [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[13] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [13]),
        .Q(\fch/nir_id [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[14] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [14]),
        .Q(\fch/nir_id [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[15] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [15]),
        .Q(\fch/nir_id [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[16] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [16]),
        .Q(\fch/nir_id [16]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[17] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [17]),
        .Q(\fch/nir_id [17]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[18] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [18]),
        .Q(\fch/nir_id [18]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[19] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [19]),
        .Q(\fch/nir_id [19]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[20] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\nir_id[20]_i_1_n_0 ),
        .Q(\fch/nir_id [20]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[21] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [21]),
        .Q(\fch/nir_id [21]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_id_reg[24] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [24]),
        .Q(\fch/nir_id [24]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[0] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[0]),
        .Q(\fch/nir [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[10] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[10]),
        .Q(\fch/nir [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[11] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[11]),
        .Q(\fch/nir [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[12] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[12]),
        .Q(\fch/nir [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[13] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[13]),
        .Q(\fch/nir [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[14] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[14]),
        .Q(\fch/nir [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[15] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[15]),
        .Q(\fch/nir [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[1] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[1]),
        .Q(\fch/nir [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[2] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[2]),
        .Q(\fch/nir [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[3] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[3]),
        .Q(\fch/nir [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[4] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[4]),
        .Q(\fch/nir [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[5] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[5]),
        .Q(\fch/nir [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[6] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[6]),
        .Q(\fch/nir [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[7] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[7]),
        .Q(\fch/nir [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[8] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[8]),
        .Q(\fch/nir [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/nir_reg[9] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[9]),
        .Q(\fch/nir [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[0]),
        .Q(fch_pc0[0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[10]),
        .Q(fch_pc0[10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[11]),
        .Q(fch_pc0[11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[12]),
        .Q(fch_pc0[12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[13]),
        .Q(fch_pc0[13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[14]),
        .Q(fch_pc0[14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[15]),
        .Q(fch_pc0[15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[1]),
        .Q(fch_pc0[1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[2]),
        .Q(fch_pc0[2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[3]),
        .Q(fch_pc0[3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[4]),
        .Q(fch_pc0[4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[5]),
        .Q(fch_pc0[5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[6]),
        .Q(fch_pc0[6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[7]),
        .Q(fch_pc0[7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[8]),
        .Q(fch_pc0[8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc0_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[9]),
        .Q(fch_pc0[9]),
        .R(\rgf/treg/p_0_in ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/pc10_carry 
       (.CI(\<const0> ),
        .CO({\fch/pc10_carry_n_0 ,\fch/pc10_carry_n_1 ,\fch/pc10_carry_n_2 ,\fch/pc10_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,fch_pc[1],\<const0> }),
        .O({\fch/pc10_carry_n_4 ,\fch/pc10_carry_n_5 ,\fch/pc10_carry_n_6 ,\fch/pc10_carry_n_7 }),
        .S({pc10_carry_i_1_n_0,pc10_carry_i_2_n_0,pc10_carry_i_3_n_0,pc10_carry_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/pc10_carry__0 
       (.CI(\fch/pc10_carry_n_0 ),
        .CO({\fch/pc10_carry__0_n_0 ,\fch/pc10_carry__0_n_1 ,\fch/pc10_carry__0_n_2 ,\fch/pc10_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fch/pc10_carry__0_n_4 ,\fch/pc10_carry__0_n_5 ,\fch/pc10_carry__0_n_6 ,\fch/pc10_carry__0_n_7 }),
        .S({pc10_carry__0_i_1_n_0,pc10_carry__0_i_2_n_0,pc10_carry__0_i_3_n_0,pc10_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/pc10_carry__1 
       (.CI(\fch/pc10_carry__0_n_0 ),
        .CO({\fch/pc10_carry__1_n_0 ,\fch/pc10_carry__1_n_1 ,\fch/pc10_carry__1_n_2 ,\fch/pc10_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fch/pc10_carry__1_n_4 ,\fch/pc10_carry__1_n_5 ,\fch/pc10_carry__1_n_6 ,\fch/pc10_carry__1_n_7 }),
        .S({pc10_carry__1_i_1_n_0,pc10_carry__1_i_2_n_0,pc10_carry__1_i_3_n_0,pc10_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fch/pc10_carry__2 
       (.CI(\fch/pc10_carry__1_n_0 ),
        .CO({\fch/pc10_carry__2_n_1 ,\fch/pc10_carry__2_n_2 ,\fch/pc10_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fch/pc10_carry__2_n_4 ,\fch/pc10_carry__2_n_5 ,\fch/pc10_carry__2_n_6 ,\fch/pc10_carry__2_n_7 }),
        .S({pc10_carry__2_i_1_n_0,pc10_carry__2_i_2_n_0,pc10_carry__2_i_3_n_0,pc10_carry__2_i_4_n_0}));
  FDRE \fch/pc1_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry_n_7 ),
        .Q(fch_pc1[0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__1_n_5 ),
        .Q(fch_pc1[10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__1_n_4 ),
        .Q(fch_pc1[11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__2_n_7 ),
        .Q(fch_pc1[12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__2_n_6 ),
        .Q(fch_pc1[13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__2_n_5 ),
        .Q(fch_pc1[14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__2_n_4 ),
        .Q(fch_pc1[15]),
        .R(\rgf/treg/p_0_in ));
  FDSE \fch/pc1_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry_n_6 ),
        .Q(fch_pc1[1]),
        .S(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry_n_5 ),
        .Q(fch_pc1[2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry_n_4 ),
        .Q(fch_pc1[3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__0_n_7 ),
        .Q(fch_pc1[4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__0_n_6 ),
        .Q(fch_pc1[5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__0_n_5 ),
        .Q(fch_pc1[6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__0_n_4 ),
        .Q(fch_pc1[7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__1_n_7 ),
        .Q(fch_pc1[8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/pc1_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(\fch/pc10_carry__1_n_6 ),
        .Q(fch_pc1[9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \fch/rst_n_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(\fch/rst_n_fl ),
        .R(\<const0> ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(fch_irq_lev[0]),
        .O(\fch_irq_lev[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(fch_irq_lev[1]),
        .O(\fch_irq_lev[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h5555004000400040)) 
    \fch_irq_lev[1]_i_2 
       (.I0(\pc0[15]_i_3_n_0 ),
        .I1(\fadr[15]_INST_0_i_12_n_0 ),
        .I2(\bdatw[8]_INST_0_i_15_n_0 ),
        .I3(\sr[13]_i_8_n_0 ),
        .I4(\stat[0]_i_7__0_n_0 ),
        .I5(\fch_irq_lev[1]_i_3_n_0 ),
        .O(\fch_irq_lev[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \fch_irq_lev[1]_i_3 
       (.I0(\fadr[15]_INST_0_i_17_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [1]),
        .I4(\ctl1/stat [2]),
        .I5(\fch_irq_lev[1]_i_5_n_0 ),
        .O(\fch_irq_lev[1]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \fch_irq_lev[1]_i_4 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [0]),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \fch_irq_lev[1]_i_5 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [14]),
        .O(\fch_irq_lev[1]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h2000AA20)) 
    fch_irq_req_fl_i_1
       (.I0(irq),
        .I1(irq_lev[0]),
        .I2(\rgf/sreg/sr [2]),
        .I3(\rgf/sreg/sr [3]),
        .I4(irq_lev[1]),
        .O(fch_irq_req));
  LUT3 #(
    .INIT(8'hB8)) 
    fch_issu1_fl_i_1
       (.I0(\fch/fch_issu1 ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_issu1_fl ),
        .O(\fch/fch_issu1_ir ));
  LUT6 #(
    .INIT(64'h0000000054450000)) 
    fch_issu1_inferred_i_1
       (.I0(fch_issu1_inferred_i_2_n_0),
        .I1(fch_issu1_inferred_i_3_n_0),
        .I2(fch_issu1_inferred_i_4_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_6_n_0),
        .I5(fch_issu1_inferred_i_7_n_0),
        .O(\fch/fch_issu1 ));
  LUT6 #(
    .INIT(64'hEEF0EEEEEEFFEEEE)) 
    fch_issu1_inferred_i_10
       (.I0(fdat[1]),
        .I1(fch_issu1_inferred_i_36_n_0),
        .I2(fdatx[1]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fch_issu1_inferred_i_37_n_0),
        .O(fch_issu1_inferred_i_10_n_0));
  LUT6 #(
    .INIT(64'h0414545455555555)) 
    fch_issu1_inferred_i_100
       (.I0(fdatx[11]),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[6]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_100_n_0));
  LUT6 #(
    .INIT(64'h0004400004004400)) 
    fch_issu1_inferred_i_101
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_101_n_0));
  LUT6 #(
    .INIT(64'hFEFF5455FFFFFFFF)) 
    fch_issu1_inferred_i_102
       (.I0(fdatx[9]),
        .I1(fdatx[8]),
        .I2(fdatx[6]),
        .I3(fdatx[7]),
        .I4(fch_issu1_inferred_i_166_n_0),
        .I5(fch_issu1_inferred_i_119_n_0),
        .O(fch_issu1_inferred_i_102_n_0));
  LUT6 #(
    .INIT(64'h000000005777FFFF)) 
    fch_issu1_inferred_i_103
       (.I0(fch_issu1_inferred_i_167_n_0),
        .I1(fch_issu1_inferred_i_168_n_0),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_127_n_0),
        .O(fch_issu1_inferred_i_103_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_104
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .O(fch_issu1_inferred_i_104_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_105
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_105_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    fch_issu1_inferred_i_106
       (.I0(fch_issu1_inferred_i_169_n_0),
        .I1(fch_issu1_inferred_i_170_n_0),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[13]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_106_n_0));
  LUT3 #(
    .INIT(8'h45)) 
    fch_issu1_inferred_i_107
       (.I0(\fch/fadr_1_fl ),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [1]),
        .O(fch_issu1_inferred_i_107_n_0));
  LUT6 #(
    .INIT(64'h0DFDFDFDFDFDFDFD)) 
    fch_issu1_inferred_i_108
       (.I0(fdatx[3]),
        .I1(fch_issu1_inferred_i_165_n_0),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[0]),
        .I5(fch_issu1_inferred_i_171_n_0),
        .O(fch_issu1_inferred_i_108_n_0));
  LUT4 #(
    .INIT(16'hCFA7)) 
    fch_issu1_inferred_i_109
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .O(fch_issu1_inferred_i_109_n_0));
  LUT6 #(
    .INIT(64'h10111F1110111011)) 
    fch_issu1_inferred_i_11
       (.I0(fch_issu1_inferred_i_36_n_0),
        .I1(fdat[2]),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_37_n_0),
        .O(fch_issu1_inferred_i_11_n_0));
  LUT4 #(
    .INIT(16'hFF5D)) 
    fch_issu1_inferred_i_110
       (.I0(fdat[8]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_110_n_0));
  LUT4 #(
    .INIT(16'h8088)) 
    fch_issu1_inferred_i_111
       (.I0(fdat[13]),
        .I1(fdat[12]),
        .I2(fdat[14]),
        .I3(fdat[11]),
        .O(fch_issu1_inferred_i_111_n_0));
  LUT6 #(
    .INIT(64'h0DFDFDFDFDFDFDFD)) 
    fch_issu1_inferred_i_112
       (.I0(fdat[3]),
        .I1(\nir_id[14]_i_12_n_0 ),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[0]),
        .I5(fch_issu1_inferred_i_172_n_0),
        .O(fch_issu1_inferred_i_112_n_0));
  LUT6 #(
    .INIT(64'h0454145455555555)) 
    fch_issu1_inferred_i_113
       (.I0(fdat[11]),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(fdat[6]),
        .I4(fdat[7]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_113_n_0));
  LUT4 #(
    .INIT(16'hF93B)) 
    fch_issu1_inferred_i_114
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fdat[6]),
        .O(fch_issu1_inferred_i_114_n_0));
  LUT6 #(
    .INIT(64'hFF0FFFFFFF020000)) 
    fch_issu1_inferred_i_115
       (.I0(fch_issu1_inferred_i_84_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_173_n_0),
        .I4(fch_issu1_inferred_i_119_n_0),
        .I5(fdatx[3]),
        .O(fch_issu1_inferred_i_115_n_0));
  LUT6 #(
    .INIT(64'h00000000CFCFCFEF)) 
    fch_issu1_inferred_i_116
       (.I0(fch_issu1_inferred_i_159_n_0),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .I3(fdatx[3]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_174_n_0),
        .O(fch_issu1_inferred_i_116_n_0));
  LUT4 #(
    .INIT(16'h0100)) 
    fch_issu1_inferred_i_117
       (.I0(fdatx[9]),
        .I1(fdatx[8]),
        .I2(fdatx[6]),
        .I3(fdatx[7]),
        .O(fch_issu1_inferred_i_117_n_0));
  LUT4 #(
    .INIT(16'hEFFF)) 
    fch_issu1_inferred_i_118
       (.I0(fch_issu1_inferred_i_101_n_0),
        .I1(fch_issu1_inferred_i_100_n_0),
        .I2(fdatx[12]),
        .I3(fdatx[13]),
        .O(fch_issu1_inferred_i_118_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_119
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_119_n_0));
  LUT6 #(
    .INIT(64'hEFFFEFEEEFFFEFFF)) 
    fch_issu1_inferred_i_12
       (.I0(fch_issu1_inferred_i_38_n_0),
        .I1(\rgf/sreg/sr [9]),
        .I2(fch_issu1_inferred_i_39_n_0),
        .I3(fch_issu1_inferred_i_20_n_0),
        .I4(fch_issu1_inferred_i_40_n_0),
        .I5(fch_issu1_inferred_i_41_n_0),
        .O(fch_issu1_inferred_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    fch_issu1_inferred_i_120
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .I4(fdatx[8]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_120_n_0));
  LUT4 #(
    .INIT(16'hEFFF)) 
    fch_issu1_inferred_i_121
       (.I0(fdatx[13]),
        .I1(fdatx[12]),
        .I2(fdatx[1]),
        .I3(fdatx[0]),
        .O(fch_issu1_inferred_i_121_n_0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    fch_issu1_inferred_i_122
       (.I0(fdatx[2]),
        .I1(fdatx[3]),
        .I2(fdatx[4]),
        .I3(fdatx[5]),
        .O(fch_issu1_inferred_i_122_n_0));
  LUT4 #(
    .INIT(16'h0001)) 
    fch_issu1_inferred_i_123
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .O(fch_issu1_inferred_i_123_n_0));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    fch_issu1_inferred_i_124
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fch_issu1_inferred_i_175_n_0),
        .I3(fdat[0]),
        .I4(fdat[9]),
        .I5(\nir_id[24]_i_12_n_0 ),
        .O(fch_issu1_inferred_i_124_n_0));
  LUT6 #(
    .INIT(64'hFFF3FFFBFF33FFFB)) 
    fch_issu1_inferred_i_125
       (.I0(fdat[4]),
        .I1(fdat[8]),
        .I2(fdat[5]),
        .I3(fdat[2]),
        .I4(fdat[6]),
        .I5(fdat[3]),
        .O(fch_issu1_inferred_i_125_n_0));
  LUT6 #(
    .INIT(64'h40FF40FF40FFFFFF)) 
    fch_issu1_inferred_i_126
       (.I0(fch_issu1_inferred_i_176_n_0),
        .I1(fch_issu1_inferred_i_177_n_0),
        .I2(fch_issu1_inferred_i_178_n_0),
        .I3(fdatx[9]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_168_n_0),
        .O(fch_issu1_inferred_i_126_n_0));
  LUT4 #(
    .INIT(16'h1000)) 
    fch_issu1_inferred_i_127
       (.I0(fdatx[9]),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .O(fch_issu1_inferred_i_127_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_128
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_128_n_0));
  LUT6 #(
    .INIT(64'hFEFFFFFF19FF0000)) 
    fch_issu1_inferred_i_129
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[3]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_129_n_0));
  MUXF7 fch_issu1_inferred_i_13
       (.I0(fch_issu1_inferred_i_42_n_0),
        .I1(fch_issu1_inferred_i_43_n_0),
        .O(fch_issu1_inferred_i_13_n_0),
        .S(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAA2882)) 
    fch_issu1_inferred_i_130
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[15]),
        .I5(fch_issu1_inferred_i_179_n_0),
        .O(fch_issu1_inferred_i_130_n_0));
  LUT5 #(
    .INIT(32'h2A6F2AEF)) 
    fch_issu1_inferred_i_131
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .I2(fdat[13]),
        .I3(fdat[12]),
        .I4(fdat[11]),
        .O(fch_issu1_inferred_i_131_n_0));
  LUT6 #(
    .INIT(64'h4444444440444444)) 
    fch_issu1_inferred_i_132
       (.I0(fdat[11]),
        .I1(fdat[14]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(fdat[8]),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_132_n_0));
  LUT5 #(
    .INIT(32'h44CC7FDD)) 
    fch_issu1_inferred_i_133
       (.I0(fdatx[13]),
        .I1(fdatx[15]),
        .I2(fdatx[11]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .O(fch_issu1_inferred_i_133_n_0));
  LUT6 #(
    .INIT(64'h4444444440444444)) 
    fch_issu1_inferred_i_134
       (.I0(fdatx[11]),
        .I1(fdatx[14]),
        .I2(fdatx[9]),
        .I3(fdatx[10]),
        .I4(fdatx[8]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_134_n_0));
  LUT6 #(
    .INIT(64'h5050505045555050)) 
    fch_issu1_inferred_i_135
       (.I0(fch_issu1_inferred_i_180_n_0),
        .I1(fch_issu1_inferred_i_181_n_0),
        .I2(fdatx[7]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_182_n_0),
        .O(fch_issu1_inferred_i_135_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAAA)) 
    fch_issu1_inferred_i_136
       (.I0(fch_issu1_inferred_i_145_n_0),
        .I1(fch_issu1_inferred_i_122_n_0),
        .I2(fdatx[15]),
        .I3(fdatx[11]),
        .I4(fdatx[13]),
        .I5(fch_issu1_inferred_i_183_n_0),
        .O(fch_issu1_inferred_i_136_n_0));
  LUT6 #(
    .INIT(64'hAFAEAAAEFFFFFFFF)) 
    fch_issu1_inferred_i_137
       (.I0(fch_issu1_inferred_i_150_n_0),
        .I1(fdatx[7]),
        .I2(fch_issu1_inferred_i_184_n_0),
        .I3(fdatx[8]),
        .I4(fdatx[2]),
        .I5(fch_issu1_inferred_i_185_n_0),
        .O(fch_issu1_inferred_i_137_n_0));
  LUT5 #(
    .INIT(32'h00EC0000)) 
    fch_issu1_inferred_i_138
       (.I0(fch_issu1_inferred_i_165_n_0),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[11]),
        .I4(fdatx[12]),
        .O(fch_issu1_inferred_i_138_n_0));
  LUT6 #(
    .INIT(64'hAAAA08A8AAAAA8A8)) 
    fch_issu1_inferred_i_139
       (.I0(fdatx[10]),
        .I1(fdatx[2]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[9]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_139_n_0));
  MUXF7 fch_issu1_inferred_i_14
       (.I0(fch_issu1_inferred_i_44_n_0),
        .I1(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_14_n_0),
        .S(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hC1C0C0C0C0C0C0C0)) 
    fch_issu1_inferred_i_140
       (.I0(fdatx[12]),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(\ir0_id_fl[20]_i_8_n_0 ),
        .I4(fch_issu1_inferred_i_186_n_0),
        .I5(fch_issu1_inferred_i_187_n_0),
        .O(fch_issu1_inferred_i_140_n_0));
  LUT6 #(
    .INIT(64'h0040000000000000)) 
    fch_issu1_inferred_i_141
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .I2(fdat[6]),
        .I3(fdat[7]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_141_n_0));
  LUT6 #(
    .INIT(64'h000000000441FFFF)) 
    fch_issu1_inferred_i_142
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(\nir_id[17]_i_2_n_0 ),
        .I5(fch_issu1_inferred_i_188_n_0),
        .O(fch_issu1_inferred_i_142_n_0));
  LUT6 #(
    .INIT(64'h000000000441FFFF)) 
    fch_issu1_inferred_i_143
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fch_issu1_inferred_i_119_n_0),
        .I5(fch_issu1_inferred_i_189_n_0),
        .O(fch_issu1_inferred_i_143_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_144
       (.I0(fdatx[8]),
        .I1(fdatx[10]),
        .O(fch_issu1_inferred_i_144_n_0));
  LUT6 #(
    .INIT(64'hFFFF1110FFFFFFFF)) 
    fch_issu1_inferred_i_145
       (.I0(fdatx[13]),
        .I1(fdatx[15]),
        .I2(fdatx[12]),
        .I3(fdatx[14]),
        .I4(\fch/stat [0]),
        .I5(\fch/stat [1]),
        .O(fch_issu1_inferred_i_145_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    fch_issu1_inferred_i_146
       (.I0(fdatx[7]),
        .I1(fdatx[3]),
        .I2(fdatx[10]),
        .I3(fdatx[9]),
        .I4(fdatx[8]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_146_n_0));
  LUT6 #(
    .INIT(64'hAAAA08A8AAAAA8A8)) 
    fch_issu1_inferred_i_147
       (.I0(fdatx[10]),
        .I1(fdatx[1]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[9]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_147_n_0));
  LUT6 #(
    .INIT(64'h888A8A8AAAAAAAAA)) 
    fch_issu1_inferred_i_148
       (.I0(fch_issu1_inferred_i_185_n_0),
        .I1(fch_issu1_inferred_i_190_n_0),
        .I2(fdatx[9]),
        .I3(fdatx[1]),
        .I4(fdatx[8]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_148_n_0));
  LUT6 #(
    .INIT(64'hF7550000FFFFFFFF)) 
    fch_issu1_inferred_i_149
       (.I0(fdatx[10]),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fch_issu1_inferred_i_191_n_0),
        .I4(fch_issu1_inferred_i_138_n_0),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_149_n_0));
  LUT6 #(
    .INIT(64'h0000FF0F77077707)) 
    fch_issu1_inferred_i_15
       (.I0(\fch/lir_id_0 [19]),
        .I1(\fch/fadr_1_fl ),
        .I2(fch_issu1_inferred_i_46_n_0),
        .I3(fch_issu1_inferred_i_47_n_0),
        .I4(\fch/nir_id [19]),
        .I5(fch_issu1_inferred_i_20_n_0),
        .O(fch_issu1_inferred_i_15_n_0));
  LUT3 #(
    .INIT(8'h08)) 
    fch_issu1_inferred_i_150
       (.I0(fdatx[9]),
        .I1(fdatx[10]),
        .I2(fch_issu1_inferred_i_192_n_0),
        .O(fch_issu1_inferred_i_150_n_0));
  LUT6 #(
    .INIT(64'h7777F777FF777777)) 
    fch_issu1_inferred_i_151
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .I2(fdatx[0]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_151_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    fch_issu1_inferred_i_152
       (.I0(fdatx[15]),
        .I1(fdatx[13]),
        .I2(fdatx[12]),
        .O(fch_issu1_inferred_i_152_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_153
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .O(fch_issu1_inferred_i_153_n_0));
  LUT6 #(
    .INIT(64'h40FF40FF40FFFFFF)) 
    fch_issu1_inferred_i_154
       (.I0(fch_issu1_inferred_i_193_n_0),
        .I1(fch_issu1_inferred_i_177_n_0),
        .I2(fch_issu1_inferred_i_194_n_0),
        .I3(fdatx[9]),
        .I4(fdatx[1]),
        .I5(fch_issu1_inferred_i_168_n_0),
        .O(fch_issu1_inferred_i_154_n_0));
  LUT4 #(
    .INIT(16'h4D6C)) 
    fch_issu1_inferred_i_155
       (.I0(fdatx[1]),
        .I1(fdatx[2]),
        .I2(fdatx[3]),
        .I3(fdatx[0]),
        .O(fch_issu1_inferred_i_155_n_0));
  LUT4 #(
    .INIT(16'hE551)) 
    fch_issu1_inferred_i_156
       (.I0(fdat[2]),
        .I1(fdat[0]),
        .I2(fdat[1]),
        .I3(fdat[3]),
        .O(fch_issu1_inferred_i_156_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_157
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .O(fch_issu1_inferred_i_157_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_158
       (.I0(fdatx[10]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_158_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_159
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(fch_issu1_inferred_i_159_n_0));
  LUT6 #(
    .INIT(64'hFF80FF80FFFFFF80)) 
    fch_issu1_inferred_i_16
       (.I0(fch_issu1_inferred_i_20_n_0),
        .I1(fch_issu1_inferred_i_48_n_0),
        .I2(fch_issu1_inferred_i_49_n_0),
        .I3(fch_issu1_inferred_i_50_n_0),
        .I4(fch_issu1_inferred_i_51_n_0),
        .I5(fch_issu1_inferred_i_52_n_0),
        .O(fch_issu1_inferred_i_16_n_0));
  LUT6 #(
    .INIT(64'h8000000080000040)) 
    fch_issu1_inferred_i_160
       (.I0(fdatx[9]),
        .I1(fch_issu1_inferred_i_195_n_0),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(fdatx[7]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_160_n_0));
  LUT4 #(
    .INIT(16'hEEEA)) 
    fch_issu1_inferred_i_161
       (.I0(fdatx[13]),
        .I1(fdatx[0]),
        .I2(fdatx[3]),
        .I3(fdatx[2]),
        .O(fch_issu1_inferred_i_161_n_0));
  LUT4 #(
    .INIT(16'hBFEA)) 
    fch_issu1_inferred_i_162
       (.I0(fdatx[0]),
        .I1(fdatx[3]),
        .I2(fdatx[2]),
        .I3(fdatx[1]),
        .O(fch_issu1_inferred_i_162_n_0));
  LUT6 #(
    .INIT(64'hAA00AA0000000200)) 
    fch_issu1_inferred_i_163
       (.I0(fch_issu1_inferred_i_196_n_0),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[8]),
        .I4(fdat[1]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_163_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF0F0FFFEF)) 
    fch_issu1_inferred_i_164
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[8]),
        .I3(fdatx[1]),
        .I4(fdatx[6]),
        .I5(fch_issu1_inferred_i_197_n_0),
        .O(fch_issu1_inferred_i_164_n_0));
  LUT3 #(
    .INIT(8'h10)) 
    fch_issu1_inferred_i_165
       (.I0(fdatx[6]),
        .I1(fdatx[8]),
        .I2(fdatx[7]),
        .O(fch_issu1_inferred_i_165_n_0));
  LUT6 #(
    .INIT(64'h0A2A000A2000000A)) 
    fch_issu1_inferred_i_166
       (.I0(fdatx[8]),
        .I1(fdatx[3]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_166_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFDFFFFFFD)) 
    fch_issu1_inferred_i_167
       (.I0(fdatx[8]),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .I3(fdatx[4]),
        .I4(fdatx[5]),
        .I5(fdatx[3]),
        .O(fch_issu1_inferred_i_167_n_0));
  LUT5 #(
    .INIT(32'h4FFFFFFF)) 
    fch_issu1_inferred_i_168
       (.I0(fdatx[3]),
        .I1(fdatx[5]),
        .I2(fdatx[8]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .O(fch_issu1_inferred_i_168_n_0));
  LUT6 #(
    .INIT(64'h2020222002200220)) 
    fch_issu1_inferred_i_169
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[7]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_169_n_0));
  LUT6 #(
    .INIT(64'h0100515551555155)) 
    fch_issu1_inferred_i_17
       (.I0(fch_issu1_inferred_i_53_n_0),
        .I1(\fch/nir_id [16]),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(\fch/lir_id_0 [16]),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hCFDFCFDFFFDFCFDF)) 
    fch_issu1_inferred_i_170
       (.I0(fdatx[7]),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[11]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_170_n_0));
  LUT5 #(
    .INIT(32'h08C80B8B)) 
    fch_issu1_inferred_i_171
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[5]),
        .I3(fdatx[3]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_171_n_0));
  LUT5 #(
    .INIT(32'h08C80B8B)) 
    fch_issu1_inferred_i_172
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[3]),
        .I4(fdat[4]),
        .O(fch_issu1_inferred_i_172_n_0));
  LUT4 #(
    .INIT(16'h8AAA)) 
    fch_issu1_inferred_i_173
       (.I0(fdatx[9]),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fch_issu1_inferred_i_198_n_0),
        .O(fch_issu1_inferred_i_173_n_0));
  LUT6 #(
    .INIT(64'hFFFFA0FFFFFFFCFF)) 
    fch_issu1_inferred_i_174
       (.I0(fdatx[3]),
        .I1(fdatx[4]),
        .I2(fdatx[5]),
        .I3(fdatx[8]),
        .I4(fdatx[2]),
        .I5(fdatx[6]),
        .O(fch_issu1_inferred_i_174_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_175
       (.I0(fdat[1]),
        .I1(fdat[8]),
        .O(fch_issu1_inferred_i_175_n_0));
  LUT5 #(
    .INIT(32'h5F5F5F4F)) 
    fch_issu1_inferred_i_176
       (.I0(fdatx[6]),
        .I1(fdatx[2]),
        .I2(fdatx[8]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_176_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_177
       (.I0(fdatx[6]),
        .I1(fdatx[3]),
        .O(fch_issu1_inferred_i_177_n_0));
  LUT6 #(
    .INIT(64'h000F000F000F080F)) 
    fch_issu1_inferred_i_178
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[7]),
        .I3(fdatx[6]),
        .I4(fdatx[3]),
        .I5(fdatx[2]),
        .O(fch_issu1_inferred_i_178_n_0));
  LUT5 #(
    .INIT(32'h2330C330)) 
    fch_issu1_inferred_i_179
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[5]),
        .O(fch_issu1_inferred_i_179_n_0));
  LUT5 #(
    .INIT(32'h00B0BBBB)) 
    fch_issu1_inferred_i_18
       (.I0(fdatx[10]),
        .I1(fch_issu1_inferred_i_54_n_0),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_55_n_0),
        .I4(fch_issu1_inferred_i_56_n_0),
        .O(fch_issu1_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hEEFEFEEEFEEEEEFE)) 
    fch_issu1_inferred_i_180
       (.I0(fch_issu1_inferred_i_199_n_0),
        .I1(fch_issu1_inferred_i_200_n_0),
        .I2(fdatx[11]),
        .I3(fdatx[8]),
        .I4(fdatx[9]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_180_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_181
       (.I0(fdatx[3]),
        .I1(fdatx[5]),
        .O(fch_issu1_inferred_i_181_n_0));
  LUT4 #(
    .INIT(16'h8CC0)) 
    fch_issu1_inferred_i_182
       (.I0(fdatx[3]),
        .I1(fdatx[8]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .O(fch_issu1_inferred_i_182_n_0));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    fch_issu1_inferred_i_183
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[1]),
        .I3(fdatx[8]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_183_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_184
       (.I0(fdatx[9]),
        .I1(fdatx[10]),
        .O(fch_issu1_inferred_i_184_n_0));
  LUT5 #(
    .INIT(32'h88880888)) 
    fch_issu1_inferred_i_185
       (.I0(fdatx[11]),
        .I1(fdatx[12]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .O(fch_issu1_inferred_i_185_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_186
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(fch_issu1_inferred_i_186_n_0));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    fch_issu1_inferred_i_187
       (.I0(fdatx[0]),
        .I1(fdatx[1]),
        .I2(fch_issu1_inferred_i_201_n_0),
        .I3(fch_issu1_inferred_i_104_n_0),
        .I4(fdatx[10]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_187_n_0));
  LUT6 #(
    .INIT(64'hCCCFFFCFDFFFDFFF)) 
    fch_issu1_inferred_i_188
       (.I0(fdat[7]),
        .I1(fdat[15]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_188_n_0));
  LUT6 #(
    .INIT(64'hCCCFFFCFDFFFDFFF)) 
    fch_issu1_inferred_i_189
       (.I0(fdatx[7]),
        .I1(fdatx[15]),
        .I2(fdatx[6]),
        .I3(fdatx[8]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_189_n_0));
  LUT6 #(
    .INIT(64'h20AAA0AAA8AAA0AA)) 
    fch_issu1_inferred_i_19
       (.I0(fch_issu1_inferred_i_57_n_0),
        .I1(\nir_id[17]_i_2_n_0 ),
        .I2(fdat[5]),
        .I3(fch_issu1_inferred_i_58_n_0),
        .I4(fdat[9]),
        .I5(fch_issu1_inferred_i_59_n_0),
        .O(fch_issu1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h0505055010000005)) 
    fch_issu1_inferred_i_190
       (.I0(\ir0_id_fl[21]_i_9_n_0 ),
        .I1(fdatx[3]),
        .I2(fdatx[5]),
        .I3(fdatx[4]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_190_n_0));
  LUT4 #(
    .INIT(16'h2033)) 
    fch_issu1_inferred_i_191
       (.I0(fdatx[7]),
        .I1(fdatx[9]),
        .I2(fdatx[6]),
        .I3(fdatx[8]),
        .O(fch_issu1_inferred_i_191_n_0));
  LUT6 #(
    .INIT(64'hAA0A2000AAA8000A)) 
    fch_issu1_inferred_i_192
       (.I0(fdatx[8]),
        .I1(fdatx[3]),
        .I2(fdatx[4]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_192_n_0));
  LUT5 #(
    .INIT(32'h5F5F5F4F)) 
    fch_issu1_inferred_i_193
       (.I0(fdatx[6]),
        .I1(fdatx[1]),
        .I2(fdatx[8]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .O(fch_issu1_inferred_i_193_n_0));
  LUT6 #(
    .INIT(64'h000000000008FFFF)) 
    fch_issu1_inferred_i_194
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[1]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_194_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_195
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .O(fch_issu1_inferred_i_195_n_0));
  LUT6 #(
    .INIT(64'h33333F333F3B3F33)) 
    fch_issu1_inferred_i_196
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[1]),
        .I3(fdat[7]),
        .I4(fdat[5]),
        .I5(fdat[3]),
        .O(fch_issu1_inferred_i_196_n_0));
  LUT6 #(
    .INIT(64'hCCC0C4C4CCC4C4C4)) 
    fch_issu1_inferred_i_197
       (.I0(fdatx[7]),
        .I1(fdatx[6]),
        .I2(fdatx[1]),
        .I3(fdatx[3]),
        .I4(fdatx[5]),
        .I5(fdatx[4]),
        .O(fch_issu1_inferred_i_197_n_0));
  LUT5 #(
    .INIT(32'hBB004001)) 
    fch_issu1_inferred_i_198
       (.I0(fdatx[3]),
        .I1(fdatx[5]),
        .I2(fdatx[4]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .O(fch_issu1_inferred_i_198_n_0));
  LUT5 #(
    .INIT(32'h00008FF0)) 
    fch_issu1_inferred_i_199
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .O(fch_issu1_inferred_i_199_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF14000014)) 
    fch_issu1_inferred_i_2
       (.I0(fch_issu1_inferred_i_8_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_11_n_0),
        .I5(fch_issu1_inferred_i_12_n_0),
        .O(fch_issu1_inferred_i_2_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_20
       (.I0(\fch/stat [1]),
        .I1(\fch/stat [0]),
        .O(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h88888888F8888888)) 
    fch_issu1_inferred_i_200
       (.I0(fdatx[11]),
        .I1(fdatx[15]),
        .I2(fdatx[8]),
        .I3(fdatx[9]),
        .I4(fdatx[6]),
        .I5(fdatx[5]),
        .O(fch_issu1_inferred_i_200_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_201
       (.I0(fdatx[3]),
        .I1(fdatx[2]),
        .O(fch_issu1_inferred_i_201_n_0));
  LUT5 #(
    .INIT(32'h04555555)) 
    fch_issu1_inferred_i_21
       (.I0(\fch/fadr_1_fl ),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fdat[13]),
        .O(fch_issu1_inferred_i_21_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_22
       (.I0(\fch/fadr_1_fl ),
        .I1(fdat[15]),
        .O(fch_issu1_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'h00A20000AAAAAAAA)) 
    fch_issu1_inferred_i_23
       (.I0(fch_issu1_inferred_i_60_n_0),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdatx[10]),
        .I5(fch_issu1_inferred_i_61_n_0),
        .O(fch_issu1_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hF3A200A2FFAE0CAE)) 
    fch_issu1_inferred_i_24
       (.I0(fch_issu1_inferred_i_62_n_0),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fch_issu1_inferred_i_63_n_0),
        .I5(\fch/nir_id [15]),
        .O(fch_issu1_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'h000000000000FFBA)) 
    fch_issu1_inferred_i_25
       (.I0(fch_issu1_inferred_i_64_n_0),
        .I1(fch_issu1_inferred_i_65_n_0),
        .I2(fch_issu1_inferred_i_66_n_0),
        .I3(fch_issu1_inferred_i_67_n_0),
        .I4(fch_issu1_inferred_i_68_n_0),
        .I5(fch_issu1_inferred_i_69_n_0),
        .O(fch_issu1_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'h4744777747444744)) 
    fch_issu1_inferred_i_26
       (.I0(\fch/nir_id [14]),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(fch_issu1_inferred_i_70_n_0),
        .I3(fch_issu1_inferred_i_71_n_0),
        .I4(\fch/lir_id_0 [14]),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hEE0EEE0E0000EE0E)) 
    fch_issu1_inferred_i_27
       (.I0(fch_issu1_inferred_i_72_n_0),
        .I1(fch_issu1_inferred_i_73_n_0),
        .I2(fch_issu1_inferred_i_74_n_0),
        .I3(fch_issu1_inferred_i_75_n_0),
        .I4(\fch/fadr_1_fl ),
        .I5(fch_issu1_inferred_i_20_n_0),
        .O(fch_issu1_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'h7777474447444744)) 
    fch_issu1_inferred_i_28
       (.I0(\fch/nir_id [13]),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(fch_issu1_inferred_i_76_n_0),
        .I3(fch_issu1_inferred_i_71_n_0),
        .I4(\fch/fadr_1_fl ),
        .I5(\nir_id[13]_i_2_n_0 ),
        .O(fch_issu1_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h20EF202020EF20EF)) 
    fch_issu1_inferred_i_29
       (.I0(\fch/nir_id [12]),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [1]),
        .I3(fch_issu1_inferred_i_77_n_0),
        .I4(\fch/lir_id_0 [12]),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFF6FF66FF6FFFF)) 
    fch_issu1_inferred_i_3
       (.I0(fch_issu1_inferred_i_9_n_0),
        .I1(fch_issu1_inferred_i_13_n_0),
        .I2(fch_issu1_inferred_i_14_n_0),
        .I3(fch_issu1_inferred_i_15_n_0),
        .I4(fch_issu1_inferred_i_16_n_0),
        .I5(fch_issu1_inferred_i_17_n_0),
        .O(fch_issu1_inferred_i_3_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    fch_issu1_inferred_i_30
       (.I0(fch_issu1_inferred_i_13_n_0),
        .I1(fch_issu1_inferred_i_28_n_0),
        .I2(fch_issu1_inferred_i_14_n_0),
        .I3(fch_issu1_inferred_i_24_n_0),
        .I4(fch_issu1_inferred_i_29_n_0),
        .I5(fch_issu1_inferred_i_16_n_0),
        .O(fch_issu1_inferred_i_30_n_0));
  LUT4 #(
    .INIT(16'hF99F)) 
    fch_issu1_inferred_i_31
       (.I0(fch_issu1_inferred_i_34_n_0),
        .I1(fch_issu1_inferred_i_24_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_28_n_0),
        .O(fch_issu1_inferred_i_31_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    fch_issu1_inferred_i_32
       (.I0(fch_issu1_inferred_i_29_n_0),
        .I1(fch_issu1_inferred_i_33_n_0),
        .O(fch_issu1_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'hFF4F0000FF4FFF4F)) 
    fch_issu1_inferred_i_33
       (.I0(\fch/stat [0]),
        .I1(\fch/stat [1]),
        .I2(fdat[0]),
        .I3(fch_issu1_inferred_i_36_n_0),
        .I4(fch_issu1_inferred_i_78_n_0),
        .I5(fch_issu1_inferred_i_79_n_0),
        .O(fch_issu1_inferred_i_33_n_0));
  MUXF7 fch_issu1_inferred_i_34
       (.I0(fch_issu1_inferred_i_80_n_0),
        .I1(fch_issu1_inferred_i_81_n_0),
        .O(fch_issu1_inferred_i_34_n_0),
        .S(fch_issu1_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'h00A20000AAAAAAAA)) 
    fch_issu1_inferred_i_35
       (.I0(fch_issu1_inferred_i_82_n_0),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_61_n_0),
        .O(fch_issu1_inferred_i_35_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF00005D7D)) 
    fch_issu1_inferred_i_36
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(\nir_id[14]_i_9_n_0 ),
        .I4(fdat[11]),
        .I5(fch_issu1_inferred_i_83_n_0),
        .O(fch_issu1_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'h00C0F000F0B0F000)) 
    fch_issu1_inferred_i_37
       (.I0(fch_issu1_inferred_i_84_n_0),
        .I1(fdatx[8]),
        .I2(fch_issu1_inferred_i_48_n_0),
        .I3(fdatx[11]),
        .I4(fdatx[10]),
        .I5(fdatx[9]),
        .O(fch_issu1_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'h0900000000000900)) 
    fch_issu1_inferred_i_38
       (.I0(fch_issu1_inferred_i_27_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_15_n_0),
        .I3(fch_issu1_inferred_i_17_n_0),
        .I4(fch_issu1_inferred_i_5_n_0),
        .I5(fch_issu1_inferred_i_25_n_0),
        .O(fch_issu1_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFFB0)) 
    fch_issu1_inferred_i_39
       (.I0(fch_issu1_inferred_i_85_n_0),
        .I1(fch_issu1_inferred_i_86_n_0),
        .I2(fdatx[12]),
        .I3(fdatx[15]),
        .I4(fch_issu1_inferred_i_87_n_0),
        .I5(\fch/nir_id [24]),
        .O(fch_issu1_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'hACACACACAFAFACAF)) 
    fch_issu1_inferred_i_4
       (.I0(fch_issu1_inferred_i_18_n_0),
        .I1(fch_issu1_inferred_i_19_n_0),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(fch_issu1_inferred_i_21_n_0),
        .I4(fdat[10]),
        .I5(fch_issu1_inferred_i_22_n_0),
        .O(fch_issu1_inferred_i_4_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF1011)) 
    fch_issu1_inferred_i_40
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_88_n_0),
        .I2(fch_issu1_inferred_i_89_n_0),
        .I3(fdat[12]),
        .I4(fch_issu1_inferred_i_90_n_0),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBABB)) 
    fch_issu1_inferred_i_41
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_91_n_0),
        .I2(fch_issu1_inferred_i_92_n_0),
        .I3(fch_issu1_inferred_i_93_n_0),
        .I4(fdatx[10]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_41_n_0));
  LUT6 #(
    .INIT(64'h0000F200F2F2F2F2)) 
    fch_issu1_inferred_i_42
       (.I0(fch_issu1_inferred_i_21_n_0),
        .I1(fdat[9]),
        .I2(fch_issu1_inferred_i_22_n_0),
        .I3(fch_issu1_inferred_i_94_n_0),
        .I4(fch_issu1_inferred_i_95_n_0),
        .I5(fch_issu1_inferred_i_57_n_0),
        .O(fch_issu1_inferred_i_42_n_0));
  LUT5 #(
    .INIT(32'hF4FF4444)) 
    fch_issu1_inferred_i_43
       (.I0(fdatx[9]),
        .I1(fch_issu1_inferred_i_54_n_0),
        .I2(fch_issu1_inferred_i_96_n_0),
        .I3(fdatx[14]),
        .I4(fch_issu1_inferred_i_56_n_0),
        .O(fch_issu1_inferred_i_43_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAA80888888)) 
    fch_issu1_inferred_i_44
       (.I0(fch_issu1_inferred_i_97_n_0),
        .I1(fch_issu1_inferred_i_58_n_0),
        .I2(fch_issu1_inferred_i_98_n_0),
        .I3(fch_issu1_inferred_i_99_n_0),
        .I4(fdat[11]),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_44_n_0));
  LUT6 #(
    .INIT(64'h0400FFFF04000400)) 
    fch_issu1_inferred_i_45
       (.I0(fch_issu1_inferred_i_100_n_0),
        .I1(fch_issu1_inferred_i_48_n_0),
        .I2(fch_issu1_inferred_i_101_n_0),
        .I3(fch_issu1_inferred_i_102_n_0),
        .I4(fch_issu1_inferred_i_90_n_0),
        .I5(fch_issu1_inferred_i_54_n_0),
        .O(fch_issu1_inferred_i_45_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF55003000)) 
    fch_issu1_inferred_i_46
       (.I0(fch_issu1_inferred_i_103_n_0),
        .I1(fch_issu1_inferred_i_104_n_0),
        .I2(fch_issu1_inferred_i_105_n_0),
        .I3(fdatx[11]),
        .I4(fdatx[10]),
        .I5(fch_issu1_inferred_i_106_n_0),
        .O(fch_issu1_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'h3BBBB33B33BBBBBB)) 
    fch_issu1_inferred_i_47
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_107_n_0),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .I4(fdatx[12]),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_47_n_0));
  LUT4 #(
    .INIT(16'h0080)) 
    fch_issu1_inferred_i_48
       (.I0(fdatx[14]),
        .I1(fdatx[12]),
        .I2(fdatx[13]),
        .I3(fdatx[15]),
        .O(fch_issu1_inferred_i_48_n_0));
  LUT6 #(
    .INIT(64'h5530550030303030)) 
    fch_issu1_inferred_i_49
       (.I0(fch_issu1_inferred_i_108_n_0),
        .I1(fch_issu1_inferred_i_100_n_0),
        .I2(fdatx[3]),
        .I3(fdatx[10]),
        .I4(fch_issu1_inferred_i_109_n_0),
        .I5(fdatx[11]),
        .O(fch_issu1_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h00000000770F7777)) 
    fch_issu1_inferred_i_5
       (.I0(\fch/lir_id_0 [18]),
        .I1(\fch/fadr_1_fl ),
        .I2(\fch/nir_id [18]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fch_issu1_inferred_i_23_n_0),
        .O(fch_issu1_inferred_i_5_n_0));
  LUT6 #(
    .INIT(64'hFF04040404040404)) 
    fch_issu1_inferred_i_50
       (.I0(fch_issu1_inferred_i_110_n_0),
        .I1(fdat[15]),
        .I2(fch_issu1_inferred_i_111_n_0),
        .I3(fch_issu1_inferred_i_20_n_0),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_54_n_0),
        .O(fch_issu1_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'h5530550030303030)) 
    fch_issu1_inferred_i_51
       (.I0(fch_issu1_inferred_i_112_n_0),
        .I1(fch_issu1_inferred_i_113_n_0),
        .I2(fdat[3]),
        .I3(fdat[10]),
        .I4(fch_issu1_inferred_i_114_n_0),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_51_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7F)) 
    fch_issu1_inferred_i_52
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_20_n_0),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_52_n_0));
  LUT6 #(
    .INIT(64'h000E0000EEEEEEEE)) 
    fch_issu1_inferred_i_53
       (.I0(fch_issu1_inferred_i_115_n_0),
        .I1(fch_issu1_inferred_i_106_n_0),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(\fch/fadr_1_fl ),
        .I4(fdatx[8]),
        .I5(fch_issu1_inferred_i_61_n_0),
        .O(fch_issu1_inferred_i_53_n_0));
  LUT5 #(
    .INIT(32'h0AAA8AAA)) 
    fch_issu1_inferred_i_54
       (.I0(fdatx[15]),
        .I1(fdatx[11]),
        .I2(fdatx[12]),
        .I3(fdatx[13]),
        .I4(fdatx[14]),
        .O(fch_issu1_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'h0008000B000000FF)) 
    fch_issu1_inferred_i_55
       (.I0(fch_issu1_inferred_i_116_n_0),
        .I1(fdatx[9]),
        .I2(fch_issu1_inferred_i_117_n_0),
        .I3(fch_issu1_inferred_i_118_n_0),
        .I4(fdatx[5]),
        .I5(fch_issu1_inferred_i_119_n_0),
        .O(fch_issu1_inferred_i_55_n_0));
  LUT5 #(
    .INIT(32'h55550004)) 
    fch_issu1_inferred_i_56
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_120_n_0),
        .I2(fch_issu1_inferred_i_121_n_0),
        .I3(fch_issu1_inferred_i_122_n_0),
        .I4(fdatx[14]),
        .O(fch_issu1_inferred_i_56_n_0));
  LUT6 #(
    .INIT(64'h5555555155555555)) 
    fch_issu1_inferred_i_57
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_123_n_0),
        .I2(fdat[14]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fch_issu1_inferred_i_124_n_0),
        .O(fch_issu1_inferred_i_57_n_0));
  LUT6 #(
    .INIT(64'hAAAAAA8AAAAAAAAA)) 
    fch_issu1_inferred_i_58
       (.I0(fch_issu1_inferred_i_94_n_0),
        .I1(fdat[9]),
        .I2(\nir_id[17]_i_2_n_0 ),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_58_n_0));
  LUT6 #(
    .INIT(64'h00000000F8F0FFFF)) 
    fch_issu1_inferred_i_59
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(\nir_id[14]_i_11_n_0 ),
        .I4(fdat[6]),
        .I5(fch_issu1_inferred_i_125_n_0),
        .O(fch_issu1_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBEFFFFBE)) 
    fch_issu1_inferred_i_6
       (.I0(fch_issu1_inferred_i_24_n_0),
        .I1(fch_issu1_inferred_i_25_n_0),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fch_issu1_inferred_i_27_n_0),
        .I4(fch_issu1_inferred_i_28_n_0),
        .I5(fch_issu1_inferred_i_29_n_0),
        .O(fch_issu1_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFDFFFDDFFFFFF00)) 
    fch_issu1_inferred_i_60
       (.I0(fch_issu1_inferred_i_126_n_0),
        .I1(fch_issu1_inferred_i_127_n_0),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_106_n_0),
        .I4(fdatx[5]),
        .I5(fch_issu1_inferred_i_119_n_0),
        .O(fch_issu1_inferred_i_60_n_0));
  LUT6 #(
    .INIT(64'h77BF0000FFFFFFFF)) 
    fch_issu1_inferred_i_61
       (.I0(fdatx[14]),
        .I1(fdatx[13]),
        .I2(fdatx[11]),
        .I3(fdatx[12]),
        .I4(fdatx[15]),
        .I5(fch_issu1_inferred_i_107_n_0),
        .O(fch_issu1_inferred_i_61_n_0));
  LUT5 #(
    .INIT(32'h00820000)) 
    fch_issu1_inferred_i_62
       (.I0(fch_issu1_inferred_i_48_n_0),
        .I1(fdatx[8]),
        .I2(fdatx[11]),
        .I3(fdatx[9]),
        .I4(fdatx[10]),
        .O(fch_issu1_inferred_i_62_n_0));
  LUT6 #(
    .INIT(64'h0000200200000000)) 
    fch_issu1_inferred_i_63
       (.I0(\nir_id[15]_i_2_n_0 ),
        .I1(fdat[15]),
        .I2(fdat[8]),
        .I3(fdat[11]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_63_n_0));
  LUT6 #(
    .INIT(64'h444F444F444F4444)) 
    fch_issu1_inferred_i_64
       (.I0(\fch/stat [0]),
        .I1(\fch/stat [1]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_64_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    fch_issu1_inferred_i_65
       (.I0(fdat[5]),
        .I1(fdat[2]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fch_issu1_inferred_i_128_n_0),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_65_n_0));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    fch_issu1_inferred_i_66
       (.I0(fdat[8]),
        .I1(fdat[1]),
        .I2(fdat[3]),
        .I3(fdat[4]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'h0000000000002FFF)) 
    fch_issu1_inferred_i_67
       (.I0(fch_issu1_inferred_i_129_n_0),
        .I1(fch_issu1_inferred_i_130_n_0),
        .I2(fdat[12]),
        .I3(fdat[14]),
        .I4(fch_issu1_inferred_i_131_n_0),
        .I5(fch_issu1_inferred_i_132_n_0),
        .O(fch_issu1_inferred_i_67_n_0));
  LUT6 #(
    .INIT(64'h00000000EEEEFEEE)) 
    fch_issu1_inferred_i_68
       (.I0(fch_issu1_inferred_i_133_n_0),
        .I1(fch_issu1_inferred_i_134_n_0),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fch_issu1_inferred_i_135_n_0),
        .I5(fch_issu1_inferred_i_136_n_0),
        .O(fch_issu1_inferred_i_68_n_0));
  LUT3 #(
    .INIT(8'h8A)) 
    fch_issu1_inferred_i_69
       (.I0(\fch/fadr_1_fl ),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [1]),
        .O(fch_issu1_inferred_i_69_n_0));
  LUT6 #(
    .INIT(64'h1F11444F11114444)) 
    fch_issu1_inferred_i_7
       (.I0(fch_issu1_inferred_i_30_n_0),
        .I1(fch_issu1_inferred_i_4_n_0),
        .I2(fch_issu1_inferred_i_31_n_0),
        .I3(fch_issu1_inferred_i_11_n_0),
        .I4(fch_issu1_inferred_i_26_n_0),
        .I5(fch_issu1_inferred_i_32_n_0),
        .O(fch_issu1_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'h4040004055555555)) 
    fch_issu1_inferred_i_70
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_137_n_0),
        .I2(fdatx[14]),
        .I3(fch_issu1_inferred_i_138_n_0),
        .I4(fch_issu1_inferred_i_139_n_0),
        .I5(fch_issu1_inferred_i_140_n_0),
        .O(fch_issu1_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'h1145014555555555)) 
    fch_issu1_inferred_i_71
       (.I0(\fch/fadr_1_fl ),
        .I1(fdatx[13]),
        .I2(fdatx[14]),
        .I3(fdatx[12]),
        .I4(fdatx[11]),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_71_n_0));
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_72
       (.I0(fch_issu1_inferred_i_64_n_0),
        .I1(fdat[15]),
        .I2(fdat[8]),
        .I3(fdat[4]),
        .I4(fdat[12]),
        .I5(fch_issu1_inferred_i_141_n_0),
        .O(fch_issu1_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'h00000000BB0BFFFF)) 
    fch_issu1_inferred_i_73
       (.I0(fch_issu1_inferred_i_142_n_0),
        .I1(fdat[12]),
        .I2(\nir_id[12]_i_4_n_0 ),
        .I3(fdat[11]),
        .I4(fdat[14]),
        .I5(fch_issu1_inferred_i_131_n_0),
        .O(fch_issu1_inferred_i_73_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF44004F00)) 
    fch_issu1_inferred_i_74
       (.I0(fch_issu1_inferred_i_143_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[11]),
        .I3(fdatx[14]),
        .I4(fch_issu1_inferred_i_144_n_0),
        .I5(fch_issu1_inferred_i_133_n_0),
        .O(fch_issu1_inferred_i_74_n_0));
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_75
       (.I0(fch_issu1_inferred_i_145_n_0),
        .I1(fch_issu1_inferred_i_146_n_0),
        .I2(fdatx[6]),
        .I3(fdatx[5]),
        .I4(fdatx[4]),
        .I5(fdatx[12]),
        .O(fch_issu1_inferred_i_75_n_0));
  LUT6 #(
    .INIT(64'h0051555555555555)) 
    fch_issu1_inferred_i_76
       (.I0(fdatx[15]),
        .I1(fch_issu1_inferred_i_138_n_0),
        .I2(fch_issu1_inferred_i_147_n_0),
        .I3(fch_issu1_inferred_i_148_n_0),
        .I4(fdatx[13]),
        .I5(fdatx[14]),
        .O(fch_issu1_inferred_i_76_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAA80808088)) 
    fch_issu1_inferred_i_77
       (.I0(fch_issu1_inferred_i_71_n_0),
        .I1(fch_issu1_inferred_i_140_n_0),
        .I2(fch_issu1_inferred_i_149_n_0),
        .I3(fch_issu1_inferred_i_150_n_0),
        .I4(fch_issu1_inferred_i_151_n_0),
        .I5(fdatx[15]),
        .O(fch_issu1_inferred_i_77_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF7F7F7F)) 
    fch_issu1_inferred_i_78
       (.I0(fdatx[0]),
        .I1(fdatx[14]),
        .I2(fch_issu1_inferred_i_20_n_0),
        .I3(fch_issu1_inferred_i_119_n_0),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_152_n_0),
        .O(fch_issu1_inferred_i_78_n_0));
  LUT6 #(
    .INIT(64'hFBEBEBEBAAAAAAAA)) 
    fch_issu1_inferred_i_79
       (.I0(fdatx[11]),
        .I1(fdatx[9]),
        .I2(fdatx[8]),
        .I3(fdatx[7]),
        .I4(fdatx[6]),
        .I5(fdatx[10]),
        .O(fch_issu1_inferred_i_79_n_0));
  LUT4 #(
    .INIT(16'hF66F)) 
    fch_issu1_inferred_i_8
       (.I0(fch_issu1_inferred_i_17_n_0),
        .I1(fch_issu1_inferred_i_33_n_0),
        .I2(fch_issu1_inferred_i_15_n_0),
        .I3(fch_issu1_inferred_i_34_n_0),
        .O(fch_issu1_inferred_i_8_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAAEAAAAAA)) 
    fch_issu1_inferred_i_80
       (.I0(fch_issu1_inferred_i_36_n_0),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fch_issu1_inferred_i_153_n_0),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_80_n_0));
  LUT6 #(
    .INIT(64'h00004000FFFFFFFF)) 
    fch_issu1_inferred_i_81
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(fch_issu1_inferred_i_105_n_0),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fch_issu1_inferred_i_37_n_0),
        .O(fch_issu1_inferred_i_81_n_0));
  LUT6 #(
    .INIT(64'hFFDFFFDDFFFFFF00)) 
    fch_issu1_inferred_i_82
       (.I0(fch_issu1_inferred_i_154_n_0),
        .I1(fch_issu1_inferred_i_127_n_0),
        .I2(fdatx[9]),
        .I3(fch_issu1_inferred_i_106_n_0),
        .I4(fdatx[4]),
        .I5(fch_issu1_inferred_i_119_n_0),
        .O(fch_issu1_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFD555)) 
    fch_issu1_inferred_i_83
       (.I0(\nir_id[15]_i_2_n_0 ),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_83_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_84
       (.I0(fdatx[6]),
        .I1(fdatx[7]),
        .O(fch_issu1_inferred_i_84_n_0));
  LUT6 #(
    .INIT(64'hF6F2F6EAF6EAF6EA)) 
    fch_issu1_inferred_i_85
       (.I0(fdatx[11]),
        .I1(fdatx[10]),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(fdatx[6]),
        .I5(fdatx[7]),
        .O(fch_issu1_inferred_i_85_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_86
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .O(fch_issu1_inferred_i_86_n_0));
  LUT6 #(
    .INIT(64'h5555555155555555)) 
    fch_issu1_inferred_i_87
       (.I0(fdatx[12]),
        .I1(\ir0_id_fl[20]_i_7_n_0 ),
        .I2(fdatx[11]),
        .I3(fdatx[13]),
        .I4(fdatx[14]),
        .I5(fch_issu1_inferred_i_155_n_0),
        .O(fch_issu1_inferred_i_87_n_0));
  LUT6 #(
    .INIT(64'h5555555555555545)) 
    fch_issu1_inferred_i_88
       (.I0(fdat[12]),
        .I1(fch_issu1_inferred_i_156_n_0),
        .I2(\nir_id[20]_i_4_n_0 ),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_88_n_0));
  LUT6 #(
    .INIT(64'h00A80000000A02AA)) 
    fch_issu1_inferred_i_89
       (.I0(fch_issu1_inferred_i_157_n_0),
        .I1(\nir_id[14]_i_9_n_0 ),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_89_n_0));
  LUT6 #(
    .INIT(64'h0707000F07070707)) 
    fch_issu1_inferred_i_9
       (.I0(\fch/lir_id_0 [17]),
        .I1(\fch/fadr_1_fl ),
        .I2(fch_issu1_inferred_i_35_n_0),
        .I3(\fch/nir_id [17]),
        .I4(\fch/stat [0]),
        .I5(\fch/stat [1]),
        .O(fch_issu1_inferred_i_9_n_0));
  LUT4 #(
    .INIT(16'h0440)) 
    fch_issu1_inferred_i_90
       (.I0(fdatx[13]),
        .I1(fdatx[14]),
        .I2(fdatx[12]),
        .I3(fdatx[11]),
        .O(fch_issu1_inferred_i_90_n_0));
  LUT6 #(
    .INIT(64'hFBBFBBBFAAAAAAAA)) 
    fch_issu1_inferred_i_91
       (.I0(\ir0_id_fl[20]_i_4_n_0 ),
        .I1(fch_issu1_inferred_i_158_n_0),
        .I2(fdatx[6]),
        .I3(fch_issu1_inferred_i_159_n_0),
        .I4(fdatx[3]),
        .I5(fch_issu1_inferred_i_160_n_0),
        .O(fch_issu1_inferred_i_91_n_0));
  LUT6 #(
    .INIT(64'h3FFE3FFF3FFF3FFF)) 
    fch_issu1_inferred_i_92
       (.I0(fch_issu1_inferred_i_161_n_0),
        .I1(fdatx[12]),
        .I2(fdatx[7]),
        .I3(fdatx[9]),
        .I4(\ir0_id_fl[20]_i_8_n_0 ),
        .I5(fch_issu1_inferred_i_162_n_0),
        .O(fch_issu1_inferred_i_92_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_93
       (.I0(fdatx[8]),
        .I1(fdatx[6]),
        .O(fch_issu1_inferred_i_93_n_0));
  LUT5 #(
    .INIT(32'h44444044)) 
    fch_issu1_inferred_i_94
       (.I0(fch_issu1_inferred_i_113_n_0),
        .I1(\nir_id[15]_i_2_n_0 ),
        .I2(fch_issu1_inferred_i_114_n_0),
        .I3(fdat[11]),
        .I4(fdat[10]),
        .O(fch_issu1_inferred_i_94_n_0));
  LUT6 #(
    .INIT(64'h5CCC0CCC5CCCCCCC)) 
    fch_issu1_inferred_i_95
       (.I0(fch_issu1_inferred_i_163_n_0),
        .I1(fdat[4]),
        .I2(fdat[11]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .I5(\nir_id[14]_i_12_n_0 ),
        .O(fch_issu1_inferred_i_95_n_0));
  LUT6 #(
    .INIT(64'h000000004477C0FF)) 
    fch_issu1_inferred_i_96
       (.I0(fch_issu1_inferred_i_164_n_0),
        .I1(fch_issu1_inferred_i_119_n_0),
        .I2(fch_issu1_inferred_i_165_n_0),
        .I3(fdatx[4]),
        .I4(fdatx[9]),
        .I5(fch_issu1_inferred_i_118_n_0),
        .O(fch_issu1_inferred_i_96_n_0));
  LUT6 #(
    .INIT(64'h000000007FDF57FF)) 
    fch_issu1_inferred_i_97
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fdat[11]),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_97_n_0));
  LUT6 #(
    .INIT(64'h0A2A000A2000000A)) 
    fch_issu1_inferred_i_98
       (.I0(fdat[8]),
        .I1(fdat[3]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_98_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_99
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_99_n_0));
  LUT6 #(
    .INIT(64'h8B8B8B8B888B8B8B)) 
    fch_leir_hir_i_1
       (.I0(fch_leir_hir_i_2_n_0),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(\rgf/pcnt/pc [1]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(\fch/stat [2]),
        .O(\fch/fctl/fch_leir_hir_t ));
  LUT5 #(
    .INIT(32'h00002134)) 
    fch_leir_hir_i_2
       (.I0(\fch/stat [2]),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [1]),
        .I3(\fch/fch_issu1_ir ),
        .I4(\fadr[15]_INST_0_i_4_n_0 ),
        .O(fch_leir_hir_i_2_n_0));
  LUT5 #(
    .INIT(32'h0000BF00)) 
    fch_leir_lir_i_1
       (.I0(\fch/stat [2]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\rgf/pcnt/pc [1]),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\fch/fctl/fch_leir_lir_t ));
  LUT5 #(
    .INIT(32'h00004004)) 
    fch_leir_nir_i_1
       (.I0(\fch/stat [0]),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(\fch/stat [1]),
        .I3(fch_leir_nir_i_2_n_0),
        .I4(\fadr[15]_INST_0_i_4_n_0 ),
        .O(\fch/fctl/fch_leir_nir_t ));
  LUT4 #(
    .INIT(16'h00E2)) 
    fch_leir_nir_i_2
       (.I0(\fch/fch_issu1_fl ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_issu1 ),
        .I3(\fch/stat [2]),
        .O(fch_leir_nir_i_2_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    fch_pc_nx2_carry_i_1
       (.I0(\rgf/pcnt/pc [1]),
        .O(fch_pc_nx2_carry_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    fch_pc_nx4_carry_i_1
       (.I0(\rgf/pcnt/pc [2]),
        .O(fch_pc_nx4_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_term_fl_i_1
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .O(fch_term));
  LUT4 #(
    .INIT(16'hAAAE)) 
    \grn[15]_i_1 
       (.I0(\rgf/bank02/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hEAAA)) 
    \grn[15]_i_1__0 
       (.I0(\rgf/bank13/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__0_n_0 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1__1 
       (.I0(\rgf/bank13/grn05/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0F0F1)) 
    \grn[15]_i_1__10 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn03/grn1 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__10_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__11 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn22/grn1 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__11_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__12 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn02/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__12_n_0 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__13 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank13/grn22/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__13_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__14 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/bank02/grn02/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__15 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn21/grn1 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__16 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn01/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__17 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn21/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__18 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn01/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__19 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn26/grn1 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__19_n_0 ));
  LUT4 #(
    .INIT(16'hAAEA)) 
    \grn[15]_i_1__2 
       (.I0(\rgf/bank02/grn25/grn1 ),
        .I1(\rgf/c0bus_sel_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF40FF00)) 
    \grn[15]_i_1__20 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn06/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hFF40FF00FF00FF00)) 
    \grn[15]_i_1__21 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank13/grn26/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF40)) 
    \grn[15]_i_1__22 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/bank02/grn06/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__23 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn24/grn1 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF04FF00)) 
    \grn[15]_i_1__24 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn04/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hFF04FF00FF00FF00)) 
    \grn[15]_i_1__25 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank13/grn24/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF04)) 
    \grn[15]_i_1__26 
       (.I0(\grn[15]_i_3__1_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/bank02/grn04/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF01FF00)) 
    \grn[15]_i_1__27 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank13/grn00/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF01FF00)) 
    \grn[15]_i_1__28 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank02/grn20/grn1 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hFF01FF00FF00FF00)) 
    \grn[15]_i_1__29 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank13/grn20/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__29_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn27/grn1 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF01)) 
    \grn[15]_i_1__30 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\grn[15]_i_5__0_n_0 ),
        .I3(\rgf/bank02/grn00/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__30_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF02FF00)) 
    \grn[15]_i_1__4 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn07/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__4_n_0 ));
  LUT6 #(
    .INIT(64'hFF02FF00FF00FF00)) 
    \grn[15]_i_1__5 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank13/grn27/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__5_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF00FF00FF02)) 
    \grn[15]_i_1__6 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .I3(\rgf/bank02/grn07/grn1 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__6_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__7 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn23/grn1 ),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/sreg/sr [0]),
        .O(\grn[15]_i_1__7_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0F1F0)) 
    \grn[15]_i_1__8 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn03/grn1 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__8_n_0 ));
  LUT5 #(
    .INIT(32'hF1F0F0F0)) 
    \grn[15]_i_1__9 
       (.I0(\grn[15]_i_5__0_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn23/grn1 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__9_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .O(\grn[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_3__0 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(ctl_selc0_rn),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_rn_wb [1]),
        .O(\rgf/rctl/p_0_in [1]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_3__1 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .O(\grn[15]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__10 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__11 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn04/grn1 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \grn[15]_i_3__12 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h0100000000000000)) 
    \grn[15]_i_3__13 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__14 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn24/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__15 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn26/grn1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \grn[15]_i_3__16 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn06/grn1 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \grn[15]_i_3__17 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn20/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__18 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\rgf/bank02/grn20/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__19 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn00/grn1 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \grn[15]_i_3__2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__20 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__21 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn03/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__22 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\rgf/bank02/grn23/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__23 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank02/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__24 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank13/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__25 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0000010000000000)) 
    \grn[15]_i_3__26 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__27 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank13/grn21/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__28 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank13/grn22/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__29 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\rgf/bank02/grn01/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_3__30 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [0]),
        .I5(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/bank02/grn02/grn1 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \grn[15]_i_3__4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\rgf/bank02/grn27/grn1 ));
  LUT6 #(
    .INIT(64'h1B1F5F1FFFFFFFFF)) 
    \grn[15]_i_3__5 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\rgf_selc0_wb[0]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_wb [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\grn[15]_i_3__5_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__6 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/sreg/sr [1]),
        .O(\rgf/bank02/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \grn[15]_i_3__7 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn05/grn1 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \grn[15]_i_3__8 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/grn25/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_3__9 
       (.I0(\grn[15]_i_7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank02/grn05/grn1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4 
       (.I0(\grn[15]_i_3__5_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/rctl/p_0_in [2]),
        .O(\rgf/c0bus_sel_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__0 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\rgf_selc0_rn_wb[0]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_rn_wb [0]),
        .O(\rgf/rctl/p_0_in [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_4__1 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\rgf_selc0_rn_wb[2]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_rn_wb [2]),
        .O(\rgf/rctl/p_0_in [2]));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \grn[15]_i_4__2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank02/grn07/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \grn[15]_i_4__3 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank02/grn03/grn1 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_5 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(ctl_selc0),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_wb [1]),
        .O(\rgf/rctl/p_0_in [4]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_5__0 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_3__5_n_0 ),
        .O(\grn[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \grn[15]_i_5__1 
       (.I0(\rgf/rctl/rgf_selc1_rn [0]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn04/grn1 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \grn[15]_i_6 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\grn[15]_i_7_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/sreg/sr [0]),
        .O(\rgf/bank02/grn00/grn1 ));
  LUT6 #(
    .INIT(64'h55FF55FF757FFFFF)) 
    \grn[15]_i_7 
       (.I0(\rgf/rctl/rgf_selc1 [1]),
        .I1(\rgf/rctl/rgf_selc1_wb [0]),
        .I2(\rgf/rctl/rgf_selc1_stat ),
        .I3(\rgf_selc1_wb[0]_i_1_n_0 ),
        .I4(fch_term),
        .I5(fch_wrbufn1),
        .O(\grn[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \grn[15]_i_8 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(ctl_selc1),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_wb [1]),
        .O(\rgf/rctl/rgf_selc1 [1]));
  LUT4 #(
    .INIT(16'h8880)) 
    \ir0_id_fl[20]_i_1 
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(\fch/rst_n_fl ),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/ir0_id_fl [20]),
        .O(\fch/p_0_in ));
  LUT6 #(
    .INIT(64'hF3FFC0FFD1FFD1FF)) 
    \ir0_id_fl[20]_i_2 
       (.I0(\ir0_id_fl[20]_i_3_n_0 ),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(\fch/nir_id [20]),
        .I3(ir0_inferred_i_33_n_0),
        .I4(\nir_id[20]_i_1_n_0 ),
        .I5(\fch/fadr_1_fl ),
        .O(\ir0_id_fl[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hABAAABABABABABAB)) 
    \ir0_id_fl[20]_i_3 
       (.I0(fdatx[15]),
        .I1(\ir0_id_fl[20]_i_4_n_0 ),
        .I2(\ir0_id_fl[20]_i_5_n_0 ),
        .I3(\ir0_id_fl[20]_i_6_n_0 ),
        .I4(fdatx[12]),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[20]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0FFE)) 
    \ir0_id_fl[20]_i_4 
       (.I0(fdatx[12]),
        .I1(fdatx[11]),
        .I2(fdatx[13]),
        .I3(fdatx[14]),
        .O(\ir0_id_fl[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0002002202000020)) 
    \ir0_id_fl[20]_i_5 
       (.I0(\ir0_id_fl[20]_i_7_n_0 ),
        .I1(fdatx[13]),
        .I2(fdatx[0]),
        .I3(fdatx[3]),
        .I4(fdatx[2]),
        .I5(fdatx[1]),
        .O(\ir0_id_fl[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hA2AABBBBFFFFAAAA)) 
    \ir0_id_fl[20]_i_6 
       (.I0(fdatx[9]),
        .I1(fdatx[7]),
        .I2(fdatx[6]),
        .I3(\ir0_id_fl[20]_i_8_n_0 ),
        .I4(fdatx[8]),
        .I5(fdatx[11]),
        .O(\ir0_id_fl[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \ir0_id_fl[20]_i_7 
       (.I0(\ir0_id_fl[20]_i_8_n_0 ),
        .I1(fdatx[8]),
        .I2(fdatx[9]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[20]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[20]_i_8 
       (.I0(fdatx[5]),
        .I1(fdatx[4]),
        .O(\ir0_id_fl[20]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h8880)) 
    \ir0_id_fl[21]_i_1 
       (.I0(\ir0_id_fl[21]_i_2_n_0 ),
        .I1(\fch/rst_n_fl ),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/ir0_id_fl [21]),
        .O(\fch/ir0_id ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \ir0_id_fl[21]_i_10 
       (.I0(\ir0_id_fl[20]_i_8_n_0 ),
        .I1(fdatx[3]),
        .I2(fdatx[2]),
        .I3(fch_issu1_inferred_i_104_n_0),
        .I4(fdatx[10]),
        .I5(fdatx[11]),
        .O(\ir0_id_fl[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF3FFC0FFD1FFD1FF)) 
    \ir0_id_fl[21]_i_2 
       (.I0(\ir0_id_fl[21]_i_3_n_0 ),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(\fch/nir_id [21]),
        .I3(ir0_inferred_i_33_n_0),
        .I4(\fch/lir_id_0 [21]),
        .I5(\fch/fadr_1_fl ),
        .O(\ir0_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF5554)) 
    \ir0_id_fl[21]_i_3 
       (.I0(\ir0_id_fl[21]_i_4_n_0 ),
        .I1(\ir0_id_fl[21]_i_5_n_0 ),
        .I2(fdatx[9]),
        .I3(fdatx[8]),
        .I4(\ir0_id_fl[21]_i_6_n_0 ),
        .I5(fdatx[15]),
        .O(\ir0_id_fl[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F6000000)) 
    \ir0_id_fl[21]_i_4 
       (.I0(fdatx[10]),
        .I1(fdatx[11]),
        .I2(\ir0_id_fl[21]_i_7_n_0 ),
        .I3(\ir0_id_fl[21]_i_8_n_0 ),
        .I4(fdatx[13]),
        .I5(\ir0_id_fl[21]_i_9_n_0 ),
        .O(\ir0_id_fl[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3FFFFFFFFFFFFF55)) 
    \ir0_id_fl[21]_i_5 
       (.I0(\ir0_id_fl[21]_i_10_n_0 ),
        .I1(fch_issu1_inferred_i_119_n_0),
        .I2(fdatx[7]),
        .I3(fdatx[12]),
        .I4(fdatx[13]),
        .I5(fdatx[14]),
        .O(\ir0_id_fl[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ir0_id_fl[21]_i_6 
       (.I0(fdatx[1]),
        .I1(fdatx[0]),
        .I2(fdatx[8]),
        .I3(fdatx[10]),
        .I4(fdatx[3]),
        .I5(fdatx[5]),
        .O(\ir0_id_fl[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCC10000000000000)) 
    \ir0_id_fl[21]_i_7 
       (.I0(fdatx[4]),
        .I1(fdatx[5]),
        .I2(fdatx[3]),
        .I3(fdatx[6]),
        .I4(fdatx[7]),
        .I5(fdatx[10]),
        .O(\ir0_id_fl[21]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ir0_id_fl[21]_i_8 
       (.I0(fdatx[12]),
        .I1(fdatx[14]),
        .O(\ir0_id_fl[21]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ir0_id_fl[21]_i_9 
       (.I0(fdatx[8]),
        .I1(fdatx[9]),
        .O(\ir0_id_fl[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_1
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [15]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_17_n_0),
        .O(\fch/ir0 [15]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_10
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [6]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_26_n_0),
        .O(\fch/ir0 [6]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_11
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [5]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_27_n_0),
        .O(\fch/ir0 [5]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_12
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [4]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_28_n_0),
        .O(\fch/ir0 [4]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_13
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [3]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_29_n_0),
        .O(\fch/ir0 [3]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_14
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [2]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_30_n_0),
        .O(\fch/ir0 [2]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_15
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [1]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_31_n_0),
        .O(\fch/ir0 [1]));
  LUT5 #(
    .INIT(32'h88880080)) 
    ir0_inferred_i_16
       (.I0(ir0_inferred_i_32_n_0),
        .I1(\fch/rst_n_fl ),
        .I2(\fch/ir0_fl [0]),
        .I3(\fch/ctl_fetch0_fl ),
        .I4(\fch/fch_term_fl ),
        .O(\fch/ir0 [0]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_17
       (.I0(\fch/nir [15]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[15]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[15]),
        .O(ir0_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_18
       (.I0(\fch/nir [14]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[14]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[14]),
        .O(ir0_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_19
       (.I0(\fch/nir [13]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[13]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[13]),
        .O(ir0_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_2
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [14]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_18_n_0),
        .O(\fch/ir0 [14]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_20
       (.I0(\fch/nir [12]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[12]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[12]),
        .O(ir0_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_21
       (.I0(\fch/nir [11]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[11]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[11]),
        .O(ir0_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_22
       (.I0(\fch/nir [10]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[10]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[10]),
        .O(ir0_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_23
       (.I0(\fch/nir [9]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[9]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[9]),
        .O(ir0_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_24
       (.I0(\fch/nir [8]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[8]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[8]),
        .O(ir0_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_25
       (.I0(\fch/nir [7]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[7]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[7]),
        .O(ir0_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_26
       (.I0(\fch/nir [6]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[6]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[6]),
        .O(ir0_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_27
       (.I0(\fch/nir [5]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[5]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[5]),
        .O(ir0_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_28
       (.I0(\fch/nir [4]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[4]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[4]),
        .O(ir0_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_29
       (.I0(\fch/nir [3]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[3]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[3]),
        .O(ir0_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_3
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [13]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_19_n_0),
        .O(\fch/ir0 [13]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_30
       (.I0(\fch/nir [2]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[2]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[2]),
        .O(ir0_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_31
       (.I0(\fch/nir [1]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[1]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdatx[1]),
        .O(ir0_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hFECE3202FFFFFFFF)) 
    ir0_inferred_i_32
       (.I0(fdatx[0]),
        .I1(fch_issu1_inferred_i_20_n_0),
        .I2(\fch/fadr_1_fl ),
        .I3(fdat[0]),
        .I4(\fch/nir [0]),
        .I5(ir0_inferred_i_33_n_0),
        .O(ir0_inferred_i_32_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ir0_inferred_i_33
       (.I0(\fch/fch_term_fl ),
        .I1(\fch/fch_irq_req_fl ),
        .O(ir0_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_4
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [12]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_20_n_0),
        .O(\fch/ir0 [12]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_5
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [11]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_21_n_0),
        .O(\fch/ir0 [11]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_6
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [10]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_22_n_0),
        .O(\fch/ir0 [10]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_7
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [9]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_23_n_0),
        .O(\fch/ir0 [9]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_8
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [8]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_24_n_0),
        .O(\fch/ir0 [8]));
  LUT6 #(
    .INIT(64'h0020AA2000200020)) 
    ir0_inferred_i_9
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ctl_fetch0_fl ),
        .I2(\fch/ir0_fl [7]),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(ir0_inferred_i_25_n_0),
        .O(\fch/ir0 [7]));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[20]_i_1 
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir1_id_fl [20]),
        .I2(\fch/fch_term_fl ),
        .I3(\ir1_id_fl[20]_i_2_n_0 ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(\fch/fch_issu1 ),
        .O(fch_wrbufn1));
  LUT5 #(
    .INIT(32'hCACCFAFF)) 
    \ir1_id_fl[20]_i_2 
       (.I0(\ir0_id_fl[20]_i_3_n_0 ),
        .I1(\fch/fadr_1_fl ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(\nir_id[20]_i_1_n_0 ),
        .O(\ir1_id_fl[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[21]_i_1 
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir1_id_fl [21]),
        .I2(\fch/fch_term_fl ),
        .I3(\ir1_id_fl[21]_i_2_n_0 ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(\fch/fch_issu1 ),
        .O(fch_memacc1));
  LUT5 #(
    .INIT(32'hCACCFAFF)) 
    \ir1_id_fl[21]_i_2 
       (.I0(\ir0_id_fl[21]_i_3_n_0 ),
        .I1(\fch/fadr_1_fl ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(\fch/lir_id_0 [21]),
        .O(\ir1_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_1
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_18_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [15]),
        .O(\fch/ir1 [15]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_10
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_27_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [6]),
        .O(\fch/ir1 [6]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_11
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_28_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [5]),
        .O(\fch/ir1 [5]));
  LUT6 #(
    .INIT(64'h808080AA80808080)) 
    ir1_inferred_i_12
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_29_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [4]),
        .O(\fch/ir1 [4]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_13
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_30_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [3]),
        .O(\fch/ir1 [3]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_14
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_31_n_0),
        .I2(\fch/ctl_fetch1_fl ),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/ir1_fl [2]),
        .O(\fch/ir1 [2]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_15
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_32_n_0),
        .I2(\fch/ctl_fetch1_fl ),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/ir1_fl [1]),
        .O(\fch/ir1 [1]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_16
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_33_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [0]),
        .O(\fch/ir1 [0]));
  LUT3 #(
    .INIT(8'h20)) 
    ir1_inferred_i_17
       (.I0(\fch/fch_issu1 ),
        .I1(\fch/fch_irq_req_fl ),
        .I2(\fch/fch_term_fl ),
        .O(ir1_inferred_i_17_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_18
       (.I0(fdatx[15]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[15]),
        .O(ir1_inferred_i_18_n_0));
  LUT5 #(
    .INIT(32'hF355F3F3)) 
    ir1_inferred_i_19
       (.I0(fdatx[14]),
        .I1(fdat[14]),
        .I2(\fch/fadr_1_fl ),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .O(ir1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_2
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_19_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [14]),
        .O(\fch/ir1 [14]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_20
       (.I0(fdatx[13]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[13]),
        .O(ir1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_21
       (.I0(fdatx[12]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[12]),
        .O(ir1_inferred_i_21_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_22
       (.I0(fdatx[11]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[11]),
        .O(ir1_inferred_i_22_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_23
       (.I0(fdatx[10]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[10]),
        .O(ir1_inferred_i_23_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_24
       (.I0(fdatx[9]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[9]),
        .O(ir1_inferred_i_24_n_0));
  LUT5 #(
    .INIT(32'hBBBB0FBB)) 
    ir1_inferred_i_25
       (.I0(\fch/fadr_1_fl ),
        .I1(fdat[8]),
        .I2(fdatx[8]),
        .I3(\fch/stat [1]),
        .I4(\fch/stat [0]),
        .O(ir1_inferred_i_25_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_26
       (.I0(fdatx[7]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[7]),
        .O(ir1_inferred_i_26_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_27
       (.I0(fdatx[6]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[6]),
        .O(ir1_inferred_i_27_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_28
       (.I0(fdatx[5]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[5]),
        .O(ir1_inferred_i_28_n_0));
  LUT5 #(
    .INIT(32'h0808FB08)) 
    ir1_inferred_i_29
       (.I0(fdatx[4]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[4]),
        .I4(\fch/fadr_1_fl ),
        .O(ir1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_3
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_20_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [13]),
        .O(\fch/ir1 [13]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_30
       (.I0(fdatx[3]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[3]),
        .O(ir1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h4C4440440C000000)) 
    ir1_inferred_i_31
       (.I0(\fch/fadr_1_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(fdatx[2]),
        .I5(fdat[2]),
        .O(ir1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h44C0444400C00000)) 
    ir1_inferred_i_32
       (.I0(\fch/fadr_1_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(fdatx[1]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fdat[1]),
        .O(ir1_inferred_i_32_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_33
       (.I0(fdatx[0]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[0]),
        .O(ir1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_4
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_21_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [12]),
        .O(\fch/ir1 [12]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_5
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_22_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [11]),
        .O(\fch/ir1 [11]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_6
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_23_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [10]),
        .O(\fch/ir1 [10]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_7
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_24_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [9]),
        .O(\fch/ir1 [9]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_8
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_25_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [8]),
        .O(\fch/ir1 [8]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_9
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_26_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [7]),
        .O(\fch/ir1 [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [0]),
        .O(\rgf/ivec/p_1_in [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [10]),
        .O(\rgf/ivec/p_1_in [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [11]),
        .O(\rgf/ivec/p_1_in [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [12]),
        .O(\rgf/ivec/p_1_in [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [13]),
        .O(\rgf/ivec/p_1_in [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [14]),
        .O(\rgf/ivec/p_1_in [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [15]),
        .O(\rgf/ivec/p_1_in [15]));
  LUT4 #(
    .INIT(16'h0008)) 
    \iv[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_3 
       (.I0(\grn[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [1]),
        .O(\rgf/ivec/p_1_in [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [2]),
        .O(\rgf/ivec/p_1_in [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [3]),
        .O(\rgf/ivec/p_1_in [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [4]),
        .O(\rgf/ivec/p_1_in [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [5]),
        .O(\rgf/ivec/p_1_in [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [6]),
        .O(\rgf/ivec/p_1_in [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [7]),
        .O(\rgf/ivec/p_1_in [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [8]),
        .O(\rgf/ivec/p_1_in [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [9]),
        .O(\rgf/ivec/p_1_in [9]));
  FDRE \mem/bctl/ctl/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mem/bctl/ctl/stat_nx [0]),
        .Q(\mem/bctl/ctl/p_0_in [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \mem/bctl/ctl/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mem/bctl/ctl/stat_nx [1]),
        .Q(\mem/bctl/ctl/p_0_in [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \mem/bctl/fch_term_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(\mem/bctl/fch_term_fl ),
        .R(\<const0> ));
  FDRE \mem/bctl/read_cyc_reg[0] 
       (.C(clk),
        .CE(brdy),
        .D(badr[0]),
        .Q(\mem/read_cyc [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \mem/bctl/read_cyc_reg[1] 
       (.C(clk),
        .CE(brdy),
        .D(bcmd[2]),
        .Q(\mem/read_cyc [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \mem/bctl/read_cyc_reg[2] 
       (.C(clk),
        .CE(brdy),
        .D(bcmd[0]),
        .Q(\mem/read_cyc [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \mem/bctl/read_cyc_reg[3] 
       (.C(clk),
        .CE(brdy),
        .D(\mem/mem_accslot ),
        .Q(\mem/read_cyc [3]),
        .R(\rgf/treg/p_0_in ));
  LUT6 #(
    .INIT(64'hCC70FFFFCC700000)) 
    \nir_id[12]_i_1 
       (.I0(fdat[11]),
        .I1(fdat[12]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(fdat[15]),
        .I5(\nir_id[12]_i_2_n_0 ),
        .O(\fch/lir_id_0 [12]));
  LUT6 #(
    .INIT(64'hBABABABABABBBABA)) 
    \nir_id[12]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[12]_i_3_n_0 ),
        .I2(\nir_id[14]_i_10_n_0 ),
        .I3(\nir_id[12]_i_4_n_0 ),
        .I4(fdat[0]),
        .I5(fdat[9]),
        .O(\nir_id[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h75770000FFFFFFFF)) 
    \nir_id[12]_i_3 
       (.I0(fdat[10]),
        .I1(\nir_id[13]_i_4_n_0 ),
        .I2(fdat[8]),
        .I3(fdat[0]),
        .I4(\nir_id[14]_i_8_n_0 ),
        .I5(fdat[14]),
        .O(\nir_id[12]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[12]_i_4 
       (.I0(fdat[8]),
        .I1(fdat[10]),
        .O(\nir_id[12]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[13]_i_1 
       (.I0(\nir_id[13]_i_2_n_0 ),
        .O(\fch/lir_id_0 [13]));
  LUT6 #(
    .INIT(64'h558F558F0000F000)) 
    \nir_id[13]_i_2 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(\nir_id[13]_i_3_n_0 ),
        .I5(fdat[15]),
        .O(\nir_id[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AE00FFFF)) 
    \nir_id[13]_i_3 
       (.I0(\nir_id[13]_i_4_n_0 ),
        .I1(fdat[1]),
        .I2(fdat[8]),
        .I3(fdat[10]),
        .I4(\nir_id[14]_i_8_n_0 ),
        .I5(\nir_id[13]_i_5_n_0 ),
        .O(\nir_id[13]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \nir_id[13]_i_4 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .O(\nir_id[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h888A0AAA8A8A0AAA)) 
    \nir_id[13]_i_5 
       (.I0(\nir_id[24]_i_13_n_0 ),
        .I1(\nir_id[13]_i_6_n_0 ),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[10]),
        .I5(fdat[1]),
        .O(\nir_id[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0005555010000005)) 
    \nir_id[13]_i_6 
       (.I0(\nir_id[13]_i_7_n_0 ),
        .I1(fdat[3]),
        .I2(fdat[6]),
        .I3(fdat[4]),
        .I4(fdat[5]),
        .I5(fdat[7]),
        .O(\nir_id[13]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[13]_i_7 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(\nir_id[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7477747474747474)) 
    \nir_id[14]_i_1 
       (.I0(\nir_id[14]_i_2_n_0 ),
        .I1(fdat[15]),
        .I2(\nir_id[14]_i_3_n_0 ),
        .I3(\nir_id[14]_i_4_n_0 ),
        .I4(fdat[14]),
        .I5(\nir_id[14]_i_5_n_0 ),
        .O(\fch/lir_id_0 [14]));
  LUT6 #(
    .INIT(64'hB080FFFFFFFFFFFF)) 
    \nir_id[14]_i_10 
       (.I0(\nir_id[14]_i_13_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[14]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[14]_i_11 
       (.I0(fdat[3]),
        .I1(fdat[2]),
        .O(\nir_id[14]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \nir_id[14]_i_12 
       (.I0(fdat[6]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .O(\nir_id[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h55D415D6FFFFFFFF)) 
    \nir_id[14]_i_13 
       (.I0(fdat[7]),
        .I1(fdat[5]),
        .I2(fdat[4]),
        .I3(fdat[6]),
        .I4(fdat[3]),
        .I5(fdat[8]),
        .O(\nir_id[14]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h5B1B)) 
    \nir_id[14]_i_2 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(\nir_id[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0FFF0FF70FFF0FFF)) 
    \nir_id[14]_i_3 
       (.I0(\nir_id[14]_i_6_n_0 ),
        .I1(\nir_id[20]_i_5_n_0 ),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .I4(fdat[12]),
        .I5(\nir_id[14]_i_7_n_0 ),
        .O(\nir_id[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A20002AAAAAAAA)) 
    \nir_id[14]_i_4 
       (.I0(\nir_id[14]_i_8_n_0 ),
        .I1(fdat[2]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(\nir_id[14]_i_9_n_0 ),
        .I5(fdat[10]),
        .O(\nir_id[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABAAABABAAAAA)) 
    \nir_id[14]_i_5 
       (.I0(\nir_id[14]_i_10_n_0 ),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[2]),
        .I4(fdat[7]),
        .I5(fdat[8]),
        .O(\nir_id[14]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[14]_i_6 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(\nir_id[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0008000800080000)) 
    \nir_id[14]_i_7 
       (.I0(\nir_id[14]_i_11_n_0 ),
        .I1(\nir_id[19]_i_5_n_0 ),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .I4(fdat[0]),
        .I5(fdat[1]),
        .O(\nir_id[14]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00EC0000)) 
    \nir_id[14]_i_8 
       (.I0(\nir_id[14]_i_12_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[11]),
        .I4(fdat[12]),
        .O(\nir_id[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[14]_i_9 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDFFDFFFFFFFF)) 
    \nir_id[15]_i_1 
       (.I0(fdat[10]),
        .I1(fdat[9]),
        .I2(fdat[11]),
        .I3(fdat[8]),
        .I4(fdat[15]),
        .I5(\nir_id[15]_i_2_n_0 ),
        .O(\fch/lir_id_0 [15]));
  LUT3 #(
    .INIT(8'h80)) 
    \nir_id[15]_i_2 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .O(\nir_id[15]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hEEE0)) 
    \nir_id[16]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(fdat[8]),
        .I2(\nir_id[16]_i_2_n_0 ),
        .I3(\nir_id[19]_i_3_n_0 ),
        .O(\fch/lir_id_0 [16]));
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEA0000)) 
    \nir_id[16]_i_2 
       (.I0(\nir_id[19]_i_9_n_0 ),
        .I1(fdat[0]),
        .I2(fdat[9]),
        .I3(\nir_id[16]_i_3_n_0 ),
        .I4(\nir_id[17]_i_2_n_0 ),
        .I5(fdat[3]),
        .O(\nir_id[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h8888888088888888)) 
    \nir_id[16]_i_3 
       (.I0(\nir_id[19]_i_11_n_0 ),
        .I1(fdat[9]),
        .I2(\nir_id[19]_i_12_n_0 ),
        .I3(fdat[3]),
        .I4(fdat[7]),
        .I5(fdat[8]),
        .O(\nir_id[16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hEEEE0E00EEEEEEE0)) 
    \nir_id[17]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(fdat[9]),
        .I2(\nir_id[17]_i_2_n_0 ),
        .I3(fdat[4]),
        .I4(\nir_id[19]_i_3_n_0 ),
        .I5(\nir_id[17]_i_3_n_0 ),
        .O(\fch/lir_id_0 [17]));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[17]_i_2 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00F100F1000000FF)) 
    \nir_id[17]_i_3 
       (.I0(\nir_id[19]_i_11_n_0 ),
        .I1(fdat[1]),
        .I2(\nir_id[17]_i_4_n_0 ),
        .I3(\nir_id[19]_i_9_n_0 ),
        .I4(fdat[4]),
        .I5(fdat[9]),
        .O(\nir_id[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h888A000088880000)) 
    \nir_id[17]_i_4 
       (.I0(\nir_id[17]_i_5_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[3]),
        .I3(fdat[1]),
        .I4(fdat[8]),
        .I5(\nir_id[20]_i_5_n_0 ),
        .O(\nir_id[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000F0F00080F0F)) 
    \nir_id[17]_i_5 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[1]),
        .I4(fdat[6]),
        .I5(fdat[3]),
        .O(\nir_id[17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEE2E00EEEEEEC0)) 
    \nir_id[18]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[5]),
        .I4(\nir_id[19]_i_3_n_0 ),
        .I5(\nir_id[18]_i_2_n_0 ),
        .O(\fch/lir_id_0 [18]));
  LUT6 #(
    .INIT(64'h00F100F1000000FF)) 
    \nir_id[18]_i_2 
       (.I0(\nir_id[19]_i_11_n_0 ),
        .I1(fdat[2]),
        .I2(\nir_id[18]_i_3_n_0 ),
        .I3(\nir_id[19]_i_9_n_0 ),
        .I4(fdat[5]),
        .I5(fdat[9]),
        .O(\nir_id[18]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h888A000088880000)) 
    \nir_id[18]_i_3 
       (.I0(\nir_id[18]_i_4_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[3]),
        .I3(fdat[2]),
        .I4(fdat[8]),
        .I5(\nir_id[20]_i_5_n_0 ),
        .O(\nir_id[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000000080F0F0F0F)) 
    \nir_id[18]_i_4 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[6]),
        .O(\nir_id[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hE0EEE0E0EEEEEEEE)) 
    \nir_id[19]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .I1(\nir_id[24]_i_4_n_0 ),
        .I2(\nir_id[19]_i_3_n_0 ),
        .I3(\nir_id[19]_i_4_n_0 ),
        .I4(\nir_id[19]_i_5_n_0 ),
        .I5(\nir_id[19]_i_6_n_0 ),
        .O(\fch/lir_id_0 [19]));
  LUT5 #(
    .INIT(32'h0002FFFF)) 
    \nir_id[19]_i_10 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[3]),
        .I3(\nir_id[19]_i_12_n_0 ),
        .I4(fdat[9]),
        .O(\nir_id[19]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h4FFFFFFF)) 
    \nir_id[19]_i_11 
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[8]),
        .I4(fdat[6]),
        .O(\nir_id[19]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \nir_id[19]_i_12 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .I2(fdat[6]),
        .O(\nir_id[19]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hDD557555)) 
    \nir_id[19]_i_2 
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .I2(fdat[11]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .O(\nir_id[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \nir_id[19]_i_3 
       (.I0(\nir_id[19]_i_7_n_0 ),
        .I1(\nir_id[19]_i_8_n_0 ),
        .I2(fdat[15]),
        .I3(fdat[12]),
        .I4(fdat[14]),
        .I5(fdat[13]),
        .O(\nir_id[19]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFDFF)) 
    \nir_id[19]_i_4 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .I2(fdat[10]),
        .I3(fdat[11]),
        .O(\nir_id[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[19]_i_5 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .O(\nir_id[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44454545FFFFFFFF)) 
    \nir_id[19]_i_6 
       (.I0(\nir_id[19]_i_9_n_0 ),
        .I1(\nir_id[19]_i_10_n_0 ),
        .I2(\nir_id[19]_i_11_n_0 ),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(\nir_id[17]_i_2_n_0 ),
        .O(\nir_id[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2200222202220000)) 
    \nir_id[19]_i_7 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(\nir_id[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000DFD000000000)) 
    \nir_id[19]_i_8 
       (.I0(fdat[11]),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(fdat[7]),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(\nir_id[19]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \nir_id[19]_i_9 
       (.I0(fdat[9]),
        .I1(fdat[8]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .O(\nir_id[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5455545454545454)) 
    \nir_id[20]_i_1 
       (.I0(fdat[15]),
        .I1(\nir_id[20]_i_2_n_0 ),
        .I2(\nir_id[24]_i_8_n_0 ),
        .I3(\nir_id[20]_i_3_n_0 ),
        .I4(fdat[12]),
        .I5(fdat[10]),
        .O(\nir_id[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000C04080008)) 
    \nir_id[20]_i_2 
       (.I0(fdat[1]),
        .I1(\nir_id[20]_i_4_n_0 ),
        .I2(fdat[13]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[0]),
        .O(\nir_id[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hA2AABBBBFFFFAAAA)) 
    \nir_id[20]_i_3 
       (.I0(fdat[9]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(\nir_id[20]_i_5_n_0 ),
        .I4(fdat[8]),
        .I5(fdat[11]),
        .O(\nir_id[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \nir_id[20]_i_4 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .I2(\nir_id[20]_i_5_n_0 ),
        .I3(fdat[10]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[20]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[20]_i_5 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(\nir_id[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAAA2)) 
    \nir_id[21]_i_1 
       (.I0(\nir_id[21]_i_2_n_0 ),
        .I1(\nir_id[21]_i_3_n_0 ),
        .I2(fdat[8]),
        .I3(fdat[10]),
        .I4(\nir_id[21]_i_4_n_0 ),
        .I5(fdat[15]),
        .O(\fch/lir_id_0 [21]));
  LUT6 #(
    .INIT(64'hAAAAFAABAAAAAAAA)) 
    \nir_id[21]_i_2 
       (.I0(\nir_id[21]_i_5_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(\nir_id[21]_i_6_n_0 ),
        .I5(\nir_id[21]_i_7_n_0 ),
        .O(\nir_id[21]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[21]_i_3 
       (.I0(fdat[0]),
        .I1(fdat[1]),
        .O(\nir_id[21]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[21]_i_4 
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .O(\nir_id[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF600000000000000)) 
    \nir_id[21]_i_5 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(\nir_id[21]_i_8_n_0 ),
        .I3(\nir_id[15]_i_2_n_0 ),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(\nir_id[21]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h55FFFFFE)) 
    \nir_id[21]_i_6 
       (.I0(fdat[11]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .O(\nir_id[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC000C00100000000)) 
    \nir_id[21]_i_7 
       (.I0(fdat[2]),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .I5(\nir_id[14]_i_6_n_0 ),
        .O(\nir_id[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h8988000000000000)) 
    \nir_id[21]_i_8 
       (.I0(fdat[5]),
        .I1(fdat[6]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[7]),
        .I5(fdat[10]),
        .O(\nir_id[21]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h0000EBFB)) 
    \nir_id[24]_i_1 
       (.I0(\fch/stat [2]),
        .I1(\fch/fch_issu1_ir ),
        .I2(\fch/stat [1]),
        .I3(fch_term),
        .I4(\nir_id[24]_i_3_n_0 ),
        .O(\fch/fctl/fch_nir_lir ));
  LUT6 #(
    .INIT(64'h0000000301020202)) 
    \nir_id[24]_i_10 
       (.I0(fdat[1]),
        .I1(\nir_id[24]_i_14_n_0 ),
        .I2(fdat[13]),
        .I3(fdat[3]),
        .I4(fdat[2]),
        .I5(fdat[0]),
        .O(\nir_id[24]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_11 
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .O(\nir_id[24]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_12 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[24]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[24]_i_13 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .O(\nir_id[24]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \nir_id[24]_i_14 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[7]),
        .I3(fdat[12]),
        .O(\nir_id[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFBBFB)) 
    \nir_id[24]_i_2 
       (.I0(\nir_id[24]_i_4_n_0 ),
        .I1(\nir_id[24]_i_5_n_0 ),
        .I2(\nir_id[24]_i_6_n_0 ),
        .I3(\nir_id[24]_i_7_n_0 ),
        .I4(\nir_id[24]_i_8_n_0 ),
        .I5(fdat[15]),
        .O(\fch/lir_id_0 [24]));
  LUT6 #(
    .INIT(64'hBFFBBFFBFFFFFFF3)) 
    \nir_id[24]_i_3 
       (.I0(\fadr[15]_INST_0_i_8_n_0 ),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(\fch/stat [0]),
        .I3(\nir_id[24]_i_9_n_0 ),
        .I4(\fadr[15]_INST_0_i_4_n_0 ),
        .I5(fch_term),
        .O(\nir_id[24]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0440)) 
    \nir_id[24]_i_4 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(\nir_id[24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3F7FFF7FFF7FFF7F)) 
    \nir_id[24]_i_5 
       (.I0(\nir_id[24]_i_10_n_0 ),
        .I1(\nir_id[24]_i_11_n_0 ),
        .I2(\nir_id[24]_i_12_n_0 ),
        .I3(fdat[9]),
        .I4(fdat[7]),
        .I5(fdat[12]),
        .O(\nir_id[24]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF11F1F1F111F1F1F)) 
    \nir_id[24]_i_6 
       (.I0(fdat[9]),
        .I1(fdat[10]),
        .I2(fdat[6]),
        .I3(fdat[4]),
        .I4(fdat[5]),
        .I5(fdat[3]),
        .O(\nir_id[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5FFFFFFFFFFFEFFF)) 
    \nir_id[24]_i_7 
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(\nir_id[24]_i_13_n_0 ),
        .I4(fdat[10]),
        .I5(fdat[9]),
        .O(\nir_id[24]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h7776)) 
    \nir_id[24]_i_8 
       (.I0(fdat[13]),
        .I1(fdat[14]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(\nir_id[24]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[24]_i_9 
       (.I0(\fch/stat [1]),
        .I1(\fch/stat [2]),
        .O(\nir_id[24]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    \pc0[0]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\pc0[15]_i_3_n_0 ),
        .I2(\fch/p_2_in [0]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\rgf/pcnt/pc [0]),
        .O(fch_pc[0]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[10]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [10]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [10]),
        .O(fch_pc[10]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[11]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [11]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [11]),
        .O(fch_pc[11]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[12]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_4 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [12]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [12]),
        .O(fch_pc[12]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[13]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__2_n_7 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [13]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [13]),
        .O(fch_pc[13]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[14]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__2_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [14]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [14]),
        .O(fch_pc[14]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[15]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__2_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [15]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [15]),
        .O(fch_pc[15]));
  LUT6 #(
    .INIT(64'h11515151FFFFFFFF)) 
    \pc0[15]_i_2 
       (.I0(\fadr[15]_INST_0_i_7_n_0 ),
        .I1(\fadr[15]_INST_0_i_6_n_0 ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(\fch/stat [2]),
        .I5(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\pc0[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBB2BFFFF)) 
    \pc0[15]_i_3 
       (.I0(irq_lev[1]),
        .I1(\rgf/sreg/sr [3]),
        .I2(\rgf/sreg/sr [2]),
        .I3(irq_lev[0]),
        .I4(irq),
        .O(\pc0[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \pc0[15]_i_4 
       (.I0(\fch/fch_issu1 ),
        .I1(\fadr[15]_INST_0_i_8_n_0 ),
        .O(\pc0[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hE2F0E2F0E2FFE200)) 
    \pc0[1]_i_1 
       (.I0(\fch/fch_pc_nx4_carry_n_7 ),
        .I1(\pc0[15]_i_2_n_0 ),
        .I2(\fch/p_2_in [1]),
        .I3(\pc0[15]_i_3_n_0 ),
        .I4(\rgf/pcnt/pc [1]),
        .I5(\pc0[15]_i_4_n_0 ),
        .O(fch_pc[1]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[2]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [2]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [2]),
        .O(fch_pc[2]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[3]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [3]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [3]),
        .O(fch_pc[3]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[4]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry_n_4 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [4]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [4]),
        .O(fch_pc[4]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[5]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_7 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [5]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [5]),
        .O(fch_pc[5]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[6]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [6]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [6]),
        .O(fch_pc[6]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[7]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [7]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [7]),
        .O(fch_pc[7]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[8]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_4 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [8]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [8]),
        .O(fch_pc[8]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    \pc0[9]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_7 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [9]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [9]),
        .O(fch_pc[9]));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_1
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [7]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [7]),
        .O(pc10_carry__0_i_1_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_2
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [6]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [6]),
        .O(pc10_carry__0_i_2_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_3
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_7 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [5]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [5]),
        .O(pc10_carry__0_i_3_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__0_i_4
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry_n_4 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [4]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [4]),
        .O(pc10_carry__0_i_4_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_1
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [11]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [11]),
        .O(pc10_carry__1_i_1_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_2
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [10]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [10]),
        .O(pc10_carry__1_i_2_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_3
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_7 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [9]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [9]),
        .O(pc10_carry__1_i_3_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__1_i_4
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__0_n_4 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [8]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [8]),
        .O(pc10_carry__1_i_4_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_1
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__2_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [15]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [15]),
        .O(pc10_carry__2_i_1_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_2
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__2_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [14]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [14]),
        .O(pc10_carry__2_i_2_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_3
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__2_n_7 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [13]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [13]),
        .O(pc10_carry__2_i_3_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry__2_i_4
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry__1_n_4 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [12]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [12]),
        .O(pc10_carry__2_i_4_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry_i_1
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry_n_5 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [3]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [3]),
        .O(pc10_carry_i_1_n_0));
  LUT6 #(
    .INIT(64'hEF40EF4FEF40E040)) 
    pc10_carry_i_2
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\fch/fch_pc_nx4_carry_n_6 ),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [2]),
        .I4(\pc0[15]_i_4_n_0 ),
        .I5(\rgf/pcnt/pc [2]),
        .O(pc10_carry_i_2_n_0));
  LUT6 #(
    .INIT(64'h01FB010B01FBF1FB)) 
    pc10_carry_i_3
       (.I0(\pc0[15]_i_4_n_0 ),
        .I1(\rgf/pcnt/pc [1]),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\fch/p_2_in [1]),
        .I4(\pc0[15]_i_2_n_0 ),
        .I5(\fch/fch_pc_nx4_carry_n_7 ),
        .O(pc10_carry_i_3_n_0));
  LUT5 #(
    .INIT(32'hF4F7B080)) 
    pc10_carry_i_4
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\pc0[15]_i_3_n_0 ),
        .I2(\fch/p_2_in [0]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\rgf/pcnt/pc [0]),
        .O(pc10_carry_i_4_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[0]_i_2_n_0 ),
        .O(\rgf/pcnt/p_1_in [0]));
  LUT6 #(
    .INIT(64'hF4F7FFFFB0800000)) 
    \pc[0]_i_2 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(\pc0[15]_i_3_n_0 ),
        .I2(\fch/p_2_in [0]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc[15]_i_8_n_0 ),
        .I5(\rgf/pcnt/pc [0]),
        .O(\pc[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[10]_i_2_n_0 ),
        .O(\rgf/pcnt/p_1_in [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[10]_i_2 
       (.I0(fch_pc[10]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [10]),
        .O(\pc[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[11]_i_2_n_0 ),
        .O(\rgf/pcnt/p_1_in [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[11]_i_2 
       (.I0(fch_pc[11]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [11]),
        .O(\pc[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[12]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[12]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [12]),
        .O(\rgf/rgf_c1bus_0 [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[12]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [12]),
        .O(\rgf/rgf_c0bus_0 [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[12]_i_4 
       (.I0(fch_pc[12]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [12]),
        .O(\pc[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[13]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[13]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [13]),
        .O(\rgf/rgf_c1bus_0 [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[13]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [13]),
        .O(\rgf/rgf_c0bus_0 [13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[13]_i_4 
       (.I0(fch_pc[13]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [13]),
        .O(\pc[13]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[14]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[14]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [14]),
        .O(\rgf/rgf_c1bus_0 [14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[14]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [14]),
        .O(\rgf/rgf_c0bus_0 [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[14]_i_4 
       (.I0(fch_pc[14]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [14]),
        .O(\pc[14]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[15]_i_6_n_0 ),
        .O(\rgf/pcnt/p_1_in [15]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[15]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [15]),
        .O(\rgf/rgf_c1bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_4 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[15]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [15]),
        .O(\rgf/rgf_c0bus_0 [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_5 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[15]_i_6 
       (.I0(fch_pc[15]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [15]),
        .O(\pc[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hE4E0A0E0FFFFFFFF)) 
    \pc[15]_i_7 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\rgf_selc0_wb[0]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_wb [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\pc[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \pc[15]_i_8 
       (.I0(fch_term),
        .I1(\fadr[15]_INST_0_i_4_n_0 ),
        .O(\pc[15]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[1]_i_2_n_0 ),
        .O(\rgf/pcnt/p_1_in [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[1]_i_2 
       (.I0(fch_pc[1]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [1]),
        .O(\pc[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[2]_i_2_n_0 ),
        .O(\rgf/pcnt/p_1_in [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[2]_i_2 
       (.I0(fch_pc[2]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [2]),
        .O(\pc[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[3]_i_2_n_0 ),
        .O(\rgf/pcnt/p_1_in [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[3]_i_2 
       (.I0(fch_pc[3]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [3]),
        .O(\pc[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[4]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[4]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [4]),
        .O(\rgf/rgf_c1bus_0 [4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[4]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [4]),
        .O(\rgf/rgf_c0bus_0 [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[4]_i_4 
       (.I0(fch_pc[4]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [4]),
        .O(\pc[4]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[5]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [5]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[5]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[5]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [5]),
        .O(\rgf/rgf_c1bus_0 [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[5]_i_3 
       (.I0(fch_pc[5]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [5]),
        .O(\pc[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[6]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[6]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[6]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [6]),
        .O(\rgf/rgf_c0bus_0 [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[6]_i_3 
       (.I0(fch_pc[6]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [6]),
        .O(\pc[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[7]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[7]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[7]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [7]),
        .O(\rgf/rgf_c0bus_0 [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[7]_i_3 
       (.I0(fch_pc[7]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [7]),
        .O(\pc[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[8]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[8]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [8]),
        .O(\rgf/rgf_c1bus_0 [8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[8]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [8]),
        .O(\rgf/rgf_c0bus_0 [8]));
  LUT6 #(
    .INIT(64'hB8BBFFFFB8880000)) 
    \pc[8]_i_4 
       (.I0(\pc[8]_i_5_n_0 ),
        .I1(\pc0[15]_i_3_n_0 ),
        .I2(\fch/p_2_in [8]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc[15]_i_8_n_0 ),
        .I5(\rgf/pcnt/pc [8]),
        .O(\pc[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEAAAA0222AAAA)) 
    \pc[8]_i_5 
       (.I0(\fch/p_2_in [8]),
        .I1(\fadr[15]_INST_0_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_6_n_0 ),
        .I3(\pc[8]_i_6_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fch/fch_pc_nx4_carry__0_n_4 ),
        .O(\pc[8]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \pc[8]_i_6 
       (.I0(\fch/stat [2]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .O(\pc[8]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [1]),
        .I4(\pc[9]_i_2_n_0 ),
        .O(\rgf/pcnt/p_1_in [9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc[9]_i_2 
       (.I0(fch_pc[9]),
        .I1(\pc[15]_i_8_n_0 ),
        .I2(\rgf/pcnt/pc [9]),
        .O(\pc[9]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \read_cyc[3]_i_1 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(\mem/mem_accslot ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[0]_INST_0_i_1 
       (.I0(\badr[0]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [0]),
        .I2(\rgf/bank02/p_0_in [0]),
        .I3(\badr[0]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [0]),
        .I5(\rgf/a0bus_out/badr[0]_INST_0_i_8_n_0 ),
        .O(a0bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[0]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [0]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [0]),
        .I4(fch_pc0[0]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[10]_INST_0_i_1 
       (.I0(\badr[10]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [10]),
        .I2(\rgf/bank02/p_0_in [10]),
        .I3(\badr[10]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [10]),
        .I5(\rgf/a0bus_out/badr[10]_INST_0_i_8_n_0 ),
        .O(a0bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[10]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc0[10]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[11]_INST_0_i_1 
       (.I0(\badr[11]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [11]),
        .I2(\rgf/bank02/p_0_in [11]),
        .I3(\badr[11]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [11]),
        .I5(\rgf/a0bus_out/badr[11]_INST_0_i_8_n_0 ),
        .O(a0bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[11]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc0[11]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[11]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[12]_INST_0_i_1 
       (.I0(\badr[12]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [12]),
        .I2(\rgf/bank02/p_0_in [12]),
        .I3(\badr[12]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [12]),
        .I5(\rgf/a0bus_out/badr[12]_INST_0_i_8_n_0 ),
        .O(a0bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[12]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc0[12]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[13]_INST_0_i_1 
       (.I0(\badr[13]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [13]),
        .I2(\rgf/bank02/p_0_in [13]),
        .I3(\badr[13]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [13]),
        .I5(\rgf/a0bus_out/badr[13]_INST_0_i_8_n_0 ),
        .O(a0bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[13]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc0[13]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[14]_INST_0_i_1 
       (.I0(\badr[14]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [14]),
        .I2(\rgf/bank02/p_0_in [14]),
        .I3(\badr[14]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [14]),
        .I5(\rgf/a0bus_out/badr[14]_INST_0_i_8_n_0 ),
        .O(a0bus_0[14]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[14]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc0[14]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[14]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[15]_INST_0_i_1 
       (.I0(\badr[15]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [15]),
        .I2(\rgf/bank02/p_0_in [15]),
        .I3(\badr[15]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [15]),
        .I5(\rgf/a0bus_out/badr[15]_INST_0_i_8_n_0 ),
        .O(a0bus_0[15]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[15]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc0[15]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[15]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[1]_INST_0_i_1 
       (.I0(\badr[1]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [1]),
        .I2(\rgf/bank02/p_0_in [1]),
        .I3(\badr[1]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [1]),
        .I5(\rgf/a0bus_out/badr[1]_INST_0_i_8_n_0 ),
        .O(a0bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[1]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc0[1]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[2]_INST_0_i_1 
       (.I0(\badr[2]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [2]),
        .I2(\rgf/bank02/p_0_in [2]),
        .I3(\badr[2]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [2]),
        .I5(\rgf/a0bus_out/badr[2]_INST_0_i_8_n_0 ),
        .O(a0bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[2]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc0[2]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[3]_INST_0_i_1 
       (.I0(\badr[3]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [3]),
        .I2(\rgf/bank02/p_0_in [3]),
        .I3(\badr[3]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [3]),
        .I5(\rgf/a0bus_out/badr[3]_INST_0_i_8_n_0 ),
        .O(a0bus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[3]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc0[3]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[4]_INST_0_i_1 
       (.I0(\badr[4]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [4]),
        .I2(\rgf/bank02/p_0_in [4]),
        .I3(\badr[4]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [4]),
        .I5(\rgf/a0bus_out/badr[4]_INST_0_i_8_n_0 ),
        .O(a0bus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[4]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc0[4]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[4]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[5]_INST_0_i_1 
       (.I0(\badr[5]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [5]),
        .I2(\rgf/bank02/p_0_in [5]),
        .I3(\badr[5]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [5]),
        .I5(\rgf/a0bus_out/badr[5]_INST_0_i_8_n_0 ),
        .O(a0bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[5]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc0[5]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[5]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[6]_INST_0_i_1 
       (.I0(\badr[6]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [6]),
        .I2(\rgf/bank02/p_0_in [6]),
        .I3(\badr[6]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [6]),
        .I5(\rgf/a0bus_out/badr[6]_INST_0_i_8_n_0 ),
        .O(a0bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[6]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc0[6]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[7]_INST_0_i_1 
       (.I0(\badr[7]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [7]),
        .I2(\rgf/bank02/p_0_in [7]),
        .I3(\badr[7]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [7]),
        .I5(\rgf/a0bus_out/badr[7]_INST_0_i_8_n_0 ),
        .O(a0bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[7]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc0[7]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[8]_INST_0_i_1 
       (.I0(\badr[8]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [8]),
        .I2(\rgf/bank02/p_0_in [8]),
        .I3(\badr[8]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [8]),
        .I5(\rgf/a0bus_out/badr[8]_INST_0_i_8_n_0 ),
        .O(a0bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[8]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc0[8]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[9]_INST_0_i_1 
       (.I0(\badr[9]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in [9]),
        .I2(\rgf/bank02/p_0_in [9]),
        .I3(\badr[9]_INST_0_i_6_n_0 ),
        .I4(\rgf/a0bus_b13 [9]),
        .I5(\rgf/a0bus_out/badr[9]_INST_0_i_8_n_0 ),
        .O(a0bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[9]_INST_0_i_8 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc0[9]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[9]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/rgf_c0bus_wb[12]_i_35 
       (.I0(\rgf/a0bus_out/badr[15]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_37_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_38_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_33_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_34_n_0 ),
        .I5(\badr[15]_INST_0_i_6_n_0 ),
        .O(\rgf/a0bus_out/rgf_c0bus_wb[12]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[0]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [0]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [0]),
        .I4(fch_pc1[0]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[0]_INST_0_i_2 
       (.I0(\badr[0]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [0]),
        .I2(\rgf/bank02/p_0_in0_in [0]),
        .I3(\badr[0]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [0]),
        .I5(\rgf/a1bus_out/badr[0]_INST_0_i_14_n_0 ),
        .O(a1bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[10]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc1[10]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[10]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[10]_INST_0_i_2 
       (.I0(\badr[10]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [10]),
        .I2(\rgf/bank02/p_0_in0_in [10]),
        .I3(\badr[10]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [10]),
        .I5(\rgf/a1bus_out/badr[10]_INST_0_i_14_n_0 ),
        .O(a1bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[11]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc1[11]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[11]_INST_0_i_2 
       (.I0(\badr[11]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [11]),
        .I2(\rgf/bank02/p_0_in0_in [11]),
        .I3(\badr[11]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [11]),
        .I5(\rgf/a1bus_out/badr[11]_INST_0_i_14_n_0 ),
        .O(a1bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[12]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc1[12]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[12]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[12]_INST_0_i_2 
       (.I0(\badr[12]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [12]),
        .I2(\rgf/bank02/p_0_in0_in [12]),
        .I3(\badr[12]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [12]),
        .I5(\rgf/a1bus_out/badr[12]_INST_0_i_14_n_0 ),
        .O(a1bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[13]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc1[13]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[13]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[13]_INST_0_i_2 
       (.I0(\badr[13]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [13]),
        .I2(\rgf/bank02/p_0_in0_in [13]),
        .I3(\badr[13]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [13]),
        .I5(\rgf/a1bus_out/badr[13]_INST_0_i_14_n_0 ),
        .O(a1bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[14]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc1[14]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[14]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[14]_INST_0_i_2 
       (.I0(\badr[14]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [14]),
        .I2(\rgf/bank02/p_0_in0_in [14]),
        .I3(\badr[14]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [14]),
        .I5(\rgf/a1bus_out/badr[14]_INST_0_i_14_n_0 ),
        .O(a1bus_0[14]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[15]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc1[15]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[15]_INST_0_i_2 
       (.I0(\badr[15]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [15]),
        .I2(\rgf/bank02/p_0_in0_in [15]),
        .I3(\badr[15]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [15]),
        .I5(\rgf/a1bus_out/badr[15]_INST_0_i_14_n_0 ),
        .O(a1bus_0[15]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[1]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc1[1]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[1]_INST_0_i_2 
       (.I0(\badr[1]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [1]),
        .I2(\rgf/bank02/p_0_in0_in [1]),
        .I3(\badr[1]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [1]),
        .I5(\rgf/a1bus_out/badr[1]_INST_0_i_14_n_0 ),
        .O(a1bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[2]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc1[2]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[2]_INST_0_i_2 
       (.I0(\badr[2]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [2]),
        .I2(\rgf/bank02/p_0_in0_in [2]),
        .I3(\badr[2]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [2]),
        .I5(\rgf/a1bus_out/badr[2]_INST_0_i_14_n_0 ),
        .O(a1bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[3]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc1[3]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[3]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[3]_INST_0_i_2 
       (.I0(\badr[3]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [3]),
        .I2(\rgf/bank02/p_0_in0_in [3]),
        .I3(\badr[3]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [3]),
        .I5(\rgf/a1bus_out/badr[3]_INST_0_i_14_n_0 ),
        .O(a1bus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[4]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc1[4]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[4]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[4]_INST_0_i_2 
       (.I0(\badr[4]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [4]),
        .I2(\rgf/bank02/p_0_in0_in [4]),
        .I3(\badr[4]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [4]),
        .I5(\rgf/a1bus_out/badr[4]_INST_0_i_14_n_0 ),
        .O(a1bus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[5]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc1[5]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[5]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[5]_INST_0_i_2 
       (.I0(\badr[5]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [5]),
        .I2(\rgf/bank02/p_0_in0_in [5]),
        .I3(\badr[5]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [5]),
        .I5(\rgf/a1bus_out/badr[5]_INST_0_i_14_n_0 ),
        .O(a1bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[6]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc1[6]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[6]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[6]_INST_0_i_2 
       (.I0(\badr[6]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [6]),
        .I2(\rgf/bank02/p_0_in0_in [6]),
        .I3(\badr[6]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [6]),
        .I5(\rgf/a1bus_out/badr[6]_INST_0_i_14_n_0 ),
        .O(a1bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[7]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc1[7]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[7]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[7]_INST_0_i_2 
       (.I0(\badr[7]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [7]),
        .I2(\rgf/bank02/p_0_in0_in [7]),
        .I3(\badr[7]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [7]),
        .I5(\rgf/a1bus_out/badr[7]_INST_0_i_14_n_0 ),
        .O(a1bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[8]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc1[8]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[8]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[8]_INST_0_i_2 
       (.I0(\badr[8]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [8]),
        .I2(\rgf/bank02/p_0_in0_in [8]),
        .I3(\badr[8]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [8]),
        .I5(\rgf/a1bus_out/badr[8]_INST_0_i_14_n_0 ),
        .O(a1bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[9]_INST_0_i_14 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc1[9]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[9]_INST_0_i_2 
       (.I0(\badr[9]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [9]),
        .I2(\rgf/bank02/p_0_in0_in [9]),
        .I3(\badr[9]_INST_0_i_12_n_0 ),
        .I4(\rgf/a1bus_b13 [9]),
        .I5(\rgf/a1bus_out/badr[9]_INST_0_i_14_n_0 ),
        .O(a1bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[10]_i_25 
       (.I0(\rgf/a1bus_out/badr[15]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_26_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_27_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_58_n_0 ),
        .I5(\badr[15]_INST_0_i_12_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[10]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[0]_INST_0_i_4 
       (.I0(\rgf/treg/tr [0]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [0]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[0]_INST_0_i_6 
       (.I0(\bbus_o[0]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_20_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[0]_INST_0_i_7 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [0]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [0]),
        .I4(fch_pc0[0]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[0]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[1]_INST_0_i_3 
       (.I0(\rgf/treg/tr [1]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [1]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[1]_INST_0_i_5 
       (.I0(\bbus_o[1]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_15_n_0 ),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_17_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_18_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_19_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[1]_INST_0_i_6 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc0[1]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[1]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[2]_INST_0_i_4 
       (.I0(\rgf/treg/tr [2]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [2]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[2]_INST_0_i_6 
       (.I0(\bbus_o[2]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_18_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_19_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_20_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[2]_INST_0_i_7 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc0[2]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[2]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[3]_INST_0_i_4 
       (.I0(\rgf/treg/tr [3]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [3]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[3]_INST_0_i_6 
       (.I0(\bbus_o[3]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_18_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_19_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_20_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[3]_INST_0_i_7 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc0[3]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[3]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[4]_INST_0_i_4 
       (.I0(\rgf/treg/tr [4]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [4]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[4]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[4]_INST_0_i_6 
       (.I0(\bbus_o[4]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_18_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_19_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_20_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[4]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[4]_INST_0_i_7 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc0[4]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[4]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[5]_INST_0_i_13 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc0[5]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[5]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[5]_INST_0_i_4 
       (.I0(\rgf/treg/tr [5]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [5]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[5]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[5]_INST_0_i_7 
       (.I0(\rgf/b0bus_out/bbus_o[5]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_17_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_18_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[5]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[6]_INST_0_i_13 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc0[6]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[6]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[6]_INST_0_i_4 
       (.I0(\rgf/treg/tr [6]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [6]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[6]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[6]_INST_0_i_7 
       (.I0(\rgf/b0bus_out/bbus_o[6]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17_n_0 ),
        .I5(\bbus_o[6]_INST_0_i_18_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[6]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[7]_INST_0_i_13 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc0[7]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[7]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[7]_INST_0_i_4 
       (.I0(\rgf/treg/tr [7]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [7]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[7]_INST_0_i_7 
       (.I0(\rgf/b0bus_out/bbus_o[7]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17_n_0 ),
        .I5(\bbus_o[7]_INST_0_i_18_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[7]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[10]_INST_0_i_18 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc0[10]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[10]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[10]_INST_0_i_6 
       (.I0(\rgf/bank02/p_0_in2_in [10]),
        .I1(\rgf/bank02/p_1_in3_in [10]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [10]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [10]),
        .O(\rgf/b0bus_out/bdatw[10]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[10]_INST_0_i_7 
       (.I0(\rgf/b0bus_out/bdatw[10]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [10]),
        .I2(\rgf/bank13/p_0_in2_in [10]),
        .I3(\rgf/b0bus_sel_cr [0]),
        .I4(\rgf/sreg/sr [10]),
        .O(\rgf/b0bus_out/bdatw[10]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[11]_INST_0_i_21 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc0[11]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[11]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bdatw[11]_INST_0_i_6 
       (.I0(\rgf/treg/tr [11]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [11]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bdatw[11]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bdatw[11]_INST_0_i_9 
       (.I0(\rgf/b0bus_out/bdatw[11]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_22_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_23_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_24_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_25_n_0 ),
        .I5(\bdatw[11]_INST_0_i_26_n_0 ),
        .O(\rgf/b0bus_out/bdatw[11]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[12]_INST_0_i_22 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc0[12]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[12]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bdatw[12]_INST_0_i_6 
       (.I0(\rgf/treg/tr [12]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [12]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bdatw[12]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bdatw[12]_INST_0_i_9 
       (.I0(\rgf/b0bus_out/bdatw[12]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_23_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_24_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_25_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_26_n_0 ),
        .I5(\bdatw[12]_INST_0_i_27_n_0 ),
        .O(\rgf/b0bus_out/bdatw[12]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[13]_INST_0_i_22 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc0[13]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[13]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bdatw[13]_INST_0_i_6 
       (.I0(\rgf/treg/tr [13]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [13]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bdatw[13]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bdatw[13]_INST_0_i_9 
       (.I0(\rgf/b0bus_out/bdatw[13]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_23_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_24_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_25_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_26_n_0 ),
        .I5(\bdatw[13]_INST_0_i_27_n_0 ),
        .O(\rgf/b0bus_out/bdatw[13]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[14]_INST_0_i_23 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc0[14]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[14]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bdatw[14]_INST_0_i_6 
       (.I0(\rgf/treg/tr [14]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [14]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bdatw[14]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bdatw[14]_INST_0_i_9 
       (.I0(\rgf/b0bus_out/bdatw[14]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_27_n_0 ),
        .I5(\bdatw[14]_INST_0_i_28_n_0 ),
        .O(\rgf/b0bus_out/bdatw[14]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bdatw[15]_INST_0_i_11 
       (.I0(\rgf/b0bus_out/bdatw[15]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_37_n_0 ),
        .I5(\bdatw[15]_INST_0_i_38_n_0 ),
        .O(\rgf/b0bus_out/bdatw[15]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[15]_INST_0_i_33 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc0[15]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[15]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bdatw[15]_INST_0_i_8 
       (.I0(\rgf/treg/tr [15]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [15]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bdatw[15]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[8]_INST_0_i_22 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc0[8]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[8]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[8]_INST_0_i_6 
       (.I0(\rgf/bank02/p_0_in2_in [8]),
        .I1(\rgf/bank02/p_1_in3_in [8]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [8]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [8]),
        .O(\rgf/b0bus_out/bdatw[8]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[8]_INST_0_i_7 
       (.I0(\rgf/b0bus_out/bdatw[8]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [8]),
        .I2(\rgf/bank13/p_0_in2_in [8]),
        .I3(\rgf/b0bus_sel_cr [0]),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf/b0bus_out/bdatw[8]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[9]_INST_0_i_17 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc0[9]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[9]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[9]_INST_0_i_5 
       (.I0(\rgf/bank02/p_0_in2_in [9]),
        .I1(\rgf/bank02/p_1_in3_in [9]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [9]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [9]),
        .O(\rgf/b0bus_out/bdatw[9]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[9]_INST_0_i_6 
       (.I0(\rgf/b0bus_out/bdatw[9]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [9]),
        .I2(\rgf/bank13/p_0_in2_in [9]),
        .I3(\rgf/b0bus_sel_cr [0]),
        .I4(\rgf/sreg/sr [9]),
        .O(\rgf/b0bus_out/bdatw[9]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_10 
       (.I0(\rgf/treg/tr [10]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [10]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_13 
       (.I0(\rgf/b1bus_out/bdatw[10]_INST_0_i_27_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_28_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_29_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_30_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_31_n_0 ),
        .I5(\bdatw[10]_INST_0_i_32_n_0 ),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_27 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc1[10]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_35 
       (.I0(\rgf/treg/tr [2]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [2]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_38 
       (.I0(\rgf/b1bus_out/bdatw[10]_INST_0_i_62_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_63_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_64_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_65_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_66_n_0 ),
        .I5(\bdatw[10]_INST_0_i_67_n_0 ),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_62 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc1[2]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_12 
       (.I0(\rgf/treg/tr [11]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [11]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_15 
       (.I0(\rgf/b1bus_out/bdatw[11]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_37_n_0 ),
        .I5(\bdatw[11]_INST_0_i_38_n_0 ),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_33 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc1[11]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_41 
       (.I0(\rgf/treg/tr [3]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [3]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_44 
       (.I0(\rgf/b1bus_out/bdatw[11]_INST_0_i_66_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_67_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_68_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_69_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_70_n_0 ),
        .I5(\bdatw[11]_INST_0_i_71_n_0 ),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_66 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc1[3]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_12 
       (.I0(\rgf/treg/tr [12]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [12]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_15 
       (.I0(\rgf/b1bus_out/bdatw[12]_INST_0_i_32_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_33_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_34_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_35_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_36_n_0 ),
        .I5(\bdatw[12]_INST_0_i_37_n_0 ),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_32 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc1[12]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_40 
       (.I0(\rgf/treg/tr [4]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [4]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_43 
       (.I0(\rgf/b1bus_out/bdatw[12]_INST_0_i_65_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_66_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_67_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_68_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_69_n_0 ),
        .I5(\bdatw[12]_INST_0_i_70_n_0 ),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_65 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc1[4]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_65_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_12 
       (.I0(\rgf/treg/tr [13]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [13]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_15 
       (.I0(\rgf/b1bus_out/bdatw[13]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_37_n_0 ),
        .I5(\bdatw[13]_INST_0_i_38_n_0 ),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_33 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc1[13]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_41 
       (.I0(\rgf/treg/tr [5]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [5]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_44 
       (.I0(\rgf/b1bus_out/bdatw[13]_INST_0_i_62_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_63_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_64_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_65_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_66_n_0 ),
        .I5(\bdatw[13]_INST_0_i_67_n_0 ),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_62 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc1[5]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_12 
       (.I0(\rgf/treg/tr [14]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [14]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_15 
       (.I0(\rgf/b1bus_out/bdatw[14]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_36_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_39_n_0 ),
        .I5(\bdatw[14]_INST_0_i_40_n_0 ),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_35 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc1[14]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_43 
       (.I0(\rgf/treg/tr [6]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [6]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_46 
       (.I0(\rgf/b1bus_out/bdatw[14]_INST_0_i_64_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_65_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_66_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_67_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_68_n_0 ),
        .I5(\bdatw[14]_INST_0_i_69_n_0 ),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_64 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc1[6]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_14 
       (.I0(\rgf/treg/tr [15]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [15]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_147 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc1[7]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_17 
       (.I0(\rgf/b1bus_out/bdatw[15]_INST_0_i_54_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_55_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_56_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_58_n_0 ),
        .I5(\bdatw[15]_INST_0_i_59_n_0 ),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_54 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc1[15]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_62 
       (.I0(\rgf/treg/tr [7]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [7]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_65 
       (.I0(\rgf/b1bus_out/bdatw[15]_INST_0_i_147_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_148_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_149_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_150_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_151_n_0 ),
        .I5(\bdatw[15]_INST_0_i_152_n_0 ),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_65_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_10 
       (.I0(\rgf/treg/tr [8]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [8]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_13 
       (.I0(\rgf/b1bus_out/bdatw[8]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_32_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_33_n_0 ),
        .I5(\bdatw[8]_INST_0_i_34_n_0 ),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_29 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc1[8]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_37 
       (.I0(\rgf/treg/tr [0]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [0]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_40 
       (.I0(\rgf/b1bus_out/bdatw[8]_INST_0_i_68_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_69_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_70_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_71_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_72_n_0 ),
        .I5(\bdatw[8]_INST_0_i_73_n_0 ),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_68 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [0]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [0]),
        .I4(fch_pc1[0]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_12 
       (.I0(\rgf/b1bus_out/bdatw[9]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_28_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29_n_0 ),
        .I5(\bdatw[9]_INST_0_i_30_n_0 ),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_25 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc1[9]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_32 
       (.I0(\rgf/treg/tr [1]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [1]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_35 
       (.I0(\rgf/b1bus_out/bdatw[9]_INST_0_i_59_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_60_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_61_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_62_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_63_n_0 ),
        .I5(\bdatw[9]_INST_0_i_64_n_0 ),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_59 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc1[1]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_9 
       (.I0(\rgf/treg/tr [9]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [9]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [0]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [0]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [10]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [10]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [10]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [10]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [11]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [11]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [11]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [11]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [12]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [12]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [12]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [12]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [13]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [13]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [13]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [13]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [14]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [14]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [14]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [14]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_19 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_20 
       (.I0(\rgf/bank02/gr00 [15]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [15]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_21 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_22 
       (.I0(\rgf/bank02/gr04 [15]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [15]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_1_in [15]));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_71 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(ctl_sela0_rn[0]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_72 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[0]),
        .I4(\badr[15]_INST_0_i_28_n_0 ),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_73 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_74 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\badr[15]_INST_0_i_191_n_0 ),
        .I5(ctl_sela0_rn[2]),
        .O(\bank02/a0buso/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_75 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_76 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_77 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_78 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [1]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [1]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [2]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [2]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [3]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [3]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [3]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [3]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [4]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [4]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [5]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [5]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [5]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [5]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [6]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [6]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [6]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [6]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [7]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [7]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [7]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [7]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [8]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [8]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [8]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [8]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [9]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [9]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [9]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [9]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_4 
       (.I0(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_17_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [0]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [0]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [10]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [10]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [10]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [10]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [11]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [11]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [11]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [11]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [12]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [12]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [12]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [12]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [13]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [13]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [13]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [13]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [14]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [14]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [14]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [14]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_23 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_24 
       (.I0(\rgf/bank02/gr20 [15]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [15]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_25 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_26 
       (.I0(\rgf/bank02/gr24 [15]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [15]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/p_0_in [15]));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_79 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_sela0_rn[2]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(ctl_sela0_rn[0]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_80 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[0]),
        .I4(\badr[15]_INST_0_i_28_n_0 ),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso2l/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_81 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_82 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\badr[15]_INST_0_i_191_n_0 ),
        .I5(ctl_sela0_rn[2]),
        .O(\bank02/a0buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_83 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso2l/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_84 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso2l/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_85 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_86 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank02/a0buso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [1]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [1]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [2]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [2]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [3]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [3]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [3]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [3]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [4]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [4]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [5]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [5]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [5]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [5]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [6]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [6]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [6]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [6]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [7]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [7]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [7]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [7]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [8]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [8]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [8]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [8]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [9]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [9]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [9]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [9]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_5 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in [9]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_33 
       (.I0(\rgf/bank02/gr04 [0]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [0]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [10]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [10]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [10]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [10]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [11]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [11]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_33 
       (.I0(\rgf/bank02/gr04 [11]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [11]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [12]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [12]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [12]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [12]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [13]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [13]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [13]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [13]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [14]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [14]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [14]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [14]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_43_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_44_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_45_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [15]));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_124 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(ctl_sela1_rn),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_125 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_52_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_126 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_127 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_235_n_0 ),
        .I5(\badr[15]_INST_0_i_40_n_0 ),
        .O(\bank02/a1buso/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_128 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_129 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_130 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(ctl_sela1_rn),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_131 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_43 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_44 
       (.I0(\rgf/bank02/gr00 [15]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [15]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_45 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_46 
       (.I0(\rgf/bank02/gr04 [15]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [15]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [1]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [1]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [2]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [2]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [3]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [3]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_33 
       (.I0(\rgf/bank02/gr04 [3]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [3]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [4]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [4]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [5]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [5]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [5]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [5]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [6]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [6]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [6]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [6]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [7]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [7]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_33 
       (.I0(\rgf/bank02/gr04 [7]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [7]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [8]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [8]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [8]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [8]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_10 
       (.I0(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [9]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [9]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/a1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/a1buso/gr1_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [9]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [9]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_34 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [0]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [0]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [10]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [10]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [10]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [10]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_34 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [11]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [11]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [11]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [11]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [12]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [12]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [12]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [12]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [13]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [13]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [13]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [13]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [14]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [14]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [14]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [14]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_47_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_48_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_49_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_50_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [15]));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_132 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(ctl_sela1_rn),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_133 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_52_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso2l/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_134 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_135 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_235_n_0 ),
        .I5(\badr[15]_INST_0_i_40_n_0 ),
        .O(\bank02/a1buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_136 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso2l/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_137 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso2l/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_138 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(ctl_sela1_rn),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_139 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank02/a1buso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_47 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_48 
       (.I0(\rgf/bank02/gr20 [15]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [15]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_49 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_50 
       (.I0(\rgf/bank02/gr24 [15]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [15]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [1]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [1]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [2]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [2]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_34 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [3]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [3]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [3]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [3]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [4]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [4]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [5]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [5]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [5]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [5]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [6]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [6]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [6]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [6]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_34 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [7]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [7]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [7]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [7]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [8]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [8]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [8]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [8]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_11 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [9]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [9]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\bank02/a1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\bank02/a1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [9]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [9]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/b0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/b0buso/gr7_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_21 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\rgf/bank02/gr01 [0]),
        .I2(\rgf/bank_sel [0]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_9 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [0]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [0]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_21_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_20 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\rgf/bank02/gr01 [1]),
        .I2(\rgf/bank_sel [0]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_8 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [1]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [1]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/b0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/b0buso/gr7_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/b0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/b0buso/gr7_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_11 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_21 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\rgf/bank02/gr01 [2]),
        .I2(\rgf/bank_sel [0]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [2]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [2]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_21_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [3]),
        .I1(\bank02/b0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [3]),
        .I3(\bank02/b0buso/gr7_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_21 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\rgf/bank02/gr01 [3]),
        .I2(\rgf/bank_sel [0]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_9 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [3]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [3]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_21_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/b0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/b0buso/gr7_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_11 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_24 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\rgf/bank02/gr01 [4]),
        .I2(\rgf/bank_sel [0]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [4]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [4]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_10 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [5]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [5]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_19 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_5 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/gr00 [5]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [5]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_9 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_10 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [6]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [6]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_19 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_5 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/gr00 [6]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [6]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_9 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_10 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [7]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [7]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_19 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_5 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/gr00 [7]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [7]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_10_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_9 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_17 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_41_n_0 ),
        .I1(\rgf/bank02/gr00 [10]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [10]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_42_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_41 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_42 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [10]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [10]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_69_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_69 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_69_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_17 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_18 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [11]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [11]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_45 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_7 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank02/gr00 [11]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [11]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_18 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_19 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [12]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [12]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_44_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_44 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_7 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank02/gr00 [12]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [12]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_18 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_19 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [13]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [13]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_45 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_7 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank02/gr00 [13]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [13]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_19 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_20 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [14]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [14]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_47_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_47 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_7 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/gr00 [14]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [14]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [14]));
  LUT5 #(
    .INIT(32'h00000100)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_193 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso/gr2_bus1 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_194 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_25 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_26 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_27 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_81_n_0 ),
        .I5(\bdatw[15]_INST_0_i_76_n_0 ),
        .O(\bank02/b0buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_28 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [15]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [15]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_84_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_78 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\bdatw[15]_INST_0_i_76_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank02/b0buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_79 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_189_n_0 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[8]_INST_0_i_5_n_0 ),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\bank02/b0buso/gr5_bus1 ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_82 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_83 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank02/b0buso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_84 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_9 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/gr00 [15]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [15]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_21 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_47_n_0 ),
        .I1(\rgf/bank02/gr00 [8]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [8]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_48_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_47 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_48 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [8]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [8]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_75_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_75 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_16 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank02/gr00 [9]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [9]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_39 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_40 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [9]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [9]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_67_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_67 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [0]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [0]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_13 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/b0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/b0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_14 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_22 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\rgf/bank02/gr21 [0]),
        .I2(\bdatw[15]_INST_0_i_123_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_11 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [1]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [1]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_21_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_12 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/b0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/b0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_13 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_21 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\rgf/bank02/gr21 [1]),
        .I2(\bdatw[15]_INST_0_i_123_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [2]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [2]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_13 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/b0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/b0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_14 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_22 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\rgf/bank02/gr21 [2]),
        .I2(\bdatw[15]_INST_0_i_123_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [3]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [3]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_13 
       (.I0(\rgf/bank02/gr20 [3]),
        .I1(\bank02/b0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [3]),
        .I3(\bank02/b0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_14 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_22 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\rgf/bank02/gr21 [3]),
        .I2(\bdatw[15]_INST_0_i_123_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [4]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [4]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_13 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/b0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/b0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_14 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_25 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\rgf/bank02/gr21 [4]),
        .I2(\bdatw[15]_INST_0_i_123_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_11 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [5]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [5]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_20 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_6 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/gr20 [5]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [5]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [6]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_20 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_6 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/gr20 [6]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [6]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [7]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_20 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_6 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/gr20 [7]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [7]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_16 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank02/gr20 [10]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [10]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_39 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_40 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [10]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_68 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_68_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_20 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [11]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_46 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_8 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/gr20 [11]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [11]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_20 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_21 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [12]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_45 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_8 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_20_n_0 ),
        .I1(\rgf/bank02/gr20 [12]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [12]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_21_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_20 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_21 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [13]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_46 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_8 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_20_n_0 ),
        .I1(\rgf/bank02/gr20 [13]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [13]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_21_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_21 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_22 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_48_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_48 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_8 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank02/gr20 [14]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [14]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_10 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/gr20 [15]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [15]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [15]));
  LUT5 #(
    .INIT(32'h00000400)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_195 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso2l/gr2_bus1 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_196 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso2l/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_30 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_31 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_81_n_0 ),
        .I5(\bdatw[15]_INST_0_i_76_n_0 ),
        .O(\bank02/b0buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_32 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_89_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_85 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\bdatw[15]_INST_0_i_76_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank02/b0buso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_86 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_189_n_0 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[8]_INST_0_i_5_n_0 ),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\bank02/b0buso2l/gr5_bus1 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_87 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank02/b0buso2l/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_88 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank02/b0buso2l/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_89 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_20 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_45_n_0 ),
        .I1(\rgf/bank02/gr20 [8]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [8]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_45 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_46 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [8]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_74_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_74 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_15 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank02/gr20 [9]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [9]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_38_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_37 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_38 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [9]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_66_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_66 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_11 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank02/gr00 [10]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [10]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_23 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_24 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [10]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [10]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_47_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_36 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_54_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_55_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_56_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_57_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_47 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_54 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_55 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_56 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_57 
       (.I0(\rgf/bank02/gr04 [2]),
        .I1(\bank02/b1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [2]),
        .I3(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_13 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/gr00 [11]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [11]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_30_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_30 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [11]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [11]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_51_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_42 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_58_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_59_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_60_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_61_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_51 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_58 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_59 
       (.I0(\rgf/bank02/gr00 [3]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [3]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_60 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_61 
       (.I0(\rgf/bank02/gr04 [3]),
        .I1(\bank02/b1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [3]),
        .I3(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_28_n_0 ),
        .I1(\rgf/bank02/gr00 [12]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [12]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_29_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_28 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_29 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [12]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [12]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_50_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_41 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_57_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_58_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_59_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_60_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_50 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_57 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_58 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_59 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_60 
       (.I0(\rgf/bank02/gr04 [4]),
        .I1(\bank02/b1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [4]),
        .I3(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_13 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/gr00 [13]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [13]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_30_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_30 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [13]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [13]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_51_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_42 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_58_n_0 ),
        .I1(\rgf/bank02/gr00 [5]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [5]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_59_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_51 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_58 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_59 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [5]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [5]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_68 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_13 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/gr00 [14]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [14]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_31 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_32 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [14]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [14]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_53_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_44 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_60_n_0 ),
        .I1(\rgf/bank02/gr00 [6]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [6]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_61_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_53 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_60 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_60_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_61 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [6]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [6]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_70_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_70 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_113 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_230_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_114 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_231_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_118 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_119 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_233_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_120 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_120_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_143 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_143_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_144 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [7]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [7]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_247_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_15 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_46_n_0 ),
        .I1(\rgf/bank02/gr00 [15]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [15]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_49_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_234 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_293_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_235 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_294_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_247 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_247_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_46 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_47 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_116_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_48 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\bdatw[15]_INST_0_i_39_n_0 ),
        .I5(ctl_selb1_rn[2]),
        .O(\bank02/b1buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_49 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [15]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [15]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_120_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_63 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_143_n_0 ),
        .I1(\rgf/bank02/gr00 [7]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [7]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_144_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_11 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/gr00 [8]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [8]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [8]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [8]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_53_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_38 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_60_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_61_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_62_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_63_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_53 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_60 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_61 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_62 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_63 
       (.I0(\rgf/bank02/gr04 [0]),
        .I1(\bank02/b1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [0]),
        .I3(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_10 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank02/gr00 [9]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [9]),
        .I4(\bank02/b1buso/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_21 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_22 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [9]),
        .I2(\bank02/b1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [9]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_33 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_51_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_52_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_53_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_54_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_45 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_51 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/b1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_52 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_53 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_54 
       (.I0(\rgf/bank02/gr04 [1]),
        .I1(\bank02/b1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [1]),
        .I3(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_12 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/gr20 [10]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [10]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_25 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_26 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [10]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_48_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_37 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_58_n_0 ),
        .I1(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_59_n_0 ),
        .I2(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_60_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_61_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_48 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_58 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_59 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_60 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_60_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_61 
       (.I0(\rgf/bank02/gr24 [2]),
        .I1(\bank02/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [2]),
        .I3(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_14 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/gr20 [11]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [11]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_31 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_32 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [11]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_52_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_62_n_0 ),
        .I1(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_63_n_0 ),
        .I2(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_64_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_65_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_52 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_62 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_63 
       (.I0(\rgf/bank02/gr20 [3]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [3]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_64 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_65 
       (.I0(\rgf/bank02/gr24 [3]),
        .I1(\bank02/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [3]),
        .I3(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/gr20 [12]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [12]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_31_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_30 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_31 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [12]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_51_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_42 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_61_n_0 ),
        .I1(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_62_n_0 ),
        .I2(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_63_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_64_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_51 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_61 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_62 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_63 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_64 
       (.I0(\rgf/bank02/gr24 [4]),
        .I1(\bank02/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [4]),
        .I3(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_14 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/gr20 [13]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [13]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_31 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_32 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [13]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_52_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_43 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_60_n_0 ),
        .I1(\rgf/bank02/gr20 [5]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [5]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_61_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_52 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_60 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_60_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_61 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [5]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [5]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_69_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_69 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/gr20 [14]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [14]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_34_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_34 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_54_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_45 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_62_n_0 ),
        .I1(\rgf/bank02/gr20 [6]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [6]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_63_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_54 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_62 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_63 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [6]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_71_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_71 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_121 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_230_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_122 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_231_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso2l/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_124 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso2l/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_125 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_233_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso2l/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_126 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_126_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_145 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_145_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_146 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [7]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_248_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_16 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_50_n_0 ),
        .I1(\rgf/bank02/gr20 [15]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [15]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_53_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_236 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_293_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso2l/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_237 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_294_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso2l/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_248 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_248_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_50 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_51 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_116_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank02/b1buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_52 
       (.I0(\bdatw[15]_INST_0_i_123_n_0 ),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\bdatw[15]_INST_0_i_39_n_0 ),
        .I5(ctl_selb1_rn[2]),
        .O(\bank02/b1buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_53 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_126_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_64 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_145_n_0 ),
        .I1(\rgf/bank02/gr20 [7]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [7]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_146_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_12 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_27_n_0 ),
        .I1(\rgf/bank02/gr20 [8]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [8]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_27 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_28 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [8]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_54_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_64_n_0 ),
        .I1(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_65_n_0 ),
        .I2(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_66_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_67_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_54 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_64 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_65 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_65_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_66 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_67 
       (.I0(\rgf/bank02/gr24 [0]),
        .I1(\bank02/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [0]),
        .I3(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_11 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank02/gr20 [9]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [9]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\bank02/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [9]),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_34 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_55_n_0 ),
        .I1(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_56_n_0 ),
        .I2(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_57_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_58_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_46 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_55 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_56 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_57 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\bank02/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\bank02/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_58 
       (.I0(\rgf/bank02/gr24 [1]),
        .I1(\bank02/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [1]),
        .I3(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/bbus_o[0]_INST_0_i_5 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_14_n_0 ),
        .O(\rgf/b0bus_b02 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/bbus_o[1]_INST_0_i_4 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10_n_0 ),
        .I3(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_11_n_0 ),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_12_n_0 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_13_n_0 ),
        .O(\rgf/b0bus_b02 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/bbus_o[2]_INST_0_i_5 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_14_n_0 ),
        .O(\rgf/b0bus_b02 [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/bbus_o[3]_INST_0_i_5 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_14_n_0 ),
        .O(\rgf/b0bus_b02 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/bbus_o[4]_INST_0_i_5 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_13_n_0 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_14_n_0 ),
        .O(\rgf/b0bus_b02 [4]));
  FDRE \rgf/bank02/grn00/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [0]),
        .Q(\rgf/bank02/gr00 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [10]),
        .Q(\rgf/bank02/gr00 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [11]),
        .Q(\rgf/bank02/gr00 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [12]),
        .Q(\rgf/bank02/gr00 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [13]),
        .Q(\rgf/bank02/gr00 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [14]),
        .Q(\rgf/bank02/gr00 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [15]),
        .Q(\rgf/bank02/gr00 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [1]),
        .Q(\rgf/bank02/gr00 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [2]),
        .Q(\rgf/bank02/gr00 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [3]),
        .Q(\rgf/bank02/gr00 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [4]),
        .Q(\rgf/bank02/gr00 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [5]),
        .Q(\rgf/bank02/gr00 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [6]),
        .Q(\rgf/bank02/gr00 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [7]),
        .Q(\rgf/bank02/gr00 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [8]),
        .Q(\rgf/bank02/gr00 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn00/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [9]),
        .Q(\rgf/bank02/gr00 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr01 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn01/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\bank02/grn01/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr01 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr02 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn02/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\bank02/grn02/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr02 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr03 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn03/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\bank02/grn03/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr03 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr04 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn04/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\bank02/grn04/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr04 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr05 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn05/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\bank02/grn05/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr05 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr06 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn06/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\bank02/grn06/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr06 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr07 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn07/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\bank02/grn07/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr07 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr20 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn20/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\bank02/grn20/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr20 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr21 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn21/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\bank02/grn21/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr21 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr22 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn22/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\bank02/grn22/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr22 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr23 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn23/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\bank02/grn23/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr23 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr24 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn24/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\bank02/grn24/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr24 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr25 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn25/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\bank02/grn25/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr25 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr26 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn26/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\bank02/grn26/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr26 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank02/gr27 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank02/grn27/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\bank02/grn27/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank02/gr27 [9]),
        .R(\rgf/treg/p_0_in ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [0]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [0]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [0]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [0]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [0]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [0]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [0]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [0]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [10]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [10]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [10]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [10]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [11]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [11]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [11]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [11]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [12]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [12]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [12]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [12]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [13]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [13]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [13]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [13]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [14]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [14]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [14]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [14]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_100 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(ctl_sela0_rn[0]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_101 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela0_rn[2]),
        .I3(ctl_sela0_rn[0]),
        .I4(\badr[15]_INST_0_i_28_n_0 ),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_29 
       (.I0(\rgf/bank13/gr04 [15]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [15]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_30 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_31 
       (.I0(\rgf/bank13/gr00 [15]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [15]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_32 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_94 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_95 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_96 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_97 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_98 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_99 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\badr[15]_INST_0_i_191_n_0 ),
        .I5(ctl_sela0_rn[2]),
        .O(\bank13/a0buso/gr7_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [1]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [1]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [1]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [1]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [1]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [1]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [1]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [1]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [2]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [2]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [2]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [2]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [2]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [2]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [2]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [2]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [3]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [3]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [3]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [3]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [3]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [3]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [3]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [3]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [4]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [4]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [4]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [4]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [4]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [4]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [4]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [4]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [5]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [5]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [5]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [5]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [5]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [5]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [6]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [6]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [6]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [6]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [7]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [7]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [7]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [7]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [8]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [8]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [8]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [8]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [9]),
        .I1(\bank13/a0buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [9]),
        .I3(\bank13/a0buso/gr3_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_24 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\bank13/a0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\bank13/a0buso/gr1_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_25 
       (.I0(\rgf/bank13/gr00 [9]),
        .I1(\bank13/a0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [9]),
        .I3(\bank13/a0buso/gr7_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\bank13/a0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\bank13/a0buso/gr5_bus1 ),
        .O(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_37 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\rgf_c0bus_wb[12]_i_39_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_40_n_0 ),
        .O(\rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_38 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\rgf_c0bus_wb[12]_i_41_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_42_n_0 ),
        .O(\rgf/bank13/a0buso/i_/rgf_c0bus_wb[12]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\badr[0]_INST_0_i_44_n_0 ),
        .I5(\badr[0]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\badr[0]_INST_0_i_46_n_0 ),
        .I5(\badr[0]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\badr[10]_INST_0_i_43_n_0 ),
        .I5(\badr[10]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\badr[10]_INST_0_i_45_n_0 ),
        .I5(\badr[10]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\badr[11]_INST_0_i_44_n_0 ),
        .I5(\badr[11]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\badr[11]_INST_0_i_46_n_0 ),
        .I5(\badr[11]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\badr[12]_INST_0_i_43_n_0 ),
        .I5(\badr[12]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\badr[12]_INST_0_i_45_n_0 ),
        .I5(\badr[12]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\badr[13]_INST_0_i_43_n_0 ),
        .I5(\badr[13]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\badr[13]_INST_0_i_45_n_0 ),
        .I5(\badr[13]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\badr[14]_INST_0_i_43_n_0 ),
        .I5(\badr[14]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\badr[14]_INST_0_i_45_n_0 ),
        .I5(\badr[14]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_102 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso2l/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_103 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(ctl_sela0_rn[0]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_106 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\badr[15]_INST_0_i_191_n_0 ),
        .I5(ctl_sela0_rn[2]),
        .O(\bank13/a0buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_107 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(ctl_sela0_rn[2]),
        .I5(\badr[15]_INST_0_i_191_n_0 ),
        .O(\bank13/a0buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_33 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\badr[15]_INST_0_i_104_n_0 ),
        .I5(\badr[15]_INST_0_i_105_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_34 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\badr[15]_INST_0_i_108_n_0 ),
        .I5(\badr[15]_INST_0_i_109_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\badr[1]_INST_0_i_43_n_0 ),
        .I5(\badr[1]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\badr[1]_INST_0_i_45_n_0 ),
        .I5(\badr[1]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\badr[2]_INST_0_i_43_n_0 ),
        .I5(\badr[2]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\badr[2]_INST_0_i_45_n_0 ),
        .I5(\badr[2]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\badr[3]_INST_0_i_44_n_0 ),
        .I5(\badr[3]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\badr[3]_INST_0_i_46_n_0 ),
        .I5(\badr[3]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\badr[4]_INST_0_i_43_n_0 ),
        .I5(\badr[4]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\badr[4]_INST_0_i_45_n_0 ),
        .I5(\badr[4]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\badr[5]_INST_0_i_43_n_0 ),
        .I5(\badr[5]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\badr[5]_INST_0_i_45_n_0 ),
        .I5(\badr[5]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\badr[6]_INST_0_i_43_n_0 ),
        .I5(\badr[6]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\badr[6]_INST_0_i_45_n_0 ),
        .I5(\badr[6]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\badr[7]_INST_0_i_44_n_0 ),
        .I5(\badr[7]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\badr[7]_INST_0_i_46_n_0 ),
        .I5(\badr[7]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\badr[8]_INST_0_i_43_n_0 ),
        .I5(\badr[8]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\badr[8]_INST_0_i_45_n_0 ),
        .I5(\badr[8]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_27 
       (.I0(\bank13/a0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/a0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\badr[9]_INST_0_i_43_n_0 ),
        .I5(\badr[9]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_28 
       (.I0(\bank13/a0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/a0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\badr[9]_INST_0_i_45_n_0 ),
        .I5(\badr[9]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_38 
       (.I0(\rgf/bank13/gr04 [0]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [0]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_39 
       (.I0(\rgf/bank13/gr02 [0]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [0]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_40 
       (.I0(\rgf/bank13/gr00 [0]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [0]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_41 
       (.I0(\rgf/bank13/gr06 [0]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [0]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [10]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [10]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [10]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [10]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_38 
       (.I0(\rgf/bank13/gr04 [11]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [11]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_39 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_40 
       (.I0(\rgf/bank13/gr00 [11]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [11]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_41 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [12]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [12]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [12]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [12]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [13]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [13]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [13]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [13]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [14]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [14]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [14]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [14]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_149 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(ctl_sela1_rn),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_150 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_151 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_152 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_153 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_154 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_235_n_0 ),
        .I5(\badr[15]_INST_0_i_40_n_0 ),
        .O(\bank13/a1buso/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_155 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(ctl_sela1_rn),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_156 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_40_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_52_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_53 
       (.I0(\rgf/bank13/gr04 [15]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [15]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_54 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_55 
       (.I0(\rgf/bank13/gr00 [15]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [15]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_56 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [1]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [1]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [1]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [1]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [1]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [1]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [1]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [1]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [2]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [2]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [2]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [2]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [2]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [2]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [2]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [2]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_38 
       (.I0(\rgf/bank13/gr04 [3]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [3]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_39 
       (.I0(\rgf/bank13/gr02 [3]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [3]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_40 
       (.I0(\rgf/bank13/gr00 [3]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [3]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41 
       (.I0(\rgf/bank13/gr06 [3]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [3]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [4]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [4]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [4]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [4]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [4]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [4]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [4]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [4]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [5]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [5]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [5]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [5]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [5]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [5]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [6]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [6]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [6]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [6]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_38 
       (.I0(\rgf/bank13/gr04 [7]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [7]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_39 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_40 
       (.I0(\rgf/bank13/gr00 [7]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [7]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_41 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [8]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [8]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [8]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [8]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_37 
       (.I0(\rgf/bank13/gr04 [9]),
        .I1(\bank13/a1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr03 [9]),
        .I3(\bank13/a1buso/gr3_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\bank13/a1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\bank13/a1buso/gr1_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_39 
       (.I0(\rgf/bank13/gr00 [9]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [9]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_40 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_26 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\rgf_c1bus_wb[10]_i_28_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_29_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_27 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\rgf_c1bus_wb[10]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_31_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\badr[0]_INST_0_i_49_n_0 ),
        .I5(\badr[0]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\badr[0]_INST_0_i_51_n_0 ),
        .I5(\badr[0]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\badr[10]_INST_0_i_47_n_0 ),
        .I5(\badr[10]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\badr[10]_INST_0_i_49_n_0 ),
        .I5(\badr[10]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\badr[11]_INST_0_i_52_n_0 ),
        .I5(\badr[11]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_43 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\badr[11]_INST_0_i_54_n_0 ),
        .I5(\badr[11]_INST_0_i_55_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\badr[12]_INST_0_i_47_n_0 ),
        .I5(\badr[12]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\badr[12]_INST_0_i_49_n_0 ),
        .I5(\badr[12]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\badr[13]_INST_0_i_47_n_0 ),
        .I5(\badr[13]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\badr[13]_INST_0_i_49_n_0 ),
        .I5(\badr[13]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\badr[14]_INST_0_i_47_n_0 ),
        .I5(\badr[14]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\badr[14]_INST_0_i_49_n_0 ),
        .I5(\badr[14]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_157 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso2l/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_158 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(ctl_sela1_rn),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_161 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_235_n_0 ),
        .I5(\badr[15]_INST_0_i_40_n_0 ),
        .O(\bank13/a1buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_162 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\badr[15]_INST_0_i_40_n_0 ),
        .I5(\badr[15]_INST_0_i_235_n_0 ),
        .O(\bank13/a1buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_57 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\badr[15]_INST_0_i_159_n_0 ),
        .I5(\badr[15]_INST_0_i_160_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_58 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\badr[15]_INST_0_i_163_n_0 ),
        .I5(\badr[15]_INST_0_i_164_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\badr[1]_INST_0_i_47_n_0 ),
        .I5(\badr[1]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\badr[1]_INST_0_i_49_n_0 ),
        .I5(\badr[1]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\badr[2]_INST_0_i_47_n_0 ),
        .I5(\badr[2]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\badr[2]_INST_0_i_49_n_0 ),
        .I5(\badr[2]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\badr[3]_INST_0_i_51_n_0 ),
        .I5(\badr[3]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_43 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\badr[3]_INST_0_i_53_n_0 ),
        .I5(\badr[3]_INST_0_i_54_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\badr[4]_INST_0_i_47_n_0 ),
        .I5(\badr[4]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\badr[4]_INST_0_i_49_n_0 ),
        .I5(\badr[4]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\badr[5]_INST_0_i_47_n_0 ),
        .I5(\badr[5]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\badr[5]_INST_0_i_49_n_0 ),
        .I5(\badr[5]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\badr[6]_INST_0_i_47_n_0 ),
        .I5(\badr[6]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\badr[6]_INST_0_i_49_n_0 ),
        .I5(\badr[6]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\badr[7]_INST_0_i_52_n_0 ),
        .I5(\badr[7]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_43 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\badr[7]_INST_0_i_54_n_0 ),
        .I5(\badr[7]_INST_0_i_55_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\badr[8]_INST_0_i_47_n_0 ),
        .I5(\badr[8]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\badr[8]_INST_0_i_49_n_0 ),
        .I5(\badr[8]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_41 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\badr[9]_INST_0_i_47_n_0 ),
        .I5(\badr[9]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_42 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\badr[9]_INST_0_i_49_n_0 ),
        .I5(\badr[9]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18 
       (.I0(\rgf/bank13/gr06 [0]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [0]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19 
       (.I0(\rgf/bank13/gr00 [0]),
        .I1(\bank13/b0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [0]),
        .I3(\bank13/b0buso/gr7_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_20 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [0]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [0]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26 
       (.I0(\rgf/bank13/gr02 [0]),
        .I1(\rgf/bank13/gr01 [0]),
        .I2(\bdatw[15]_INST_0_i_238_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_17 
       (.I0(\rgf/bank13/gr06 [1]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [1]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_18 
       (.I0(\rgf/bank13/gr00 [1]),
        .I1(\bank13/b0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [1]),
        .I3(\bank13/b0buso/gr7_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_19 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [1]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [1]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_25_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_25 
       (.I0(\rgf/bank13/gr02 [1]),
        .I1(\rgf/bank13/gr01 [1]),
        .I2(\bdatw[15]_INST_0_i_238_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_18 
       (.I0(\rgf/bank13/gr06 [2]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [2]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_19 
       (.I0(\rgf/bank13/gr00 [2]),
        .I1(\bank13/b0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [2]),
        .I3(\bank13/b0buso/gr7_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_20 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [2]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [2]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_26 
       (.I0(\rgf/bank13/gr02 [2]),
        .I1(\rgf/bank13/gr01 [2]),
        .I2(\bdatw[15]_INST_0_i_238_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_18 
       (.I0(\rgf/bank13/gr06 [3]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [3]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_19 
       (.I0(\rgf/bank13/gr00 [3]),
        .I1(\bank13/b0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [3]),
        .I3(\bank13/b0buso/gr7_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_20 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [3]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [3]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_26 
       (.I0(\rgf/bank13/gr02 [3]),
        .I1(\rgf/bank13/gr01 [3]),
        .I2(\bdatw[15]_INST_0_i_238_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_18 
       (.I0(\rgf/bank13/gr06 [4]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [4]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_19 
       (.I0(\rgf/bank13/gr00 [4]),
        .I1(\bank13/b0buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [4]),
        .I3(\bank13/b0buso/gr7_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_20 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [4]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [4]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_32_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004000)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_30 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\bdatw[15]_INST_0_i_76_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank13/b0buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_31 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_189_n_0 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[8]_INST_0_i_5_n_0 ),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\bank13/b0buso/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_32 
       (.I0(\rgf/bank13/gr02 [4]),
        .I1(\rgf/bank13/gr01 [4]),
        .I2(\bdatw[15]_INST_0_i_238_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_14 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [5]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [5]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_15 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [5]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [5]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [5]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [5]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_14 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [6]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [6]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [6]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [6]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_22 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_14 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [7]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [7]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [7]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [7]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_22 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_19 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_43_n_0 ),
        .I1(\rgf/bank13/gr00 [10]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [10]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_43 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_44 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [10]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [10]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_70_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_70 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_22 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [11]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [11]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_23 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [11]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [11]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_48 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_23 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [12]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [12]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_24 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [12]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [12]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_46 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_47 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_23 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [13]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [13]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_24 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [13]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [13]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_47 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_48 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_24 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [14]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [14]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_49_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_25 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [14]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [14]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_49 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_50 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_197 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso/gr2_bus1 ));
  LUT5 #(
    .INIT(32'h00000400)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_198 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso/gr1_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_34 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_92_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_35 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_95_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_90 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_91 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank13/b0buso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_92 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h0000400000000000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_93 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_81_n_0 ),
        .I5(\bdatw[15]_INST_0_i_76_n_0 ),
        .O(\bank13/b0buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_94 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_95 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_95_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_23 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_49_n_0 ),
        .I1(\rgf/bank13/gr00 [8]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [8]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_49 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_50 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [8]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [8]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_76_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_76 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_18 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_41_n_0 ),
        .I1(\rgf/bank13/gr00 [9]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [9]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_41 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_42 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [9]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [9]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_68 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bbus_o[0]_INST_0_i_23_n_0 ),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [0]),
        .I5(\bbus_o[0]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_17 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_25_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_25 
       (.I0(\rgf/bank13/gr22 [0]),
        .I1(\rgf/bank13/gr21 [0]),
        .I2(\rgf/bank_sel [3]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_15 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bbus_o[1]_INST_0_i_22_n_0 ),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [1]),
        .I5(\bbus_o[1]_INST_0_i_23_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_24 
       (.I0(\rgf/bank13/gr22 [1]),
        .I1(\rgf/bank13/gr21 [1]),
        .I2(\rgf/bank_sel [3]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bbus_o[2]_INST_0_i_23_n_0 ),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [2]),
        .I5(\bbus_o[2]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_17 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_25_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_25 
       (.I0(\rgf/bank13/gr22 [2]),
        .I1(\rgf/bank13/gr21 [2]),
        .I2(\rgf/bank_sel [3]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bbus_o[3]_INST_0_i_23_n_0 ),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [3]),
        .I5(\bbus_o[3]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_17 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_25_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_25 
       (.I0(\rgf/bank13/gr22 [3]),
        .I1(\rgf/bank13/gr21 [3]),
        .I2(\rgf/bank_sel [3]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bbus_o[4]_INST_0_i_26_n_0 ),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [4]),
        .I5(\bbus_o[4]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_17 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_27 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_189_n_0 ),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[8]_INST_0_i_5_n_0 ),
        .I4(\bdatw[15]_INST_0_i_19_n_0 ),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\bank13/b0buso2l/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_29 
       (.I0(\rgf/bank13/gr22 [4]),
        .I1(\rgf/bank13/gr21 [4]),
        .I2(\rgf/bank_sel [3]),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_23_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_17 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_23 
       (.I0(\rgf/bank13/gr22 [5]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [5]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [5]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [5]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_23_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_23 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [6]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [6]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_16 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_23_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_23 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [7]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [7]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_20 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_45_n_0 ),
        .I1(\rgf/bank13/gr20 [10]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [10]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_45 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [10]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_46 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_71_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_71 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [10]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_71_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_24 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_49_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_25 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_49 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [11]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_50 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [11]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_25 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_26 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_49_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_48 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [12]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_49 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [12]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_25 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_49_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_26 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_49 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [13]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_50 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [13]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_26 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_51_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_27 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_51 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [14]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_52 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [14]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_100 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso2l/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_101 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [15]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_101_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_199 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[0]),
        .I3(ctl_selb0_rn[1]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso2l/gr2_bus1 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_200 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso2l/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_201 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\bdatw[15]_INST_0_i_76_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank13/b0buso2l/gr6_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_36 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_98_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_37 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_101_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_96 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_80_n_0 ),
        .O(\bank13/b0buso2l/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_97 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(\bdatw[15]_INST_0_i_76_n_0 ),
        .I4(ctl_selb0_rn[0]),
        .I5(\bdatw[15]_INST_0_i_81_n_0 ),
        .O(\bank13/b0buso2l/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_98 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [15]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_99 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(ctl_selb0_rn[1]),
        .I3(ctl_selb0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_81_n_0 ),
        .I5(\bdatw[15]_INST_0_i_76_n_0 ),
        .O(\bank13/b0buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_24 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_51_n_0 ),
        .I1(\rgf/bank13/gr20 [8]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [8]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_51 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [8]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_52 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_77_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_77 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [8]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_19 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_43_n_0 ),
        .I1(\rgf/bank13/gr20 [9]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [9]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_43 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [9]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_44 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_69_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_69 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [9]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_69_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_28 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [10]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [10]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_49_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_29 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [10]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [10]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_49 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_50 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_63 
       (.I0(\bdatw[10]_INST_0_i_72_n_0 ),
        .I1(\bdatw[10]_INST_0_i_73_n_0 ),
        .I2(\bank13/b1buso/gr1_bus1 ),
        .I3(\rgf/bank13/gr01 [2]),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [2]),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_64 
       (.I0(\bdatw[10]_INST_0_i_74_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [2]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .I4(\rgf/bank13/gr05 [2]),
        .I5(\bdatw[10]_INST_0_i_75_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_34 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [11]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [11]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_35 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [11]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [11]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_54_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_53 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_54 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_67 
       (.I0(\bdatw[11]_INST_0_i_72_n_0 ),
        .I1(\bdatw[11]_INST_0_i_73_n_0 ),
        .I2(\bank13/b1buso/gr1_bus1 ),
        .I3(\rgf/bank13/gr01 [3]),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [3]),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_68 
       (.I0(\bdatw[11]_INST_0_i_74_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [3]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .I4(\rgf/bank13/gr05 [3]),
        .I5(\bdatw[11]_INST_0_i_75_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_68_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_33 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [12]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [12]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_34 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [12]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [12]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_52 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_52_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_53 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_66 
       (.I0(\bdatw[12]_INST_0_i_71_n_0 ),
        .I1(\bdatw[12]_INST_0_i_72_n_0 ),
        .I2(\bank13/b1buso/gr1_bus1 ),
        .I3(\rgf/bank13/gr01 [4]),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [4]),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_67 
       (.I0(\bdatw[12]_INST_0_i_73_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [4]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .I4(\rgf/bank13/gr05 [4]),
        .I5(\bdatw[12]_INST_0_i_74_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_34 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [13]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [13]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_35 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [13]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [13]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_54_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_53 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_54 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_54_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_63 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [5]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [5]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_70_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_63_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_64 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [5]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [5]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_71_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_70 
       (.I0(\rgf/bank13/gr02 [5]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [5]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_70_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_71 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_71_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_36 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [14]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [14]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_55_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [14]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [14]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_56_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_55 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_56 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_65 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [6]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [6]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_72_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_65_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_66 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [6]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [6]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_73_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_72 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_72_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_73 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_130 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_131 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_233_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_132 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_133 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\bdatw[15]_INST_0_i_39_n_0 ),
        .I5(ctl_selb1_rn[2]),
        .O(\bank13/b1buso/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_134 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_116_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_135 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_135_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_148 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [7]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [7]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_249_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_148_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_149 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [7]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [7]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_250_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_239 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_293_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_240 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_294_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_241 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_230_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_242 
       (.I0(\bdatw[15]_INST_0_i_238_n_0 ),
        .I1(\bdatw[15]_INST_0_i_231_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_249 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_249_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_250 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_250_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_55 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_132_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_55_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_56 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_135_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_30 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [8]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [8]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_55_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_31 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [8]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [8]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_56_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_55 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_56 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_69 
       (.I0(\bdatw[8]_INST_0_i_78_n_0 ),
        .I1(\bdatw[8]_INST_0_i_79_n_0 ),
        .I2(\bank13/b1buso/gr1_bus1 ),
        .I3(\rgf/bank13/gr01 [0]),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [0]),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_70 
       (.I0(\bdatw[8]_INST_0_i_80_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [0]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .I4(\rgf/bank13/gr05 [0]),
        .I5(\bdatw[8]_INST_0_i_81_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_26 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [9]),
        .I2(\bank13/b1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [9]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27 
       (.I0(\bank13/b1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [9]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [9]),
        .I4(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_47 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\bank13/b1buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\bank13/b1buso/gr1_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_48 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\bank13/b1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_60 
       (.I0(\bdatw[9]_INST_0_i_70_n_0 ),
        .I1(\bdatw[9]_INST_0_i_71_n_0 ),
        .I2(\bank13/b1buso/gr1_bus1 ),
        .I3(\rgf/bank13/gr01 [1]),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_61 
       (.I0(\bdatw[9]_INST_0_i_72_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [1]),
        .I3(\bank13/b1buso/gr5_bus1 ),
        .I4(\rgf/bank13/gr05 [1]),
        .I5(\bdatw[9]_INST_0_i_73_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_61_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_30 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_51_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_31 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_51 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [10]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_52 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [10]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_65 
       (.I0(\bdatw[10]_INST_0_i_76_n_0 ),
        .I1(\bdatw[10]_INST_0_i_77_n_0 ),
        .I2(\bank13/b1buso2l/gr1_bus1 ),
        .I3(\rgf/bank13/gr21 [2]),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [2]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_66 
       (.I0(\bdatw[10]_INST_0_i_78_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [2]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [2]),
        .I5(\bdatw[10]_INST_0_i_79_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_66_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_36 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_55_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_37 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_56_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_55 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [11]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_56 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [11]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_69 
       (.I0(\bdatw[11]_INST_0_i_76_n_0 ),
        .I1(\bdatw[11]_INST_0_i_77_n_0 ),
        .I2(\bank13/b1buso2l/gr1_bus1 ),
        .I3(\rgf/bank13/gr21 [3]),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [3]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_70 
       (.I0(\bdatw[11]_INST_0_i_78_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [3]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [3]),
        .I5(\bdatw[11]_INST_0_i_79_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_35 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_54_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_36 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_55_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_54 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [12]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_55 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [12]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_68 
       (.I0(\bdatw[12]_INST_0_i_75_n_0 ),
        .I1(\bdatw[12]_INST_0_i_76_n_0 ),
        .I2(\bank13/b1buso2l/gr1_bus1 ),
        .I3(\rgf/bank13/gr21 [4]),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [4]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_69 
       (.I0(\bdatw[12]_INST_0_i_77_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [4]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [4]),
        .I5(\bdatw[12]_INST_0_i_78_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_69_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_36 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_55_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_37 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_56_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_55 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [13]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_56 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [13]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_65 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_72_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_65_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_66 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_73_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_72 
       (.I0(\rgf/bank13/gr22 [5]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [5]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_72_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_73 
       (.I0(\rgf/bank13/gr26 [5]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [5]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_73_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_57_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_39 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_58_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_57 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [14]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_58 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [14]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_67 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_74_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_68 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_75_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_68_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_74 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [6]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_74_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_75 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [6]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_136 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso2l/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_137 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_233_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso2l/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_138 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [15]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_138_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_139 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_117_n_0 ),
        .I2(\bdatw[15]_INST_0_i_40_n_0 ),
        .I3(ctl_selb1_0),
        .I4(\bdatw[15]_INST_0_i_39_n_0 ),
        .I5(ctl_selb1_rn[2]),
        .O(\bank13/b1buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_140 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_116_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso2l/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_141 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [15]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_141_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_150 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_251_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_150_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_151 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_252_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_243 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_293_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso2l/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_244 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_294_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso2l/gr1_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_245 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_230_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_246 
       (.I0(\rgf/bank_sel [3]),
        .I1(\bdatw[15]_INST_0_i_231_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[15]_INST_0_i_40_n_0 ),
        .I4(ctl_selb1_0),
        .I5(\bdatw[15]_INST_0_i_39_n_0 ),
        .O(\bank13/b1buso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_251 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [7]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_251_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_252 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [7]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_252_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_57 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_138_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_57_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_58 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_141_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_32 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_57_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_33 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_58_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_57 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [8]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_58 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [8]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_71 
       (.I0(\bdatw[8]_INST_0_i_82_n_0 ),
        .I1(\bdatw[8]_INST_0_i_83_n_0 ),
        .I2(\bank13/b1buso2l/gr1_bus1 ),
        .I3(\rgf/bank13/gr21 [0]),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [0]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_72 
       (.I0(\bdatw[8]_INST_0_i_84_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [0]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [0]),
        .I5(\bdatw[8]_INST_0_i_85_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_72_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_28 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/b1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_49_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29 
       (.I0(\bank13/b1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_49 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\bank13/b1buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [9]),
        .I3(\bank13/b1buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_50 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\bank13/b1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [9]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_62 
       (.I0(\bdatw[9]_INST_0_i_74_n_0 ),
        .I1(\bdatw[9]_INST_0_i_75_n_0 ),
        .I2(\bank13/b1buso2l/gr1_bus1 ),
        .I3(\rgf/bank13/gr21 [1]),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_63 
       (.I0(\bdatw[9]_INST_0_i_76_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [1]),
        .I3(\bank13/b1buso2l/gr5_bus1 ),
        .I4(\rgf/bank13/gr25 [1]),
        .I5(\bdatw[9]_INST_0_i_77_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[0]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_42_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43_n_0 ),
        .O(\rgf/a1bus_b13 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[0]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[10]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[10]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[11]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_42_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_43_n_0 ),
        .O(\rgf/a1bus_b13 [11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[11]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[12]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[12]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[13]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[13]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[14]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[14]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[15]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_53_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_54_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_55_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_56_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_57_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_58_n_0 ),
        .O(\rgf/a1bus_b13 [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[15]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_32_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_33_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_34_n_0 ),
        .O(\rgf/a0bus_b13 [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[1]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[1]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[2]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[2]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[3]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_43_n_0 ),
        .O(\rgf/a1bus_b13 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[3]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[4]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[4]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[5]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[5]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[6]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[6]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[7]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_42_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_43_n_0 ),
        .O(\rgf/a1bus_b13 [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[7]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[8]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[8]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[9]_INST_0_i_13 
       (.I0(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_42_n_0 ),
        .O(\rgf/a1bus_b13 [9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[9]_INST_0_i_7 
       (.I0(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_28_n_0 ),
        .O(\rgf/a0bus_b13 [9]));
  FDRE \rgf/bank13/grn00/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr00 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn00/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\bank13/grn00/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr00 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr01 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn01/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\bank13/grn01/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr01 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr02 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn02/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\bank13/grn02/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr02 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr03 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn03/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\bank13/grn03/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr03 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr04 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn04/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\bank13/grn04/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr04 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr05 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn05/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\bank13/grn05/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr05 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr06 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn06/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\bank13/grn06/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr06 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr07 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn07/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\bank13/grn07/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr07 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr20 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn20/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\bank13/grn20/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr20 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr21 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn21/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\bank13/grn21/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr21 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr22 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn22/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\bank13/grn22/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr22 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr23 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn23/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\bank13/grn23/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr23 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr24 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn24/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\bank13/grn24/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr24 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr25 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn25/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\bank13/grn25/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr25 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr26 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn26/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\bank13/grn26/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr26 [9]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[0]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [0]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[10]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [10]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[11]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [11]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[12]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [12]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[13]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [13]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[14]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [14]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[15]_i_2_n_0 ),
        .Q(\rgf/bank13/gr27 [15]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[1]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [1]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[2]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [2]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[3]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [3]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[4]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [4]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[5]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [5]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[6]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [6]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[7]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [7]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[8]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [8]),
        .R(\rgf/treg/p_0_in ));
  FDRE \rgf/bank13/grn27/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\bank13/grn27/grn[9]_i_1_n_0 ),
        .Q(\rgf/bank13/gr27 [9]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [0]),
        .Q(\rgf/ivec/iv [0]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [10]),
        .Q(\rgf/ivec/iv [10]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [11]),
        .Q(\rgf/ivec/iv [11]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [12]),
        .Q(\rgf/ivec/iv [12]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [13]),
        .Q(\rgf/ivec/iv [13]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [14]),
        .Q(\rgf/ivec/iv [14]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [15]),
        .Q(\rgf/ivec/iv [15]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [1]),
        .Q(\rgf/ivec/iv [1]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [2]),
        .Q(\rgf/ivec/iv [2]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [3]),
        .Q(\rgf/ivec/iv [3]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [4]),
        .Q(\rgf/ivec/iv [4]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [5]),
        .Q(\rgf/ivec/iv [5]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [6]),
        .Q(\rgf/ivec/iv [6]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [7]),
        .Q(\rgf/ivec/iv [7]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [8]),
        .Q(\rgf/ivec/iv [8]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [9]),
        .Q(\rgf/ivec/iv [9]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [0]),
        .Q(\rgf/pcnt/pc [0]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [10]),
        .Q(\rgf/pcnt/pc [10]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [11]),
        .Q(\rgf/pcnt/pc [11]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [12]),
        .Q(\rgf/pcnt/pc [12]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [13]),
        .Q(\rgf/pcnt/pc [13]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [14]),
        .Q(\rgf/pcnt/pc [14]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [15]),
        .Q(\rgf/pcnt/pc [15]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [1]),
        .Q(\rgf/pcnt/pc [1]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [2]),
        .Q(\rgf/pcnt/pc [2]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [3]),
        .Q(\rgf/pcnt/pc [3]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [4]),
        .Q(\rgf/pcnt/pc [4]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [5]),
        .Q(\rgf/pcnt/pc [5]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [6]),
        .Q(\rgf/pcnt/pc [6]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [7]),
        .Q(\rgf/pcnt/pc [7]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [8]),
        .Q(\rgf/pcnt/pc [8]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [9]),
        .Q(\rgf/pcnt/pc [9]),
        .R(\rgf/treg/p_0_in ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf/rctl/badr[15]_INST_0_i_209 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .O(\rgf/bank_sel [3]));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf/rctl/bdatw[15]_INST_0_i_115 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [1]),
        .O(\rgf/bank_sel [0]));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[0]),
        .Q(\rgf/rctl/rgf_c0bus_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[10] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[10]),
        .Q(\rgf/rctl/rgf_c0bus_wb [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[11] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[11]),
        .Q(\rgf/rctl/rgf_c0bus_wb [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[12] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[12]),
        .Q(\rgf/rctl/rgf_c0bus_wb [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[13] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[13]),
        .Q(\rgf/rctl/rgf_c0bus_wb [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[14] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[14]),
        .Q(\rgf/rctl/rgf_c0bus_wb [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[15] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[15]),
        .Q(\rgf/rctl/rgf_c0bus_wb [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[1]),
        .Q(\rgf/rctl/rgf_c0bus_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[2]),
        .Q(\rgf/rctl/rgf_c0bus_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[3] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[3]),
        .Q(\rgf/rctl/rgf_c0bus_wb [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[4] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[4]),
        .Q(\rgf/rctl/rgf_c0bus_wb [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[5] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[5]),
        .Q(\rgf/rctl/rgf_c0bus_wb [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[6] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[6]),
        .Q(\rgf/rctl/rgf_c0bus_wb [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[7] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[7]),
        .Q(\rgf/rctl/rgf_c0bus_wb [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[8] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[8]),
        .Q(\rgf/rctl/rgf_c0bus_wb [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[9] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[9]),
        .Q(\rgf/rctl/rgf_c0bus_wb [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[0]),
        .Q(\rgf/rctl/rgf_c1bus_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[10] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[10]),
        .Q(\rgf/rctl/rgf_c1bus_wb [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[11] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[11]),
        .Q(\rgf/rctl/rgf_c1bus_wb [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[12] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[12]),
        .Q(\rgf/rctl/rgf_c1bus_wb [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[13] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[13]),
        .Q(\rgf/rctl/rgf_c1bus_wb [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[14] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[14]),
        .Q(\rgf/rctl/rgf_c1bus_wb [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[15] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[15]),
        .Q(\rgf/rctl/rgf_c1bus_wb [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[1]),
        .Q(\rgf/rctl/rgf_c1bus_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[2]),
        .Q(\rgf/rctl/rgf_c1bus_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[3] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[3]),
        .Q(\rgf/rctl/rgf_c1bus_wb [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[4] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[4]),
        .Q(\rgf/rctl/rgf_c1bus_wb [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[5] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[5]),
        .Q(\rgf/rctl/rgf_c1bus_wb [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[6] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[6]),
        .Q(\rgf/rctl/rgf_c1bus_wb [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[7] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[7]),
        .Q(\rgf/rctl/rgf_c1bus_wb [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[8] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[8]),
        .Q(\rgf/rctl/rgf_c1bus_wb [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[9] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[9]),
        .Q(\rgf/rctl/rgf_c1bus_wb [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_rn_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(\rgf_selc0_rn_wb[0]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc0_rn_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_rn_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(ctl_selc0_rn),
        .Q(\rgf/rctl/rgf_selc0_rn_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_rn_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(\rgf_selc0_rn_wb[2]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc0_rn_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_stat_reg 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(\rgf/rctl/p_2_in ),
        .Q(\rgf/rctl/rgf_selc0_stat ),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(\rgf_selc0_wb[0]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc0_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(ctl_selc0),
        .Q(\rgf/rctl/rgf_selc0_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_rn_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(ctl_selc1_rn[0]),
        .Q(\rgf/rctl/rgf_selc1_rn_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_rn_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(\rgf_selc1_rn_wb[1]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc1_rn_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_rn_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(ctl_selc1_rn[2]),
        .Q(\rgf/rctl/rgf_selc1_rn_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_stat_reg 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(rgf_selc1_stat_i_2_n_0),
        .Q(\rgf/rctl/rgf_selc1_stat ),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(\rgf_selc1_wb[0]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc1_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(ctl_selc1),
        .Q(\rgf/rctl/rgf_selc1_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[0]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [0]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[10]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [10]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[11]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [11]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[12]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [12]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[13]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [13]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[14]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [14]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[15]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [15]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[1]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [1]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[2]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [2]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[3]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [3]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[4]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [4]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[5]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [5]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[6]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [6]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[7]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [7]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[8]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [8]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[9]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [9]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [0]),
        .Q(\rgf/sreg/sr [0]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [10]),
        .Q(\rgf/sreg/sr [10]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [11]),
        .Q(\rgf/sreg/sr [11]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [12]),
        .Q(\rgf/sreg/sr [12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [13]),
        .Q(\rgf/sreg/sr [13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [14]),
        .Q(\rgf/sreg/sr [14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [15]),
        .Q(\rgf/sreg/sr [15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [1]),
        .Q(\rgf/sreg/sr [1]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [2]),
        .Q(\rgf/sreg/sr [2]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [3]),
        .Q(\rgf/sreg/sr [3]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [4]),
        .Q(\rgf/sreg/sr [4]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [5]),
        .Q(\rgf/sreg/sr [5]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [6]),
        .Q(\rgf/sreg/sr [6]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [7]),
        .Q(\rgf/sreg/sr [7]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [8]),
        .Q(\rgf/sreg/sr [8]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in [9]),
        .Q(\rgf/sreg/sr [9]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [0]),
        .Q(\rgf/treg/tr [0]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [10]),
        .Q(\rgf/treg/tr [10]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [11]),
        .Q(\rgf/treg/tr [11]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [12]),
        .Q(\rgf/treg/tr [12]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [13]),
        .Q(\rgf/treg/tr [13]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [14]),
        .Q(\rgf/treg/tr [14]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [15]),
        .Q(\rgf/treg/tr [15]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [1]),
        .Q(\rgf/treg/tr [1]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [2]),
        .Q(\rgf/treg/tr [2]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [3]),
        .Q(\rgf/treg/tr [3]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [4]),
        .Q(\rgf/treg/tr [4]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [5]),
        .Q(\rgf/treg/tr [5]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [6]),
        .Q(\rgf/treg/tr [6]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [7]),
        .Q(\rgf/treg/tr [7]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [8]),
        .Q(\rgf/treg/tr [8]),
        .R(\rgf/treg/p_0_in ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [9]),
        .Q(\rgf/treg/tr [9]),
        .R(\rgf/treg/p_0_in ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[0]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry_n_7 ),
        .I2(\rgf_c0bus_wb[0]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[0]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_4_n_0 ),
        .O(c0bus[0]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[0]_i_10 
       (.I0(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h0800FFFF)) 
    \rgf_c0bus_wb[0]_i_11 
       (.I0(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000CA00FF00CA)) 
    \rgf_c0bus_wb[0]_i_12 
       (.I0(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hCECE333F020E020E)) 
    \rgf_c0bus_wb[0]_i_13 
       (.I0(a0bus_0[8]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[0]),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00F7F7F7)) 
    \rgf_c0bus_wb[0]_i_14 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(a0bus_0[15]),
        .I2(tout__1_carry_i_11_n_0),
        .I3(\rgf/sreg/sr [6]),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[0]_i_15 
       (.I0(a0bus_0[0]),
        .I1(a0bus_0[1]),
        .I2(a0bus_0[2]),
        .I3(a0bus_0[3]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000FFF0F55335533)) 
    \rgf_c0bus_wb[0]_i_16 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \rgf_c0bus_wb[0]_i_17 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[0]_i_2 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[0]),
        .I2(bdatr[0]),
        .I3(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E000E0)) 
    \rgf_c0bus_wb[0]_i_4 
       (.I0(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[0]_i_5 
       (.I0(bdatr[0]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[8]),
        .O(\rgf_c0bus_wb[0]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h82A22000)) 
    \rgf_c0bus_wb[0]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[0]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF2A20)) 
    \rgf_c0bus_wb[0]_i_7 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(a0bus_0[0]),
        .I4(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \rgf_c0bus_wb[0]_i_8 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF350035)) 
    \rgf_c0bus_wb[0]_i_9 
       (.I0(\rgf_c0bus_wb[4]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[10]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__1_n_5 ),
        .I2(\rgf_c0bus_wb[10]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[10]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .O(c0bus[10]));
  LUT6 #(
    .INIT(64'hFF47FFFFFF47FF00)) 
    \rgf_c0bus_wb[10]_i_10 
       (.I0(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[10]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[10]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h003AF03A0F3AFF3A)) 
    \rgf_c0bus_wb[10]_i_12 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[10]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[10]_i_14 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[10]_i_15 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hBFAA)) 
    \rgf_c0bus_wb[10]_i_16 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[9]),
        .I3(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hC0CFA0A0C0CFAFAF)) 
    \rgf_c0bus_wb[10]_i_17 
       (.I0(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[10]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[10]_i_19 
       (.I0(a0bus_0[8]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[10]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[10]_i_2 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .I3(bdatr[10]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(cbus_i[10]),
        .O(\rgf_c0bus_wb[10]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE1)) 
    \rgf_c0bus_wb[10]_i_20 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[10]_i_21 
       (.I0(a0bus_0[10]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[10]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c0bus_wb[10]_i_22 
       (.I0(a0bus_0[3]),
        .I1(a0bus_0[4]),
        .I2(a0bus_0[5]),
        .I3(a0bus_0[6]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[10]_i_23 
       (.I0(a0bus_0[12]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[10]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c0bus_wb[10]_i_4 
       (.I0(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_10_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[10]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[10]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[10]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c0bus_wb[10]_i_6 
       (.I0(a0bus_0[2]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEECCCCCFEEFFCCCF)) 
    \rgf_c0bus_wb[10]_i_7 
       (.I0(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[10]_i_8 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h00A3)) 
    \rgf_c0bus_wb[10]_i_9 
       (.I0(\rgf_c0bus_wb[10]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[11]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__1_n_4 ),
        .I2(\rgf_c0bus_wb[11]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_4_n_0 ),
        .O(c0bus[11]));
  LUT6 #(
    .INIT(64'hF7550000FFFFFFFF)) 
    \rgf_c0bus_wb[11]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA03F300F0)) 
    \rgf_c0bus_wb[11]_i_11 
       (.I0(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[11]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h55550F0F333300FF)) 
    \rgf_c0bus_wb[11]_i_13 
       (.I0(a0bus_0[11]),
        .I1(a0bus_0[12]),
        .I2(a0bus_0[13]),
        .I3(a0bus_0[14]),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5FFF0F3F3FFF0)) 
    \rgf_c0bus_wb[11]_i_14 
       (.I0(a0bus_0[11]),
        .I1(a0bus_0[12]),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[11]_i_15 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[11]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I1(a0bus_0[15]),
        .O(\rgf_c0bus_wb[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[11]_i_17 
       (.I0(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c0bus_wb[11]_i_18 
       (.I0(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[11]_i_2 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .I3(bdatr[11]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(cbus_i[11]),
        .O(\rgf_c0bus_wb[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFE00000)) 
    \rgf_c0bus_wb[11]_i_3 
       (.I0(a0bus_0[3]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00FF000E0000000E)) 
    \rgf_c0bus_wb[11]_i_4 
       (.I0(\rgf_c0bus_wb[11]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_10_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[11]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[11]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[11]_i_6 
       (.I0(a0bus_0[11]),
        .I1(\bdatw[11]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \rgf_c0bus_wb[11]_i_7 
       (.I0(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0A2A)) 
    \rgf_c0bus_wb[11]_i_8 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[11]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[10]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEEEFEEEEEE)) 
    \rgf_c0bus_wb[12]_i_1 
       (.I0(\rgf_c0bus_wb[12]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .O(c0bus[12]));
  LUT3 #(
    .INIT(8'hE0)) 
    \rgf_c0bus_wb[12]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c0bus_wb[12]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_12 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[12]_i_13 
       (.I0(\rgf_c0bus_wb[12]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_14 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[12]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_16 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_c0bus_wb[12]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_29_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02AA)) 
    \rgf_c0bus_wb[12]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c0bus_wb[12]_i_19 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF444F444FFFFF444)) 
    \rgf_c0bus_wb[12]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__2_n_7 ),
        .I2(cbus_i[12]),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(bdatr[12]),
        .I5(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hA8FF)) 
    \rgf_c0bus_wb[12]_i_20 
       (.I0(\rgf_c0bus_wb[12]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5FFF0F3F3FFF0)) 
    \rgf_c0bus_wb[12]_i_21 
       (.I0(a0bus_0[12]),
        .I1(a0bus_0[13]),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h4555BAAA)) 
    \rgf_c0bus_wb[12]_i_22 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[12]_i_23 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[12]_i_24 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[12]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF033F055)) 
    \rgf_c0bus_wb[12]_i_25 
       (.I0(a0bus_0[3]),
        .I1(a0bus_0[4]),
        .I2(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF00B8B8B8B8)) 
    \rgf_c0bus_wb[12]_i_26 
       (.I0(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h00FF3535)) 
    \rgf_c0bus_wb[12]_i_27 
       (.I0(a0bus_0[5]),
        .I1(a0bus_0[6]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c0bus_wb[12]_i_28 
       (.I0(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAABFFFFFFFF)) 
    \rgf_c0bus_wb[12]_i_29 
       (.I0(tout__1_carry_i_11_n_0),
        .I1(\badr[15]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/p_1_in [15]),
        .I3(\rgf/bank02/p_0_in [15]),
        .I4(\rgf/a0bus_out/rgf_c0bus_wb[12]_i_35_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFE0FFFFFFE00000)) 
    \rgf_c0bus_wb[12]_i_3 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hF077F000)) 
    \rgf_c0bus_wb[12]_i_30 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_36_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAEAAAAA)) 
    \rgf_c0bus_wb[12]_i_31 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[12]_i_32 
       (.I0(a0bus_0[7]),
        .I1(a0bus_0[8]),
        .I2(a0bus_0[9]),
        .I3(a0bus_0[10]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h55550F0F333300FF)) 
    \rgf_c0bus_wb[12]_i_33 
       (.I0(a0bus_0[3]),
        .I1(a0bus_0[4]),
        .I2(a0bus_0[5]),
        .I3(a0bus_0[6]),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c0bus_wb[12]_i_34 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[12]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[12]_i_36 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[0]),
        .O(\rgf_c0bus_wb[12]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c0bus_wb[12]_i_39 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(ctl_sela0_rn[0]),
        .I3(\badr[15]_INST_0_i_28_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr01 [15]),
        .O(\rgf_c0bus_wb[12]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0E0E0E0E02020E00)) 
    \rgf_c0bus_wb[12]_i_4 
       (.I0(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c0bus_wb[12]_i_40 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[2]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[0]),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr02 [15]),
        .O(\rgf_c0bus_wb[12]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c0bus_wb[12]_i_41 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(\badr[15]_INST_0_i_28_n_0 ),
        .I2(ctl_sela0_rn[0]),
        .I3(ctl_sela0_rn[2]),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr05 [15]),
        .O(\rgf_c0bus_wb[12]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c0bus_wb[12]_i_42 
       (.I0(\badr[15]_INST_0_i_191_n_0 ),
        .I1(ctl_sela0_rn[0]),
        .I2(\badr[15]_INST_0_i_28_n_0 ),
        .I3(ctl_sela0_rn[2]),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr06 [15]),
        .O(\rgf_c0bus_wb[12]_i_42_n_0 ));
  LUT4 #(
    .INIT(16'h0E04)) 
    \rgf_c0bus_wb[12]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8F8F8F008F8F8F8F)) 
    \rgf_c0bus_wb[12]_i_6 
       (.I0(a0bus_0[11]),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[12]_i_7 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\rgf_c0bus_wb[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF028AFF8A028A02)) 
    \rgf_c0bus_wb[12]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[12]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[12]_i_9 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[12]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[12]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[13]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__2_n_6 ),
        .I2(\rgf_c0bus_wb[13]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .O(c0bus[13]));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[13]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[13]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F5F305F)) 
    \rgf_c0bus_wb[13]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \rgf_c0bus_wb[13]_i_12 
       (.I0(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF000F0FF33553355)) 
    \rgf_c0bus_wb[13]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h01510000FFFFFFFF)) 
    \rgf_c0bus_wb[13]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h2227772700000000)) 
    \rgf_c0bus_wb[13]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_16 
       (.I0(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[13]_i_17 
       (.I0(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[13]_i_18 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[13]_i_19 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[13]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[13]_i_2 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .I3(bdatr[13]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(cbus_i[13]),
        .O(\rgf_c0bus_wb[13]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_20 
       (.I0(a0bus_0[13]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[14]),
        .O(\rgf_c0bus_wb[13]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[13]_i_21 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_22 
       (.I0(a0bus_0[2]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[13]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_23 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[13]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_24 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[13]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_25 
       (.I0(a0bus_0[10]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[13]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_26 
       (.I0(a0bus_0[8]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[13]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_27 
       (.I0(a0bus_0[6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[13]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[13]_i_28 
       (.I0(a0bus_0[4]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[13]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hABFEAB32A8CEA802)) 
    \rgf_c0bus_wb[13]_i_29 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[13]),
        .I5(a0bus_0[14]),
        .O(\rgf_c0bus_wb[13]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFE00000)) 
    \rgf_c0bus_wb[13]_i_3 
       (.I0(a0bus_0[5]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hE000E0E0E000E000)) 
    \rgf_c0bus_wb[13]_i_4 
       (.I0(\rgf_c0bus_wb[13]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb_reg[13]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[13]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[13]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[13]_i_6 
       (.I0(a0bus_0[13]),
        .I1(\bdatw[13]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000033330000550F)) 
    \rgf_c0bus_wb[13]_i_7 
       (.I0(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h3323332003230320)) 
    \rgf_c0bus_wb[13]_i_9 
       (.I0(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[14]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__2_n_5 ),
        .I2(\rgf_c0bus_wb[14]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .O(c0bus[14]));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[14]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[14]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[14]_i_11 
       (.I0(tout__1_carry_i_11_n_0),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000AACCAACC)) 
    \rgf_c0bus_wb[14]_i_13 
       (.I0(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA5595)) 
    \rgf_c0bus_wb[14]_i_14 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[14]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c0bus_wb[14]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rgf_c0bus_wb[14]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(a0bus_0[15]),
        .O(\rgf_c0bus_wb[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[14]_i_18 
       (.I0(\rgf_c0bus_wb[14]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8F0F0F0)) 
    \rgf_c0bus_wb[14]_i_19 
       (.I0(a0bus_0[14]),
        .I1(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[14]_i_2 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .I3(bdatr[14]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(cbus_i[14]),
        .O(\rgf_c0bus_wb[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_20 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[14]_i_21 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_22 
       (.I0(a0bus_0[1]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[14]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_23 
       (.I0(a0bus_0[4]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[14]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_24 
       (.I0(a0bus_0[6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[14]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[14]_i_25 
       (.I0(a0bus_0[12]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[14]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[14]_i_26 
       (.I0(a0bus_0[14]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .O(\rgf_c0bus_wb[14]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_27 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[14]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_28 
       (.I0(a0bus_0[14]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[14]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_29 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFE0FFFFFFE00000)) 
    \rgf_c0bus_wb[14]_i_3 
       (.I0(a0bus_0[6]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_30 
       (.I0(a0bus_0[1]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[14]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[14]_i_31 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[14]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_32 
       (.I0(a0bus_0[11]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[14]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_33 
       (.I0(a0bus_0[9]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[14]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_34 
       (.I0(a0bus_0[7]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[14]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[14]_i_35 
       (.I0(a0bus_0[5]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[14]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hE000E0E0E000E000)) 
    \rgf_c0bus_wb[14]_i_4 
       (.I0(\rgf_c0bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[14]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[14]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[14]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[14]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[14]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF0501111F050FF11)) 
    \rgf_c0bus_wb[14]_i_7 
       (.I0(\rgf_c0bus_wb[14]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hC0CF50500F0F0F0F)) 
    \rgf_c0bus_wb[14]_i_8 
       (.I0(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0545554505405540)) 
    \rgf_c0bus_wb[14]_i_9 
       (.I0(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[15]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/p_0_in ),
        .I2(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_5_n_0 ),
        .O(c0bus[15]));
  LUT6 #(
    .INIT(64'hFF10B0FFB010B010)) 
    \rgf_c0bus_wb[15]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h82880808)) 
    \rgf_c0bus_wb[15]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[15]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[15]_i_12 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(a0bus_0[14]),
        .I2(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[15]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c0bus_wb[15]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h8AFF)) 
    \rgf_c0bus_wb[15]_i_15 
       (.I0(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF003A003A00)) 
    \rgf_c0bus_wb[15]_i_16 
       (.I0(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I5(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c0bus_wb[15]_i_17 
       (.I0(\ctl0/stat [1]),
        .I1(\ctl0/stat [0]),
        .I2(\fch/ir0 [15]),
        .O(\rgf_c0bus_wb[15]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4500)) 
    \rgf_c0bus_wb[15]_i_18 
       (.I0(\ccmd[0]_INST_0_i_8_n_0 ),
        .I1(\ccmd[0]_INST_0_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_36_n_0 ),
        .I3(\ccmd[0]_INST_0_i_3_n_0 ),
        .I4(\ccmd[0]_INST_0_i_5_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055550001)) 
    \rgf_c0bus_wb[15]_i_19 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [11]),
        .I3(\ctl0/stat [1]),
        .I4(\fch/ir0 [12]),
        .I5(\ccmd[0]_INST_0_i_14_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c0bus_wb[15]_i_2 
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAEA000000000000)) 
    \rgf_c0bus_wb[15]_i_20 
       (.I0(\rgf_c0bus_wb[15]_i_37_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\ccmd[0]_INST_0_i_19_n_0 ),
        .I4(\ccmd[0]_INST_0_i_6_n_0 ),
        .I5(\ccmd[0]_INST_0_i_5_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[15]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .I2(tout__1_carry_i_11_n_0),
        .O(\rgf_c0bus_wb[15]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[15]_i_22 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[15]_i_23 
       (.I0(a0bus_0[2]),
        .I1(a0bus_0[3]),
        .I2(a0bus_0[4]),
        .I3(a0bus_0[5]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h45BA)) 
    \rgf_c0bus_wb[15]_i_24 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h550F3300550F33FF)) 
    \rgf_c0bus_wb[15]_i_25 
       (.I0(a0bus_0[0]),
        .I1(a0bus_0[1]),
        .I2(a0bus_0[15]),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[15]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[15]_i_26 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \rgf_c0bus_wb[15]_i_27 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[15]_i_28 
       (.I0(a0bus_0[6]),
        .I1(a0bus_0[7]),
        .I2(a0bus_0[8]),
        .I3(a0bus_0[9]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[15]_i_29 
       (.I0(a0bus_0[10]),
        .I1(a0bus_0[11]),
        .I2(a0bus_0[12]),
        .I3(a0bus_0[13]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFE0FFFFFFE00000)) 
    \rgf_c0bus_wb[15]_i_3 
       (.I0(a0bus_0[7]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_30 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c0bus_wb[15]_i_31 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h3A)) 
    \rgf_c0bus_wb[15]_i_32 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_33 
       (.I0(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hAA59)) 
    \rgf_c0bus_wb[15]_i_34 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[15]_i_35 
       (.I0(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \rgf_c0bus_wb[15]_i_36 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [11]),
        .I3(\ccmd[0]_INST_0_i_11_n_0 ),
        .I4(\fch/ir0 [12]),
        .I5(\fch/ir0 [14]),
        .O(\rgf_c0bus_wb[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_c0bus_wb[15]_i_37 
       (.I0(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\bdatw[15]_INST_0_i_20_n_0 ),
        .I4(\fadr[15]_INST_0_i_11_n_0 ),
        .I5(\ccmd[2]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[15]_i_38 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[15]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_39 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[15]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF8A)) 
    \rgf_c0bus_wb[15]_i_4 
       (.I0(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_40 
       (.I0(a0bus_0[5]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[15]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_41 
       (.I0(a0bus_0[11]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[15]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_42 
       (.I0(a0bus_0[13]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[15]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[15]_i_43 
       (.I0(a0bus_0[14]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[15]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h88888F8888888888)) 
    \rgf_c0bus_wb[15]_i_5 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[15]),
        .I2(\mem/read_cyc [3]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(bdatr[15]),
        .O(\rgf_c0bus_wb[15]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c0bus_wb[15]_i_6 
       (.I0(\ctl0/stat [2]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011111151)) 
    \rgf_c0bus_wb[15]_i_7 
       (.I0(\ccmd[2]_INST_0_i_3_n_0 ),
        .I1(\ctl0/stat [2]),
        .I2(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I3(\fadr[15]_INST_0_i_14_n_0 ),
        .I4(\fadr[15]_INST_0_i_15_n_0 ),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF51)) 
    \rgf_c0bus_wb[15]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_18_n_0 ),
        .I1(\ccmd[0]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I4(\ctl0/stat [2]),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h15)) 
    \rgf_c0bus_wb[15]_i_9 
       (.I0(tout__1_carry_i_10_n_0),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\bbus_o[7]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[1]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry_n_6 ),
        .I2(\rgf_c0bus_wb[1]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_4_n_0 ),
        .O(c0bus[1]));
  LUT6 #(
    .INIT(64'hDDD0DDD0DDDDDDD0)) 
    \rgf_c0bus_wb[1]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[1]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hC0CCC00088CC88CC)) 
    \rgf_c0bus_wb[1]_i_12 
       (.I0(\rgf_c0bus_wb[1]_i_16_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \rgf_c0bus_wb[1]_i_13 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000444EEE4E)) 
    \rgf_c0bus_wb[1]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[1]_i_15 
       (.I0(a0bus_0[1]),
        .I1(a0bus_0[2]),
        .I2(a0bus_0[3]),
        .I3(a0bus_0[4]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFFAACCAACC)) 
    \rgf_c0bus_wb[1]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hF000F0FF33553355)) 
    \rgf_c0bus_wb[1]_i_17 
       (.I0(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c0bus_wb[1]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h740374CF773377FF)) 
    \rgf_c0bus_wb[1]_i_19 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[13]),
        .I5(a0bus_0[14]),
        .O(\rgf_c0bus_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF22F222F222F2)) 
    \rgf_c0bus_wb[1]_i_2 
       (.I0(bdatr[1]),
        .I1(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(cbus_i[1]),
        .O(\rgf_c0bus_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBAAA4555FFFFFFFF)) 
    \rgf_c0bus_wb[1]_i_20 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[1]_i_3 
       (.I0(\rgf_c0bus_wb[1]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A0000)) 
    \rgf_c0bus_wb[1]_i_4 
       (.I0(\rgf_c0bus_wb[1]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_11_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[1]_i_5 
       (.I0(bdatr[1]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[9]),
        .O(\rgf_c0bus_wb[1]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h57F7)) 
    \rgf_c0bus_wb[1]_i_6 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC300EFEEC300E322)) 
    \rgf_c0bus_wb[1]_i_7 
       (.I0(a0bus_0[9]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(a0bus_0[1]),
        .I3(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I4(tout__1_carry_i_10_n_0),
        .I5(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h6080E000)) 
    \rgf_c0bus_wb[1]_i_8 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[1]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[0]),
        .O(\rgf_c0bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[2]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry_n_5 ),
        .I2(\rgf_c0bus_wb[2]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .O(c0bus[2]));
  LUT6 #(
    .INIT(64'hA8A8A8202020A820)) 
    \rgf_c0bus_wb[2]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[2]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hDC1CD010)) 
    \rgf_c0bus_wb[2]_i_12 
       (.I0(\rgf_c0bus_wb[10]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[2]_i_2 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[2]),
        .I2(\rgf_c0bus_wb[2]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(bdatr[2]),
        .I5(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[2]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFF00020000000200)) 
    \rgf_c0bus_wb[2]_i_4 
       (.I0(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[2]_i_5 
       (.I0(bdatr[2]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[10]),
        .O(\rgf_c0bus_wb[2]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF757)) 
    \rgf_c0bus_wb[2]_i_6 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(a0bus_0[2]),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCECE020E333F020E)) 
    \rgf_c0bus_wb[2]_i_7 
       (.I0(a0bus_0[10]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I5(a0bus_0[2]),
        .O(\rgf_c0bus_wb[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h8A222000)) 
    \rgf_c0bus_wb[2]_i_8 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(a0bus_0[2]),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCFEECFCCCFEECFFF)) 
    \rgf_c0bus_wb[2]_i_9 
       (.I0(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[3]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry_n_4 ),
        .I2(\rgf_c0bus_wb[3]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .O(c0bus[3]));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[3]_i_10 
       (.I0(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFF8A0000)) 
    \rgf_c0bus_wb[3]_i_11 
       (.I0(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFEEFFE2)) 
    \rgf_c0bus_wb[3]_i_12 
       (.I0(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0E0E0E00FFFFFFFF)) 
    \rgf_c0bus_wb[3]_i_13 
       (.I0(\rgf_c0bus_wb[3]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h303F303FA0A0AFAF)) 
    \rgf_c0bus_wb[3]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[3]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h40004404FFFFFFFF)) 
    \rgf_c0bus_wb[3]_i_16 
       (.I0(\rgf_c0bus_wb[3]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3FA0AFA0AF)) 
    \rgf_c0bus_wb[3]_i_17 
       (.I0(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBEEEEBEEE)) 
    \rgf_c0bus_wb[3]_i_18 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[3]_i_2 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[3]),
        .I2(\rgf_c0bus_wb[3]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(bdatr[3]),
        .I5(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[3]_i_3 
       (.I0(\rgf_c0bus_wb[3]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF888A)) 
    \rgf_c0bus_wb[3]_i_4 
       (.I0(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_12_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[3]_i_5 
       (.I0(bdatr[3]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[11]),
        .O(\rgf_c0bus_wb[3]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c0bus_wb[3]_i_6 
       (.I0(a0bus_0[3]),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCECE333F020E020E)) 
    \rgf_c0bus_wb[3]_i_7 
       (.I0(a0bus_0[11]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[3]),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[3]_i_8 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[3]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[3]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[4]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__0_n_7 ),
        .I2(\rgf_c0bus_wb[4]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .O(c0bus[4]));
  LUT5 #(
    .INIT(32'h474700FF)) 
    \rgf_c0bus_wb[4]_i_10 
       (.I0(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hBBBBBBAB)) 
    \rgf_c0bus_wb[4]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h88CCC0CC8800C0CC)) 
    \rgf_c0bus_wb[4]_i_12 
       (.I0(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00660F66)) 
    \rgf_c0bus_wb[4]_i_13 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[4]_i_14 
       (.I0(a0bus_0[4]),
        .I1(a0bus_0[5]),
        .I2(a0bus_0[6]),
        .I3(a0bus_0[7]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hAABAAAAA)) 
    \rgf_c0bus_wb[4]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[4]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \rgf_c0bus_wb[4]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[4]_i_17 
       (.I0(a0bus_0[12]),
        .I1(tout__1_carry_i_11_n_0),
        .O(\rgf_c0bus_wb[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[4]_i_2 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[4]),
        .I2(bdatr[4]),
        .I3(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD3200000)) 
    \rgf_c0bus_wb[4]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A0000)) 
    \rgf_c0bus_wb[4]_i_4 
       (.I0(\rgf_c0bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_11_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[4]_i_5 
       (.I0(bdatr[4]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[12]),
        .O(\rgf_c0bus_wb[4]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[4]_i_6 
       (.I0(\ccmd[1]_INST_0_i_1_n_0 ),
        .I1(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \rgf_c0bus_wb[4]_i_7 
       (.I0(\ctl0/stat [2]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0080C080CCCCCCCC)) 
    \rgf_c0bus_wb[4]_i_8 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[4]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[5]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__0_n_6 ),
        .I2(\rgf_c0bus_wb[5]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .O(c0bus[5]));
  LUT6 #(
    .INIT(64'h8888888A8888AA8A)) 
    \rgf_c0bus_wb[5]_i_10 
       (.I0(\rgf_c0bus_wb[5]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[5]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8800C0CC88CCC0CC)) 
    \rgf_c0bus_wb[5]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h01510000FFFFFFFF)) 
    \rgf_c0bus_wb[5]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[5]_i_14 
       (.I0(a0bus_0[5]),
        .I1(a0bus_0[6]),
        .I2(a0bus_0[7]),
        .I3(a0bus_0[8]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[5]_i_15 
       (.I0(a0bus_0[9]),
        .I1(a0bus_0[10]),
        .I2(a0bus_0[11]),
        .I3(a0bus_0[12]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[5]_i_2 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[5]),
        .I2(bdatr[5]),
        .I3(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[5]_i_3 
       (.I0(\rgf_c0bus_wb[5]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A0000)) 
    \rgf_c0bus_wb[5]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_11_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[5]_i_5 
       (.I0(bdatr[5]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[13]),
        .O(\rgf_c0bus_wb[5]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c0bus_wb[5]_i_6 
       (.I0(a0bus_0[5]),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC300E322C300EFEE)) 
    \rgf_c0bus_wb[5]_i_7 
       (.I0(a0bus_0[13]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(a0bus_0[5]),
        .I3(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I4(tout__1_carry_i_10_n_0),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[5]_i_8 
       (.I0(a0bus_0[5]),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[5]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[6]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__0_n_5 ),
        .I2(\rgf_c0bus_wb[6]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .O(c0bus[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFF55544454)) 
    \rgf_c0bus_wb[6]_i_10 
       (.I0(\rgf_c0bus_wb[6]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7444747474444444)) 
    \rgf_c0bus_wb[6]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[6]_i_12 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[6]_i_13 
       (.I0(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0100FFFF)) 
    \rgf_c0bus_wb[6]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[6]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[5]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hC5C0C5CF)) 
    \rgf_c0bus_wb[6]_i_16 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[6]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \rgf_c0bus_wb[6]_i_2 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[6]),
        .I2(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(bdatr[6]),
        .I5(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFD0)) 
    \rgf_c0bus_wb[6]_i_3 
       (.I0(\rgf_c0bus_wb[6]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0020F02000200020)) 
    \rgf_c0bus_wb[6]_i_4 
       (.I0(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[6]_i_5 
       (.I0(bdatr[6]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[14]),
        .O(\rgf_c0bus_wb[6]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hD1FF)) 
    \rgf_c0bus_wb[6]_i_6 
       (.I0(a0bus_0[6]),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hC300E322C300EFEE)) 
    \rgf_c0bus_wb[6]_i_7 
       (.I0(a0bus_0[14]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(a0bus_0[6]),
        .I3(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I4(tout__1_carry_i_10_n_0),
        .I5(\bbus_o[6]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c0bus_wb[6]_i_8 
       (.I0(a0bus_0[6]),
        .I1(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCFFFCDFDCCFCCDFD)) 
    \rgf_c0bus_wb[6]_i_9 
       (.I0(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF4FF)) 
    \rgf_c0bus_wb[7]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__0_n_4 ),
        .I2(\rgf_c0bus_wb[7]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_4_n_0 ),
        .O(c0bus[7]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_10 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hA20A0800)) 
    \rgf_c0bus_wb[7]_i_11 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\bbus_o[7]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[7]),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h7575757530303033)) 
    \rgf_c0bus_wb[7]_i_12 
       (.I0(\rgf_c0bus_wb[7]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c0bus_wb[7]_i_13 
       (.I0(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I1(a0bus_0[6]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hBFAE)) 
    \rgf_c0bus_wb[7]_i_14 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[7]_i_15 
       (.I0(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_16 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c0bus_wb[7]_i_17 
       (.I0(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h8AAA)) 
    \rgf_c0bus_wb[7]_i_18 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[7]_i_19 
       (.I0(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF22F222F222F2)) 
    \rgf_c0bus_wb[7]_i_2 
       (.I0(bdatr[7]),
        .I1(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(cbus_i[7]),
        .O(\rgf_c0bus_wb[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000000004544FFFF)) 
    \rgf_c0bus_wb[7]_i_3 
       (.I0(\rgf_c0bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00F0F0F020202020)) 
    \rgf_c0bus_wb[7]_i_4 
       (.I0(\rgf_c0bus_wb[7]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_15_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[7]_i_5 
       (.I0(bdatr[7]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[15]),
        .O(\rgf_c0bus_wb[7]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c0bus_wb[7]_i_6 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .O(\rgf_c0bus_wb[7]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h08C8)) 
    \rgf_c0bus_wb[7]_i_7 
       (.I0(a0bus_0[7]),
        .I1(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(\bbus_o[7]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hAABE)) 
    \rgf_c0bus_wb[7]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(a0bus_0[7]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_9 
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[8]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__1_n_7 ),
        .I2(\rgf_c0bus_wb[8]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[8]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .O(c0bus[8]));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c0bus_wb[8]_i_10 
       (.I0(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hBFAA)) 
    \rgf_c0bus_wb[8]_i_11 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[7]),
        .I3(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A8AFF8A8A8A00)) 
    \rgf_c0bus_wb[8]_i_12 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[8]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[8]_i_13 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h3F3F505F3030505F)) 
    \rgf_c0bus_wb[8]_i_14 
       (.I0(\rgf_c0bus_wb[15]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_43_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h55550F0F333300FF)) 
    \rgf_c0bus_wb[8]_i_15 
       (.I0(a0bus_0[12]),
        .I1(a0bus_0[13]),
        .I2(a0bus_0[14]),
        .I3(a0bus_0[15]),
        .I4(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c0bus_wb[8]_i_16 
       (.I0(a0bus_0[8]),
        .I1(a0bus_0[9]),
        .I2(a0bus_0[10]),
        .I3(a0bus_0[11]),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF040004000400)) 
    \rgf_c0bus_wb[8]_i_2 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .I3(bdatr[8]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(cbus_i[8]),
        .O(\rgf_c0bus_wb[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h08080808AA08AAAA)) 
    \rgf_c0bus_wb[8]_i_4 
       (.I0(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[8]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[8]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[8]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c0bus_wb[8]_i_6 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h08F8FFFF)) 
    \rgf_c0bus_wb[8]_i_7 
       (.I0(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hCA00FFFF)) 
    \rgf_c0bus_wb[8]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0511FFFF05110511)) 
    \rgf_c0bus_wb[8]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFF4)) 
    \rgf_c0bus_wb[9]_i_1 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__1_n_6 ),
        .I2(\rgf_c0bus_wb[9]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb_reg[9]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .O(c0bus[9]));
  LUT6 #(
    .INIT(64'h5510051050100010)) 
    \rgf_c0bus_wb[9]_i_10 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFA8A8FFA8A8A800)) 
    \rgf_c0bus_wb[9]_i_11 
       (.I0(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I3(a0bus_0[9]),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h4747FF00)) 
    \rgf_c0bus_wb[9]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF55335533)) 
    \rgf_c0bus_wb[9]_i_13 
       (.I0(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[9]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[9]_i_15 
       (.I0(\rgf_c0bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_16 
       (.I0(a0bus_0[7]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[9]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_17 
       (.I0(a0bus_0[9]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[9]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h56)) 
    \rgf_c0bus_wb[9]_i_18 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c0bus_wb[9]_i_19 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88888F8888888888)) 
    \rgf_c0bus_wb[9]_i_2 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(cbus_i[9]),
        .I2(\mem/read_cyc [3]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(bdatr[9]),
        .O(\rgf_c0bus_wb[9]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[9]_i_20 
       (.I0(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c0bus_wb[9]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_22 
       (.I0(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF0F02020F0002020)) 
    \rgf_c0bus_wb[9]_i_4 
       (.I0(\rgf_c0bus_wb[9]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c0bus_wb[9]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[9]),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I4(\bdatw[9]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c0bus_wb[9]_i_6 
       (.I0(a0bus_0[1]),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEECCCCFCEEFFCCFC)) 
    \rgf_c0bus_wb[9]_i_7 
       (.I0(\rgf_c0bus_wb[9]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF70FF70707070)) 
    \rgf_c0bus_wb[9]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I1(a0bus_0[8]),
        .I2(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000CA00FF00CA00)) 
    \rgf_c0bus_wb[9]_i_9 
       (.I0(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[0]_i_3 
       (.I0(\rgf_c0bus_wb[0]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .O(\rgf_c0bus_wb_reg[0]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[10]_i_3 
       (.I0(\rgf_c0bus_wb[10]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_6_n_0 ),
        .O(\rgf_c0bus_wb_reg[10]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[13]_i_8 
       (.I0(\rgf_c0bus_wb[13]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_15_n_0 ),
        .O(\rgf_c0bus_wb_reg[13]_i_8_n_0 ),
        .S(\bbus_o[4]_INST_0_i_1_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[8]_i_3 
       (.I0(\rgf_c0bus_wb[8]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_6_n_0 ),
        .O(\rgf_c0bus_wb_reg[8]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[9]_i_3 
       (.I0(\rgf_c0bus_wb[9]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_6_n_0 ),
        .O(\rgf_c0bus_wb_reg[9]_i_3_n_0 ),
        .S(\rgf_c0bus_wb[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEFEE)) 
    \rgf_c1bus_wb[0]_i_1 
       (.I0(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I3(\alu1/art/add/tout__1_carry_n_7 ),
        .I4(\rgf_c1bus_wb_reg[0]_i_4_n_0 ),
        .O(c1bus[0]));
  LUT6 #(
    .INIT(64'hF000B0F000008000)) 
    \rgf_c1bus_wb[0]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(a1bus_0[0]),
        .I4(\bdatw[8]_INST_0_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000454500FFC3C3)) 
    \rgf_c1bus_wb[0]_i_11 
       (.I0(\rgf_c1bus_wb[0]_i_16_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h007F7F7F)) 
    \rgf_c1bus_wb[0]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[10]_i_24_n_0 ),
        .I3(\rgf/sreg/sr [6]),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \rgf_c1bus_wb[0]_i_13 
       (.I0(\bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_c1bus_wb[0]_i_14 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[9]_INST_0_i_13_n_0 ),
        .I4(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000200000000000)) 
    \rgf_c1bus_wb[0]_i_15 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[0]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[0]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AEAE00AE)) 
    \rgf_c1bus_wb[0]_i_2 
       (.I0(\rgf_c1bus_wb[0]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[0]_i_3 
       (.I0(\mem/read_cyc [1]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [3]),
        .I3(bdatr[0]),
        .I4(\mem/read_cyc [0]),
        .I5(bdatr[8]),
        .O(\rgf_c1bus_wb[0]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \rgf_c1bus_wb[0]_i_5 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h57DF)) 
    \rgf_c1bus_wb[0]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hDCDCDDCC)) 
    \rgf_c1bus_wb[0]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFF77F77)) 
    \rgf_c1bus_wb[0]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDDDFFF)) 
    \rgf_c1bus_wb[0]_i_9 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF10111010)) 
    \rgf_c1bus_wb[10]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_6_n_0 ),
        .O(c1bus[10]));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[10]_i_10 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[4]),
        .I2(a1bus_0[5]),
        .I3(a1bus_0[6]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hCCC4CCC4CCC444C4)) 
    \rgf_c1bus_wb[10]_i_11 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \rgf_c1bus_wb[10]_i_12 
       (.I0(\bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF077F044)) 
    \rgf_c1bus_wb[10]_i_13 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hBAAA)) 
    \rgf_c1bus_wb[10]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(a1bus_0[15]),
        .O(\rgf_c1bus_wb[10]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[10]_i_15 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[10]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFF54FF54FFFFFF54)) 
    \rgf_c1bus_wb[10]_i_17 
       (.I0(\rgf_c1bus_wb[10]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[10]_i_18 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(a1bus_0[14]),
        .I3(a1bus_0[15]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h000800000008000F)) 
    \rgf_c1bus_wb[10]_i_19 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h1BFB)) 
    \rgf_c1bus_wb[10]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAA800000000)) 
    \rgf_c1bus_wb[10]_i_20 
       (.I0(\rgf_c1bus_wb[10]_i_24_n_0 ),
        .I1(\badr[15]_INST_0_i_9_n_0 ),
        .I2(\rgf/bank02/p_1_in1_in [15]),
        .I3(\rgf/bank02/p_0_in0_in [15]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[10]_i_25_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[10]_i_21 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[10]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[10]_i_22 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c1bus_wb[10]_i_23 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(a1bus_0[10]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\bdatw[10]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[10]_i_24 
       (.I0(\ctl1/stat [2]),
        .I1(\rgf_c1bus_wb[15]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c1bus_wb[10]_i_28 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_52_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr01 [15]),
        .O(\rgf_c1bus_wb[10]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \rgf_c1bus_wb[10]_i_29 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_40_n_0 ),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(ctl_sela1_rn),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr02 [15]),
        .O(\rgf_c1bus_wb[10]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hC8C8C8080808C808)) 
    \rgf_c1bus_wb[10]_i_3 
       (.I0(\rgf_c1bus_wb[10]_i_7_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_30 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(\badr[15]_INST_0_i_52_n_0 ),
        .I2(ctl_sela1_rn),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr05 [15]),
        .O(\rgf_c1bus_wb[10]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_31 
       (.I0(\badr[15]_INST_0_i_235_n_0 ),
        .I1(ctl_sela1_rn),
        .I2(\badr[15]_INST_0_i_52_n_0 ),
        .I3(\badr[15]_INST_0_i_40_n_0 ),
        .I4(\bdatw[15]_INST_0_i_238_n_0 ),
        .I5(\rgf/bank13/gr06 [15]),
        .O(\rgf_c1bus_wb[10]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hBFAA)) 
    \rgf_c1bus_wb[10]_i_4 
       (.I0(\rgf_c1bus_wb[10]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(a1bus_0[9]),
        .I3(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFF2FFF0FFF2FFFA)) 
    \rgf_c1bus_wb[10]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[10]_i_6 
       (.I0(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I1(bdatr[10]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(\alu1/art/add/tout__1_carry__1_n_5 ),
        .I4(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h0000ACFF)) 
    \rgf_c1bus_wb[10]_i_7 
       (.I0(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[10]_i_8 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[8]),
        .I2(a1bus_0[9]),
        .I3(a1bus_0[10]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h6566)) 
    \rgf_c1bus_wb[10]_i_9 
       (.I0(\bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\bdatw[9]_INST_0_i_13_n_0 ),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    \rgf_c1bus_wb[11]_i_1 
       (.I0(\rgf_c1bus_wb[11]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I2(\alu1/art/add/tout__1_carry__1_n_4 ),
        .I3(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I4(bdatr[11]),
        .I5(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .O(c1bus[11]));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[11]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[11]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[11]_i_11 
       (.I0(a1bus_0[11]),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[11]_i_12 
       (.I0(\rgf_c1bus_wb[13]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h000000E2)) 
    \rgf_c1bus_wb[11]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0F5F5FFF0F3F3)) 
    \rgf_c1bus_wb[11]_i_14 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[11]_i_15 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(a1bus_0[13]),
        .I3(a1bus_0[14]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[11]_i_16 
       (.I0(\bdatw[9]_INST_0_i_13_n_0 ),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[11]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_61_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_62_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_63_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_64_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[11]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[11]_i_19 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(a1bus_0[2]),
        .I3(a1bus_0[3]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220002)) 
    \rgf_c1bus_wb[11]_i_2 
       (.I0(\rgf_c1bus_wb[11]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_6_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAFEFFFFAAFE)) 
    \rgf_c1bus_wb[11]_i_3 
       (.I0(\rgf_c1bus_wb[11]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[11]_i_4 
       (.I0(a1bus_0[10]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h2220AAA822202220)) 
    \rgf_c1bus_wb[11]_i_5 
       (.I0(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A808A8AAAAAAAAA)) 
    \rgf_c1bus_wb[11]_i_6 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I4(a1bus_0[15]),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h20202023AFAFAFAF)) 
    \rgf_c1bus_wb[11]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[11]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[11]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\bdatw[11]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[11]_i_9 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F44)) 
    \rgf_c1bus_wb[12]_i_1 
       (.I0(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I1(\alu1/art/add/tout__1_carry__2_n_7 ),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(bdatr[12]),
        .I4(\rgf_c1bus_wb[12]_i_2_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .O(c1bus[12]));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c1bus_wb[12]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00470047000000FF)) 
    \rgf_c1bus_wb[12]_i_11 
       (.I0(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[12]_i_12 
       (.I0(a1bus_0[11]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h20333333)) 
    \rgf_c1bus_wb[12]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(a1bus_0[15]),
        .O(\rgf_c1bus_wb[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0002220200000000)) 
    \rgf_c1bus_wb[12]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h000002A2)) 
    \rgf_c1bus_wb[12]_i_15 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[12]_i_16 
       (.I0(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \rgf_c1bus_wb[12]_i_17 
       (.I0(a1bus_0[14]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [6]),
        .I4(a1bus_0[0]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[12]_i_18 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(a1bus_0[14]),
        .I3(a1bus_0[15]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[12]_i_19 
       (.I0(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFAAFE)) 
    \rgf_c1bus_wb[12]_i_2 
       (.I0(\rgf_c1bus_wb[12]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hE2FFE200E2FFE2FF)) 
    \rgf_c1bus_wb[12]_i_20 
       (.I0(\rgf_c1bus_wb[12]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[12]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[12]_i_21 
       (.I0(a1bus_0[0]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_22 
       (.I0(a1bus_0[1]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .O(\rgf_c1bus_wb[12]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_23 
       (.I0(a1bus_0[12]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[13]),
        .O(\rgf_c1bus_wb[12]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_24 
       (.I0(a1bus_0[5]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[6]),
        .O(\rgf_c1bus_wb[12]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_25 
       (.I0(a1bus_0[3]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[4]),
        .O(\rgf_c1bus_wb[12]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_26 
       (.I0(a1bus_0[7]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[8]),
        .O(\rgf_c1bus_wb[12]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_27 
       (.I0(a1bus_0[9]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[10]),
        .O(\rgf_c1bus_wb[12]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_28 
       (.I0(a1bus_0[4]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[3]),
        .O(\rgf_c1bus_wb[12]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAFAC8CA)) 
    \rgf_c1bus_wb[12]_i_3 
       (.I0(\rgf_c1bus_wb[12]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_9_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h80802888)) 
    \rgf_c1bus_wb[12]_i_4 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\bdatw[12]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[12]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(a1bus_0[4]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[12]_i_6 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hD0D0D000)) 
    \rgf_c1bus_wb[12]_i_7 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I3(a1bus_0[12]),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAA2AAAAAAA2AAA2)) 
    \rgf_c1bus_wb[12]_i_8 
       (.I0(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[12]_i_9 
       (.I0(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBAFFBABA)) 
    \rgf_c1bus_wb[13]_i_1 
       (.I0(\rgf_c1bus_wb[13]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I2(\alu1/art/add/tout__1_carry__2_n_6 ),
        .I3(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I4(bdatr[13]),
        .I5(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .O(c1bus[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[13]_i_10 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[13]_i_11 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[13]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h3F303F30A0A0AFAF)) 
    \rgf_c1bus_wb[13]_i_12 
       (.I0(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[13]_i_13 
       (.I0(\rgf_c1bus_wb[13]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h8BAA)) 
    \rgf_c1bus_wb[13]_i_14 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c1bus_wb[13]_i_15 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hCC9FFF9F)) 
    \rgf_c1bus_wb[13]_i_16 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .I4(a1bus_0[1]),
        .O(\rgf_c1bus_wb[13]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[13]_i_17 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(a1bus_0[4]),
        .I3(a1bus_0[5]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0303F3F305F505F5)) 
    \rgf_c1bus_wb[13]_i_18 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\rgf/sreg/sr [6]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[13]_i_19 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[7]),
        .I2(a1bus_0[8]),
        .I3(a1bus_0[9]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[13]_i_2 
       (.I0(\rgf_c1bus_wb[13]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_6_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[13]_i_20 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[11]),
        .I2(a1bus_0[12]),
        .I3(a1bus_0[13]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_21 
       (.I0(a1bus_0[2]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[3]),
        .O(\rgf_c1bus_wb[13]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_22 
       (.I0(a1bus_0[6]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[7]),
        .O(\rgf_c1bus_wb[13]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_23 
       (.I0(a1bus_0[4]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[13]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_24 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[9]),
        .O(\rgf_c1bus_wb[13]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_25 
       (.I0(a1bus_0[10]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[11]),
        .O(\rgf_c1bus_wb[13]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hEAEAEAEAFFFFFFEA)) 
    \rgf_c1bus_wb[13]_i_3 
       (.I0(\rgf_c1bus_wb[13]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFCDCFCDFCCDCCCDF)) 
    \rgf_c1bus_wb[13]_i_4 
       (.I0(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hD0FFFFFFD0D0D0D0)) 
    \rgf_c1bus_wb[13]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(a1bus_0[12]),
        .I5(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFAFFEAEFAAAFEAE)) 
    \rgf_c1bus_wb[13]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[13]_i_7 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[13]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\bdatw[13]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[13]_i_9 
       (.I0(\bdatw[13]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(a1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF54)) 
    \rgf_c1bus_wb[14]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_2_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .O(c1bus[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_10 
       (.I0(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hAA8B)) 
    \rgf_c1bus_wb[14]_i_11 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c1bus_wb[14]_i_13 
       (.I0(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF70FF70707070)) 
    \rgf_c1bus_wb[14]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[14]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[14]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[14]_i_16 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[14]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\bdatw[15]_INST_0_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c1bus_wb[14]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[14]_i_19 
       (.I0(a1bus_0[14]),
        .I1(\bdatw[14]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBABABABBBA)) 
    \rgf_c1bus_wb[14]_i_2 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[14]_i_20 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\bdatw[14]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[14]_i_21 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(a1bus_0[13]),
        .I3(a1bus_0[14]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[14]_i_22 
       (.I0(a1bus_0[2]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[1]),
        .O(\rgf_c1bus_wb[14]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hA9)) 
    \rgf_c1bus_wb[14]_i_23 
       (.I0(\bdatw[9]_INST_0_i_13_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c1bus_wb[14]_i_24 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[14]_i_25 
       (.I0(a1bus_0[14]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[14]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0505F505F303F303)) 
    \rgf_c1bus_wb[14]_i_26 
       (.I0(a1bus_0[14]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[14]_i_27 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[2]),
        .I2(a1bus_0[3]),
        .I3(a1bus_0[4]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[14]_i_28 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[6]),
        .I2(a1bus_0[7]),
        .I3(a1bus_0[8]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[14]_i_29 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[10]),
        .I2(a1bus_0[11]),
        .I3(a1bus_0[12]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF880A)) 
    \rgf_c1bus_wb[14]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c1bus_wb[14]_i_30 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[14]_i_31 
       (.I0(\rgf/sreg/sr [6]),
        .I1(a1bus_0[0]),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[14]_i_32 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(a1bus_0[0]),
        .O(\rgf_c1bus_wb[14]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h44F4444444444444)) 
    \rgf_c1bus_wb[14]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I1(\alu1/art/add/tout__1_carry__2_n_5 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[14]),
        .O(\rgf_c1bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF5454FF54)) 
    \rgf_c1bus_wb[14]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \rgf_c1bus_wb[14]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h99A99999)) 
    \rgf_c1bus_wb[14]_i_7 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\bdatw[9]_INST_0_i_13_n_0 ),
        .I4(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF077F077F0FFF000)) 
    \rgf_c1bus_wb[14]_i_8 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[14]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4FFFFFFF4FFF4)) 
    \rgf_c1bus_wb[15]_i_1 
       (.I0(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I1(\alu1/art/p_0_in ),
        .I2(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I5(bdatr[15]),
        .O(c1bus[15]));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[15]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_25_n_0 ),
        .I2(\ctl1/stat [2]),
        .O(\rgf_c1bus_wb[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00400400)) 
    \rgf_c1bus_wb[15]_i_100 
       (.I0(\rgf_c1bus_wb[15]_i_102_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_30_n_0 ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [3]),
        .I5(\rgf_c1bus_wb[15]_i_103_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_100_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[15]_i_101 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_c1bus_wb[15]_i_101_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[15]_i_102 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .O(\rgf_c1bus_wb[15]_i_102_n_0 ));
  LUT6 #(
    .INIT(64'h0C040C0000000C00)) 
    \rgf_c1bus_wb[15]_i_103 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_c1bus_wb[15]_i_103_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[15]_i_11 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[15]_i_12 
       (.I0(\bdatw[15]_INST_0_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[15]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(a1bus_0[7]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hEEE00000)) 
    \rgf_c1bus_wb[15]_i_14 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I3(\bdatw[15]_INST_0_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hC0007800)) 
    \rgf_c1bus_wb[15]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I4(\bdatw[15]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[15]_i_16 
       (.I0(a1bus_0[14]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \rgf_c1bus_wb[15]_i_17 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[15]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5DFD)) 
    \rgf_c1bus_wb[15]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFE0000FFEF)) 
    \rgf_c1bus_wb[15]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(tout__1_carry_i_9__0_n_0),
        .I5(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0D0D000)) 
    \rgf_c1bus_wb[15]_i_20 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_33_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_34_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000222F)) 
    \rgf_c1bus_wb[15]_i_21 
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_36_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\rgf_c1bus_wb[15]_i_37_n_0 ),
        .I4(\fch/ir1 [15]),
        .I5(\ctl1/stat [2]),
        .O(\rgf_c1bus_wb[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAABAAABAAAAA)) 
    \rgf_c1bus_wb[15]_i_22 
       (.I0(\rgf_c1bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAA2220)) 
    \rgf_c1bus_wb[15]_i_23 
       (.I0(\rgf_c1bus_wb[15]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_44_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_45_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAAABAAAAAAAA)) 
    \rgf_c1bus_wb[15]_i_24 
       (.I0(\ctl1/stat [1]),
        .I1(\rgf_c1bus_wb[15]_i_46_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_47_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_48_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_49_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_50_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFBBB8BBB8)) 
    \rgf_c1bus_wb[15]_i_25 
       (.I0(\rgf_c1bus_wb[15]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_53_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_54_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_55_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_56_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[15]_i_26 
       (.I0(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAEAAAAAA)) 
    \rgf_c1bus_wb[15]_i_27 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(\bdatw[9]_INST_0_i_13_n_0 ),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[15]_i_28 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[11]),
        .I2(a1bus_0[12]),
        .I3(a1bus_0[13]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF20D)) 
    \rgf_c1bus_wb[15]_i_29 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\bdatw[10]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF54)) 
    \rgf_c1bus_wb[15]_i_3 
       (.I0(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[15]_i_30 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[7]),
        .I2(a1bus_0[8]),
        .I3(a1bus_0[9]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[15]_i_31 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(a1bus_0[4]),
        .I3(a1bus_0[5]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_32 
       (.I0(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_33 
       (.I0(\rgf_c1bus_wb[15]_i_59_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_60_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_61_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_62_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_34 
       (.I0(\rgf_c1bus_wb[15]_i_63_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_64_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_65_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hFF8A)) 
    \rgf_c1bus_wb[15]_i_35 
       (.I0(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFDDDDFFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_36 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [7]),
        .I4(\ctl1/stat [1]),
        .I5(\bcmd[0]_INST_0_i_23_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BABBBABA)) 
    \rgf_c1bus_wb[15]_i_37 
       (.I0(\rgf_c1bus_wb[15]_i_66_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_67_n_0 ),
        .I3(\fch/ir1 [7]),
        .I4(\ctl1/stat [1]),
        .I5(\rgf_c1bus_wb[15]_i_68_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \rgf_c1bus_wb[15]_i_38 
       (.I0(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [15]),
        .I5(\stat[0]_i_3__0_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFF0000FDFF000000)) 
    \rgf_c1bus_wb[15]_i_39 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [8]),
        .I3(\ctl1/stat [0]),
        .I4(\ctl1/stat [1]),
        .I5(\fch/ir1 [9]),
        .O(\rgf_c1bus_wb[15]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF8AAA)) 
    \rgf_c1bus_wb[15]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_19_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[15]_i_40 
       (.I0(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\ctl1/stat [0]),
        .I3(\ctl1/stat [1]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_c1bus_wb[15]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFBAAAAAAAA)) 
    \rgf_c1bus_wb[15]_i_41 
       (.I0(\fch/ir1 [11]),
        .I1(\rgf_c1bus_wb[15]_i_69_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [14]),
        .I4(\ctl1/stat [1]),
        .I5(\rgf_c1bus_wb[15]_i_70_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h0000001D00000013)) 
    \rgf_c1bus_wb[15]_i_42 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [8]),
        .I4(\ctl1/stat [1]),
        .I5(\fch/ir1 [6]),
        .O(\rgf_c1bus_wb[15]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[15]_i_43 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [8]),
        .O(\rgf_c1bus_wb[15]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFF90000FFFEFFFF)) 
    \rgf_c1bus_wb[15]_i_44 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\ctl1/stat [1]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_c1bus_wb[15]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_45 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [14]),
        .I5(\ctl1/stat [0]),
        .O(\rgf_c1bus_wb[15]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \rgf_c1bus_wb[15]_i_46 
       (.I0(\fch/ir1 [13]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [15]),
        .O(\rgf_c1bus_wb[15]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011710070)) 
    \rgf_c1bus_wb[15]_i_47 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [10]),
        .I5(\rgf_c1bus_wb[15]_i_71_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8AAA8A8)) 
    \rgf_c1bus_wb[15]_i_48 
       (.I0(\fch/ir1 [11]),
        .I1(\rgf_c1bus_wb[15]_i_72_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_73_n_0 ),
        .I3(\fadr[15]_INST_0_i_21_n_0 ),
        .I4(ctl_fetch1_fl_i_12_n_0),
        .I5(\ctl1/stat [0]),
        .O(\rgf_c1bus_wb[15]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF7F3FFF3FFF)) 
    \rgf_c1bus_wb[15]_i_49 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [12]),
        .I2(\stat[0]_i_3__0_n_0 ),
        .I3(\fch/ir1 [13]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [15]),
        .O(\rgf_c1bus_wb[15]_i_49_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[15]_i_5 
       (.I0(\mem/read_cyc [2]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [3]),
        .O(\rgf_c1bus_wb[15]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hEEEAEEEE)) 
    \rgf_c1bus_wb[15]_i_50 
       (.I0(\rgf_c1bus_wb[15]_i_74_n_0 ),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [15]),
        .O(\rgf_c1bus_wb[15]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h4444455545554444)) 
    \rgf_c1bus_wb[15]_i_51 
       (.I0(\rgf_c1bus_wb[15]_i_75_n_0 ),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [15]),
        .I4(\rgf_c1bus_wb[15]_i_76_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\rgf_c1bus_wb[15]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000002FFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_52 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat [1]),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [13]),
        .O(\rgf_c1bus_wb[15]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFF3C30)) 
    \rgf_c1bus_wb[15]_i_53 
       (.I0(\rgf_c1bus_wb[15]_i_77_n_0 ),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [12]),
        .I4(\ctl1/stat [1]),
        .I5(\fch/ir1 [14]),
        .O(\rgf_c1bus_wb[15]_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF5554)) 
    \rgf_c1bus_wb[15]_i_54 
       (.I0(\fch/ir1 [12]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [15]),
        .O(\rgf_c1bus_wb[15]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0222)) 
    \rgf_c1bus_wb[15]_i_55 
       (.I0(\rgf_c1bus_wb[15]_i_78_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [1]),
        .I4(\rgf_c1bus_wb[15]_i_79_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_80_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0D0D0F000D0D0)) 
    \rgf_c1bus_wb[15]_i_56 
       (.I0(\rgf_c1bus_wb[15]_i_81_n_0 ),
        .I1(\bcmd[0]_INST_0_i_24_n_0 ),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [2]),
        .I4(\ctl1/stat [1]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_c1bus_wb[15]_i_56_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_57 
       (.I0(a1bus_0[0]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[1]),
        .O(\rgf_c1bus_wb[15]_i_57_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c1bus_wb[15]_i_58 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[15]_i_58_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_59 
       (.I0(a1bus_0[13]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[12]),
        .O(\rgf_c1bus_wb[15]_i_59_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[15]_i_6 
       (.I0(\ctl1/stat [2]),
        .I1(tout__1_carry_i_12_n_0),
        .I2(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_60 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[15]_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_61 
       (.I0(a1bus_0[9]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[8]),
        .O(\rgf_c1bus_wb[15]_i_61_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_62 
       (.I0(a1bus_0[11]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[10]),
        .O(\rgf_c1bus_wb[15]_i_62_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_63 
       (.I0(a1bus_0[5]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[4]),
        .O(\rgf_c1bus_wb[15]_i_63_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_64 
       (.I0(a1bus_0[7]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[6]),
        .O(\rgf_c1bus_wb[15]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[15]_i_65 
       (.I0(a1bus_0[3]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .O(\rgf_c1bus_wb[15]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hF00FF002F00FF00F)) 
    \rgf_c1bus_wb[15]_i_66 
       (.I0(\rgf_c1bus_wb[15]_i_82_n_0 ),
        .I1(\bdatw[15]_INST_0_i_279_n_0 ),
        .I2(\ctl1/stat [0]),
        .I3(\ctl1/stat [1]),
        .I4(ctl_fetch1_fl_i_11_n_0),
        .I5(\rgf_c1bus_wb[15]_i_83_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF7FFFFF)) 
    \rgf_c1bus_wb[15]_i_67 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_c1bus_wb[15]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf_c1bus_wb[15]_i_68 
       (.I0(\rgf_c1bus_wb[15]_i_78_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [2]),
        .I5(\rgf_c1bus_wb[15]_i_84_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0F3FFF0F1F0F1)) 
    \rgf_c1bus_wb[15]_i_69 
       (.I0(\bdatw[15]_INST_0_i_276_n_0 ),
        .I1(\fch/ir1 [12]),
        .I2(\rgf_c1bus_wb[15]_i_85_n_0 ),
        .I3(\fch/ir1 [13]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [15]),
        .O(\rgf_c1bus_wb[15]_i_69_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFD00FFFF)) 
    \rgf_c1bus_wb[15]_i_70 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\badr[15]_INST_0_i_298_n_0 ),
        .I2(\badr[15]_INST_0_i_297_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_35_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I5(\badr[15]_INST_0_i_296_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_70_n_0 ));
  LUT5 #(
    .INIT(32'hCECECDDD)) 
    \rgf_c1bus_wb[15]_i_71 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [10]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [6]),
        .O(\rgf_c1bus_wb[15]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h000000000040FF00)) 
    \rgf_c1bus_wb[15]_i_72 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [5]),
        .I5(\rgf_c1bus_wb[15]_i_86_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h00FE001100000505)) 
    \rgf_c1bus_wb[15]_i_73 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [10]),
        .O(\rgf_c1bus_wb[15]_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA88AA88AAAA8A)) 
    \rgf_c1bus_wb[15]_i_74 
       (.I0(\rgf_c1bus_wb[15]_i_87_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_88_n_0 ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [1]),
        .O(\rgf_c1bus_wb[15]_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \rgf_c1bus_wb[15]_i_75 
       (.I0(\rgf_selc1_wb[1]_i_16_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I2(\stat[1]_i_18__0_n_0 ),
        .I3(\fch/ir1 [0]),
        .I4(\ctl1/stat [1]),
        .I5(\rgf_selc1_wb[1]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h00005AAACFCFCFCF)) 
    \rgf_c1bus_wb[15]_i_76 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [14]),
        .O(\rgf_c1bus_wb[15]_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h5515551555550000)) 
    \rgf_c1bus_wb[15]_i_77 
       (.I0(\rgf_c1bus_wb[15]_i_89_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\badr[15]_INST_0_i_294_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_90_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_91_n_0 ),
        .I5(\ctl1/stat [1]),
        .O(\rgf_c1bus_wb[15]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_c1bus_wb[15]_i_78 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [4]),
        .O(\rgf_c1bus_wb[15]_i_78_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \rgf_c1bus_wb[15]_i_79 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [10]),
        .I4(\rgf_c1bus_wb[15]_i_92_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_79_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[15]_i_8 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF77FFFF0003)) 
    \rgf_c1bus_wb[15]_i_80 
       (.I0(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_93_n_0 ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [15]),
        .I5(\ctl1/stat [1]),
        .O(\rgf_c1bus_wb[15]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h0222000002220222)) 
    \rgf_c1bus_wb[15]_i_81 
       (.I0(\fch/ir1 [10]),
        .I1(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [11]),
        .O(\rgf_c1bus_wb[15]_i_81_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[15]_i_82 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_c1bus_wb[15]_i_82_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[15]_i_83 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .O(\rgf_c1bus_wb[15]_i_83_n_0 ));
  LUT5 #(
    .INIT(32'hFFC0C088)) 
    \rgf_c1bus_wb[15]_i_84 
       (.I0(\ctl1/stat [0]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .O(\rgf_c1bus_wb[15]_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F0F07000D00)) 
    \rgf_c1bus_wb[15]_i_85 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .I2(\rgf_c1bus_wb[15]_i_94_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [10]),
        .O(\rgf_c1bus_wb[15]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hFFF7FFF7FFFFFFF7)) 
    \rgf_c1bus_wb[15]_i_86 
       (.I0(\bcmd[0]_INST_0_i_7_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\ctl1/stat [0]),
        .I3(\rgf_c1bus_wb[15]_i_43_n_0 ),
        .I4(\stat[0]_i_21__0_n_0 ),
        .I5(\fch/ir1 [4]),
        .O(\rgf_c1bus_wb[15]_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7753030)) 
    \rgf_c1bus_wb[15]_i_87 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [11]),
        .I4(\rgf_c1bus_wb[15]_i_95_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_96_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFF)) 
    \rgf_c1bus_wb[15]_i_88 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [4]),
        .I2(\fadr[15]_INST_0_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_97_n_0 ),
        .I4(\ctl1/stat [2]),
        .I5(\fch/ir1 [2]),
        .O(\rgf_c1bus_wb[15]_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000020200002200)) 
    \rgf_c1bus_wb[15]_i_89 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_c1bus_wb[15]_i_89_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[15]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hBE)) 
    \rgf_c1bus_wb[15]_i_90 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [11]),
        .O(\rgf_c1bus_wb[15]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF8)) 
    \rgf_c1bus_wb[15]_i_91 
       (.I0(\rgf_selc1_wb[0]_i_20_n_0 ),
        .I1(\stat[0]_i_21__0_n_0 ),
        .I2(\fch/ir1 [6]),
        .I3(\rgf_c1bus_wb[15]_i_98_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_99_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_100_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBEEEEB3BBEEEE)) 
    \rgf_c1bus_wb[15]_i_92 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [11]),
        .I5(\rgf_c1bus_wb[15]_i_101_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_92_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_93 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [6]),
        .O(\rgf_c1bus_wb[15]_i_93_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFEFFFEFFFF)) 
    \rgf_c1bus_wb[15]_i_94 
       (.I0(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I1(\fch/ir1 [15]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_c1bus_wb[15]_i_94_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFFFFFF)) 
    \rgf_c1bus_wb[15]_i_95 
       (.I0(\fch/ir1 [8]),
        .I1(\fadr[15]_INST_0_i_21_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\badr[15]_INST_0_i_297_n_0 ),
        .I5(\fch/ir1 [2]),
        .O(\rgf_c1bus_wb[15]_i_95_n_0 ));
  LUT6 #(
    .INIT(64'hEEEFEEEEEEEEEEEF)) 
    \rgf_c1bus_wb[15]_i_96 
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [13]),
        .I3(\rgf_selc1_wb[1]_i_16_n_0 ),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [1]),
        .O(\rgf_c1bus_wb[15]_i_96_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFDFFFF)) 
    \rgf_c1bus_wb[15]_i_97 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\stat[0]_i_34_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h8888AA880888AA88)) 
    \rgf_c1bus_wb[15]_i_98 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [4]),
        .O(\rgf_c1bus_wb[15]_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h0322033303020333)) 
    \rgf_c1bus_wb[15]_i_99 
       (.I0(\fch/ir1 [7]),
        .I1(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [11]),
        .O(\rgf_c1bus_wb[15]_i_99_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[1]_i_1 
       (.I0(\rgf_c1bus_wb[1]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I2(\alu1/art/add/tout__1_carry_n_6 ),
        .I3(\rgf_c1bus_wb[1]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_4_n_0 ),
        .O(c1bus[1]));
  LUT6 #(
    .INIT(64'h44417741447D777D)) 
    \rgf_c1bus_wb[1]_i_10 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\bdatw[8]_INST_0_i_14_n_0 ),
        .I4(a1bus_0[13]),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[1]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[1]_i_11 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[1]_i_12 
       (.I0(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[1]_i_13 
       (.I0(\rgf_c1bus_wb[5]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h5555FFF7)) 
    \rgf_c1bus_wb[1]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h000000001F100000)) 
    \rgf_c1bus_wb[1]_i_15 
       (.I0(\rgf_c1bus_wb[3]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000E200)) 
    \rgf_c1bus_wb[1]_i_16 
       (.I0(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[1]_i_17 
       (.I0(\rgf_c1bus_wb[12]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[1]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[1]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[1]_i_19 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF0E)) 
    \rgf_c1bus_wb[1]_i_2 
       (.I0(\rgf_c1bus_wb[1]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_7_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[1]_i_20 
       (.I0(a1bus_0[6]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[1]_i_3 
       (.I0(\mem/read_cyc [0]),
        .I1(bdatr[9]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[1]),
        .O(\rgf_c1bus_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF6A880000)) 
    \rgf_c1bus_wb[1]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\bdatw[9]_INST_0_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c1bus_wb[1]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0511051105000555)) 
    \rgf_c1bus_wb[1]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEEFAAAAA)) 
    \rgf_c1bus_wb[1]_i_7 
       (.I0(\rgf_c1bus_wb[1]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFE00FE000000FE00)) 
    \rgf_c1bus_wb[1]_i_8 
       (.I0(\rgf_c1bus_wb[1]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_16_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h33FF23FF03FF2323)) 
    \rgf_c1bus_wb[1]_i_9 
       (.I0(a1bus_0[9]),
        .I1(\rgf_c1bus_wb[1]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I5(\bdatw[9]_INST_0_i_13_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[2]_i_1 
       (.I0(\rgf_c1bus_wb[2]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I2(\alu1/art/add/tout__1_carry_n_5 ),
        .I3(\rgf_c1bus_wb[2]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_4_n_0 ),
        .O(c1bus[2]));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_c1bus_wb[2]_i_10 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[2]_i_11 
       (.I0(a1bus_0[10]),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c1bus_wb[2]_i_12 
       (.I0(a1bus_0[2]),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h2E)) 
    \rgf_c1bus_wb[2]_i_13 
       (.I0(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[2]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h050305F3)) 
    \rgf_c1bus_wb[2]_i_14 
       (.I0(\rgf_c1bus_wb[12]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[2]_i_15 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h55335533000FFF0F)) 
    \rgf_c1bus_wb[2]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_59_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_60_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[2]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(a1bus_0[2]),
        .O(\rgf_c1bus_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF0E000E)) 
    \rgf_c1bus_wb[2]_i_2 
       (.I0(\rgf_c1bus_wb[2]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_7_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[2]_i_3 
       (.I0(\mem/read_cyc [0]),
        .I1(bdatr[10]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[2]),
        .O(\rgf_c1bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00541154)) 
    \rgf_c1bus_wb[2]_i_4 
       (.I0(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00CF444400CF4F4F)) 
    \rgf_c1bus_wb[2]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \rgf_c1bus_wb[2]_i_6 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF80B0)) 
    \rgf_c1bus_wb[2]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFACAC0C0)) 
    \rgf_c1bus_wb[2]_i_8 
       (.I0(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h02000202FFFFFFFF)) 
    \rgf_c1bus_wb[2]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_17_n_0 ),
        .I3(\bdatw[10]_INST_0_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF10111010)) 
    \rgf_c1bus_wb[3]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_2_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_5_n_0 ),
        .O(c1bus[3]));
  LUT4 #(
    .INIT(16'hB8BB)) 
    \rgf_c1bus_wb[3]_i_10 
       (.I0(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I3(a1bus_0[15]),
        .O(\rgf_c1bus_wb[3]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[3]_i_11 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hCAFA)) 
    \rgf_c1bus_wb[3]_i_12 
       (.I0(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABAAA)) 
    \rgf_c1bus_wb[3]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFABEEAB)) 
    \rgf_c1bus_wb[3]_i_14 
       (.I0(\rgf_c1bus_wb[3]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[3]_i_15 
       (.I0(\mem/read_cyc [0]),
        .I1(bdatr[11]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[3]),
        .O(\rgf_c1bus_wb[3]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[3]_i_16 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[3]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[3]_i_17 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[3]_i_18 
       (.I0(a1bus_0[14]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[13]),
        .O(\rgf_c1bus_wb[3]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h02000202FFFFFFFF)) 
    \rgf_c1bus_wb[3]_i_19 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_22_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hCACC00000A0C0000)) 
    \rgf_c1bus_wb[3]_i_2 
       (.I0(\rgf_c1bus_wb[3]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_c1bus_wb[3]_i_20 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[3]_i_21 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[3]_i_22 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(a1bus_0[3]),
        .O(\rgf_c1bus_wb[3]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF3200)) 
    \rgf_c1bus_wb[3]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \rgf_c1bus_wb[3]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF5D)) 
    \rgf_c1bus_wb[3]_i_5 
       (.I0(\rgf_c1bus_wb[3]_i_14_n_0 ),
        .I1(\alu1/art/add/tout__1_carry_n_4 ),
        .I2(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[3]_i_6 
       (.I0(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF101FFFF)) 
    \rgf_c1bus_wb[3]_i_7 
       (.I0(\rgf_c1bus_wb[3]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[3]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[3]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[4]_i_1 
       (.I0(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I2(\alu1/art/add/tout__1_carry__0_n_7 ),
        .I3(\rgf_c1bus_wb[4]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .O(c1bus[4]));
  LUT6 #(
    .INIT(64'h1F5F1F5F115F1155)) 
    \rgf_c1bus_wb[4]_i_10 
       (.I0(\rgf_c1bus_wb[4]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[4]_i_11 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0F5F5FFF0F3F3)) 
    \rgf_c1bus_wb[4]_i_12 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000001D000000)) 
    \rgf_c1bus_wb[4]_i_13 
       (.I0(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAFFFFEFFF)) 
    \rgf_c1bus_wb[4]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[4]_i_15 
       (.I0(a1bus_0[4]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[4]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[4]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[4]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000222E2222)) 
    \rgf_c1bus_wb[4]_i_2 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[4]_i_3 
       (.I0(\mem/read_cyc [0]),
        .I1(bdatr[12]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[4]),
        .O(\rgf_c1bus_wb[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF9020B000)) 
    \rgf_c1bus_wb[4]_i_4 
       (.I0(a1bus_0[4]),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA028AAAAAAAAA)) 
    \rgf_c1bus_wb[4]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hA8080000)) 
    \rgf_c1bus_wb[4]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[4]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[4]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[4]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c1bus_wb[5]_i_1 
       (.I0(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I2(\alu1/art/add/tout__1_carry__0_n_6 ),
        .I3(\rgf_c1bus_wb[5]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_4_n_0 ),
        .O(c1bus[5]));
  LUT6 #(
    .INIT(64'h00000000AFC0A0CF)) 
    \rgf_c1bus_wb[5]_i_10 
       (.I0(\bdatw[13]_INST_0_i_16_n_0 ),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(a1bus_0[5]),
        .I5(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h2A888000)) 
    \rgf_c1bus_wb[5]_i_11 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(\bdatw[13]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(a1bus_0[5]),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[5]_i_12 
       (.I0(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000151FFFFFFFF)) 
    \rgf_c1bus_wb[5]_i_13 
       (.I0(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[5]_i_14 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[4]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[5]_i_15 
       (.I0(\rgf_c1bus_wb[5]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_16 
       (.I0(a1bus_0[11]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[12]),
        .O(\rgf_c1bus_wb[5]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_17 
       (.I0(a1bus_0[12]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[11]),
        .O(\rgf_c1bus_wb[5]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_18 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[7]),
        .O(\rgf_c1bus_wb[5]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_19 
       (.I0(a1bus_0[10]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[9]),
        .O(\rgf_c1bus_wb[5]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002F20202)) 
    \rgf_c1bus_wb[5]_i_2 
       (.I0(\rgf_c1bus_wb[5]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC000C080C0004000)) 
    \rgf_c1bus_wb[5]_i_3 
       (.I0(\mem/read_cyc [1]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [3]),
        .I3(bdatr[5]),
        .I4(\mem/read_cyc [0]),
        .I5(bdatr[13]),
        .O(\rgf_c1bus_wb[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0D02000)) 
    \rgf_c1bus_wb[5]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hDFDCDFDFDCDCDCDF)) 
    \rgf_c1bus_wb[5]_i_5 
       (.I0(\rgf_c1bus_wb[5]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF54045555)) 
    \rgf_c1bus_wb[5]_i_6 
       (.I0(\rgf_c1bus_wb[5]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hB8FF0000B8000000)) 
    \rgf_c1bus_wb[5]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBABABABFAAAAAAAA)) 
    \rgf_c1bus_wb[5]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_9 
       (.I0(\bdatw[13]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00BA0010FFFFFFFF)) 
    \rgf_c1bus_wb[6]_i_1 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_5_n_0 ),
        .O(c1bus[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00541154)) 
    \rgf_c1bus_wb[6]_i_10 
       (.I0(\rgf_c1bus_wb[6]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hE0F0000040000000)) 
    \rgf_c1bus_wb[6]_i_11 
       (.I0(\mem/read_cyc [0]),
        .I1(bdatr[14]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[6]),
        .O(\rgf_c1bus_wb[6]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[6]_i_12 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[6]_i_13 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[9]),
        .I2(a1bus_0[10]),
        .I3(a1bus_0[11]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[6]_i_14 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h02000202FFFFFFFF)) 
    \rgf_c1bus_wb[6]_i_15 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_18_n_0 ),
        .I3(\bdatw[14]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \rgf_c1bus_wb[6]_i_16 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h882A0080)) 
    \rgf_c1bus_wb[6]_i_17 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\bdatw[14]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[6]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(a1bus_0[6]),
        .O(\rgf_c1bus_wb[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h22223330AAAAFFFF)) 
    \rgf_c1bus_wb[6]_i_2 
       (.I0(\rgf_c1bus_wb[6]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[6]_i_3 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h03113300)) 
    \rgf_c1bus_wb[6]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h1101)) 
    \rgf_c1bus_wb[6]_i_5 
       (.I0(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_11_n_0 ),
        .I2(\alu1/art/add/tout__1_carry__0_n_5 ),
        .I3(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[6]_i_6 
       (.I0(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[6]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_c1bus_wb[6]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[6]_i_9 
       (.I0(\rgf_c1bus_wb[6]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4544)) 
    \rgf_c1bus_wb[7]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .O(c1bus[7]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_10 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[7]_i_11 
       (.I0(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF00DF00FF00FF00)) 
    \rgf_c1bus_wb[7]_i_12 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[7]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c1bus_wb[7]_i_13 
       (.I0(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[7]_i_14 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c1bus_wb[7]_i_15 
       (.I0(\mem/read_cyc [1]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [3]),
        .O(\rgf_c1bus_wb[7]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hAABE)) 
    \rgf_c1bus_wb[7]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(a1bus_0[7]),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h22200020)) 
    \rgf_c1bus_wb[7]_i_18 
       (.I0(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(a1bus_0[7]),
        .I3(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I4(\bdatw[15]_INST_0_i_18_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h2AA08000)) 
    \rgf_c1bus_wb[7]_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I2(\bdatw[15]_INST_0_i_18_n_0 ),
        .I3(a1bus_0[7]),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FFACFF00FFFF)) 
    \rgf_c1bus_wb[7]_i_2 
       (.I0(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[7]_i_20 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[5]),
        .I2(a1bus_0[6]),
        .I3(a1bus_0[7]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[7]_i_21 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[8]),
        .I2(a1bus_0[9]),
        .I3(a1bus_0[10]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[7]_i_22 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_c1bus_wb[7]_i_3 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8F888F8F8F888F88)) 
    \rgf_c1bus_wb[7]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h22F2FFFF22F222F2)) 
    \rgf_c1bus_wb[7]_i_5 
       (.I0(\rgf_c0bus_wb[7]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(bdatr[7]),
        .I3(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I5(\alu1/art/add/tout__1_carry__0_n_4 ),
        .O(\rgf_c1bus_wb[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF510000)) 
    \rgf_c1bus_wb[7]_i_6 
       (.I0(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[7]_i_7 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[10]),
        .I2(a1bus_0[11]),
        .I3(a1bus_0[12]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \rgf_c1bus_wb[7]_i_8 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\rgf/sreg/sr [6]),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h5D555DDD)) 
    \rgf_c1bus_wb[7]_i_9 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45554050)) 
    \rgf_c1bus_wb[8]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_2_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .O(c1bus[8]));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[8]_i_10 
       (.I0(a1bus_0[7]),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[8]_i_11 
       (.I0(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[8]_i_12 
       (.I0(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF54FF54FFFFFF54)) 
    \rgf_c1bus_wb[8]_i_13 
       (.I0(\rgf_c1bus_wb[8]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[8]_i_14 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[9]),
        .I2(a1bus_0[10]),
        .I3(a1bus_0[11]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c1bus_wb[8]_i_15 
       (.I0(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[8]_i_16 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[4]),
        .I2(a1bus_0[5]),
        .I3(a1bus_0[6]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[8]_i_17 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[8]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[8]_i_18 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h9020B000)) 
    \rgf_c1bus_wb[8]_i_19 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8]_INST_0_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[8]_i_2 
       (.I0(\bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c1bus_wb[8]_i_20 
       (.I0(a1bus_0[8]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hAEEE)) 
    \rgf_c1bus_wb[8]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hCC80CCCCCC80CC80)) 
    \rgf_c1bus_wb[8]_i_4 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[8]_i_5 
       (.I0(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .I1(bdatr[8]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(\alu1/art/add/tout__1_carry__1_n_7 ),
        .I4(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[8]_i_6 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[6]),
        .I2(a1bus_0[7]),
        .I3(a1bus_0[8]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h333300FF55550F0F)) 
    \rgf_c1bus_wb[8]_i_7 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[2]),
        .I2(a1bus_0[3]),
        .I3(a1bus_0[4]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFDFFF)) 
    \rgf_c1bus_wb[8]_i_8 
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\bdatw[10]_INST_0_i_14_n_0 ),
        .I3(a1bus_0[0]),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[8]_i_9 
       (.I0(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF10111010)) 
    \rgf_c1bus_wb[9]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_2_n_0 ),
        .I2(\bdatw[12]_INST_0_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_5_n_0 ),
        .O(c1bus[9]));
  LUT4 #(
    .INIT(16'h5404)) 
    \rgf_c1bus_wb[9]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFF5C005C00000000)) 
    \rgf_c1bus_wb[9]_i_11 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[9]_i_12 
       (.I0(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAEAEFFFFFFAE)) 
    \rgf_c1bus_wb[9]_i_13 
       (.I0(\rgf_c1bus_wb[9]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[9]_i_14 
       (.I0(a1bus_0[1]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[0]),
        .O(\rgf_c1bus_wb[9]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[9]_i_15 
       (.I0(a1bus_0[13]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[9]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[9]_i_16 
       (.I0(a1bus_0[15]),
        .I1(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h3A)) 
    \rgf_c1bus_wb[9]_i_17 
       (.I0(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_58_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0F0F555500FF3333)) 
    \rgf_c1bus_wb[9]_i_18 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[5]),
        .I2(a1bus_0[6]),
        .I3(a1bus_0[7]),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\bdatw[8]_INST_0_i_14_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h535300FF)) 
    \rgf_c1bus_wb[9]_i_19 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(\bdatw[8]_INST_0_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_57_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFE00FE000000FE00)) 
    \rgf_c1bus_wb[9]_i_2 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\bdatw[11]_INST_0_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hC06000C0)) 
    \rgf_c1bus_wb[9]_i_20 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I3(\bdatw[9]_INST_0_i_2_n_0 ),
        .I4(a1bus_0[9]),
        .O(\rgf_c1bus_wb[9]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \rgf_c1bus_wb[9]_i_21 
       (.I0(a1bus_0[9]),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[9]_i_22 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDFFD)) 
    \rgf_c1bus_wb[9]_i_23 
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(a1bus_0[9]),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h70FF7070)) 
    \rgf_c1bus_wb[9]_i_3 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF101F1010)) 
    \rgf_c1bus_wb[9]_i_4 
       (.I0(\rgf_c1bus_wb[9]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \rgf_c1bus_wb[9]_i_5 
       (.I0(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .I1(bdatr[9]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(\alu1/art/add/tout__1_carry__1_n_6 ),
        .I4(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h5455)) 
    \rgf_c1bus_wb[9]_i_6 
       (.I0(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hE020)) 
    \rgf_c1bus_wb[9]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[9]_i_8 
       (.I0(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \rgf_c1bus_wb[9]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c1bus_wb_reg[0]_i_4 
       (.I0(\rgf_c1bus_wb[0]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_11_n_0 ),
        .O(\rgf_c1bus_wb_reg[0]_i_4_n_0 ),
        .S(\rgf_c1bus_wb[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5555510055555555)) 
    \rgf_selc0_rn_wb[0]_i_1 
       (.I0(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_4_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_5_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h5555FFFFF3FFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_10 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [6]),
        .I3(brdy),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[0]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \rgf_selc0_rn_wb[0]_i_11 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [10]),
        .O(\rgf_selc0_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDDFFFFFFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_12 
       (.I0(\rgf_selc0_rn_wb[0]_i_20_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .I2(brdy),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [1]),
        .I5(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc0_rn_wb[0]_i_13 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000601000)) 
    \rgf_selc0_rn_wb[0]_i_14 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [3]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [2]),
        .I5(\fadr[15]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFEAAA)) 
    \rgf_selc0_rn_wb[0]_i_15 
       (.I0(\rgf_selc0_rn_wb[0]_i_23_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\ccmd[4]_INST_0_i_13_n_0 ),
        .I3(crdy),
        .I4(\fch/ir0 [11]),
        .I5(\rgf_selc0_rn_wb[0]_i_24_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000032C0)) 
    \rgf_selc0_rn_wb[0]_i_16 
       (.I0(brdy),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [0]),
        .I5(\fadr[15]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FBAE0000)) 
    \rgf_selc0_rn_wb[0]_i_17 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [12]),
        .I2(\rgf/sreg/sr [4]),
        .I3(\fch/ir0 [11]),
        .I4(\ccmd[1]_INST_0_i_21_n_0 ),
        .I5(\stat[0]_i_24_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[0]_i_18 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [14]),
        .O(\rgf_selc0_rn_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFF009696FFFF6666)) 
    \rgf_selc0_rn_wb[0]_i_19 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir0 [11]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\rgf_selc0_rn_wb[0]_i_25_n_0 ),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [12]),
        .O(\rgf_selc0_rn_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAA8A)) 
    \rgf_selc0_rn_wb[0]_i_2 
       (.I0(\ctl0/stat [2]),
        .I1(\ctl0/stat [1]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [15]),
        .I4(\fadr[15]_INST_0_i_14_n_0 ),
        .I5(\fadr[15]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[0]_i_20 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_rn_wb[0]_i_21 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [7]),
        .O(\rgf_selc0_rn_wb[0]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc0_rn_wb[0]_i_22 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .O(\rgf_selc0_rn_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFF0E0000FF0C0000)) 
    \rgf_selc0_rn_wb[0]_i_23 
       (.I0(\ccmd[0]_INST_0_i_30_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_26_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .I4(\fch/ir0 [10]),
        .I5(crdy),
        .O(\rgf_selc0_rn_wb[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h4F0F0F0F4FFF0F0F)) 
    \rgf_selc0_rn_wb[0]_i_24 
       (.I0(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_29_n_0 ),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [11]),
        .I5(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000AA2AAAAAAAAA)) 
    \rgf_selc0_rn_wb[0]_i_25 
       (.I0(\rgf_selc0_rn_wb[0]_i_30_n_0 ),
        .I1(\fch/ir0 [0]),
        .I2(\stat[0]_i_8__1_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_31_n_0 ),
        .I5(\stat[0]_i_7__1_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_26 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [7]),
        .O(\rgf_selc0_rn_wb[0]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h20000000)) 
    \rgf_selc0_rn_wb[0]_i_27 
       (.I0(brdy),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [3]),
        .O(\rgf_selc0_rn_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h08080C0000000C00)) 
    \rgf_selc0_rn_wb[0]_i_28 
       (.I0(crdy),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [3]),
        .O(\rgf_selc0_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h7F7DFFFFFFFDFFFF)) 
    \rgf_selc0_rn_wb[0]_i_29 
       (.I0(\rgf_selc0_rn_wb[0]_i_32_n_0 ),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [3]),
        .I5(\rgf_selc0_rn_wb[0]_i_33_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFEEAEFFBFFFBF)) 
    \rgf_selc0_rn_wb[0]_i_3 
       (.I0(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I5(\fch/ir0 [0]),
        .O(\rgf_selc0_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h57770000FFFFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_30 
       (.I0(\rgf_selc0_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_34_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I3(crdy),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(\fch/ir0 [3]),
        .O(\rgf_selc0_rn_wb[0]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hF008000C0008000C)) 
    \rgf_selc0_rn_wb[0]_i_31 
       (.I0(crdy),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .I5(\rgf_selc0_wb[1]_i_18_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc0_rn_wb[0]_i_32 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[0]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_rn_wb[0]_i_33 
       (.I0(\fch/ir0 [0]),
        .I1(brdy),
        .O(\rgf_selc0_rn_wb[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \rgf_selc0_rn_wb[0]_i_34 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [8]),
        .I4(crdy),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \rgf_selc0_rn_wb[0]_i_4 
       (.I0(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [11]),
        .I4(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_5 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [15]),
        .O(\rgf_selc0_rn_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0404040404040400)) 
    \rgf_selc0_rn_wb[0]_i_6 
       (.I0(\fch/ir0 [15]),
        .I1(\ctl0/stat [0]),
        .I2(\ctl0/stat [1]),
        .I3(\rgf_selc0_rn_wb[0]_i_15_n_0 ),
        .I4(\ctl0/stat [2]),
        .I5(\rgf_selc0_rn_wb[0]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h45454500FFFFFFFF)) 
    \rgf_selc0_rn_wb[0]_i_7 
       (.I0(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_19_n_0 ),
        .I5(\ccmd[4]_INST_0_i_8_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hBFFF)) 
    \rgf_selc0_rn_wb[0]_i_8 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [14]),
        .O(\rgf_selc0_rn_wb[0]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[0]_i_9 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .O(\rgf_selc0_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00007555)) 
    \rgf_selc0_rn_wb[1]_i_1 
       (.I0(\rgf_selc0_rn_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I2(\ccmd[4]_INST_0_i_8_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\ctl0/stat [2]),
        .I5(\rgf_selc0_rn_wb[1]_i_3_n_0 ),
        .O(ctl_selc0_rn));
  LUT6 #(
    .INIT(64'hA080808020000000)) 
    \rgf_selc0_rn_wb[1]_i_10 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [1]),
        .O(\rgf_selc0_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0202030000000300)) 
    \rgf_selc0_rn_wb[1]_i_11 
       (.I0(crdy),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [4]),
        .O(\rgf_selc0_rn_wb[1]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf_selc0_rn_wb[1]_i_12 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[1]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h44400040)) 
    \rgf_selc0_rn_wb[1]_i_13 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [4]),
        .O(\rgf_selc0_rn_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0040FFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_14 
       (.I0(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I1(\fch/ir0 [4]),
        .I2(\stat[0]_i_7__1_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .I4(\ctl0/stat [0]),
        .I5(\rgf_selc0_rn_wb[1]_i_19_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0083)) 
    \rgf_selc0_rn_wb[1]_i_15 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [11]),
        .O(\rgf_selc0_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h15555555FFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_16 
       (.I0(crdy),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [8]),
        .I5(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFE0FFFF)) 
    \rgf_selc0_rn_wb[1]_i_17 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [11]),
        .O(\rgf_selc0_rn_wb[1]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[1]_i_18 
       (.I0(\fch/ir0 [8]),
        .I1(crdy),
        .O(\rgf_selc0_rn_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFB73FBFBFFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_19 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [1]),
        .I2(\rgf_selc0_rn_wb[1]_i_20_n_0 ),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [6]),
        .I5(\stat[2]_i_10_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFF45FFFF)) 
    \rgf_selc0_rn_wb[1]_i_2 
       (.I0(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I1(\fadr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I3(\fch/ir0 [15]),
        .I4(\ctl0/stat [1]),
        .O(\rgf_selc0_rn_wb[1]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFF7E)) 
    \rgf_selc0_rn_wb[1]_i_20 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [3]),
        .O(\rgf_selc0_rn_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF10FFD0)) 
    \rgf_selc0_rn_wb[1]_i_3 
       (.I0(\rgf_selc0_rn_wb[1]_i_6_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [10]),
        .I3(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_9_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFF400F4)) 
    \rgf_selc0_rn_wb[1]_i_4 
       (.I0(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I1(\fch/ir0 [1]),
        .I2(\stat[0]_i_29__0_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\rgf_selc0_rn_wb[1]_i_10_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0028)) 
    \rgf_selc0_rn_wb[1]_i_5 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .O(\rgf_selc0_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_6 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [6]),
        .I2(brdy),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .I5(\rgf_selc0_rn_wb[1]_i_11_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF555555D55555)) 
    \rgf_selc0_rn_wb[1]_i_7 
       (.I0(\ctl0/stat [0]),
        .I1(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .I2(brdy),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [4]),
        .I5(\stat[0]_i_29__0_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0D000F0FDDDDFFFF)) 
    \rgf_selc0_rn_wb[1]_i_8 
       (.I0(\fch/ir0 [3]),
        .I1(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I2(crdy),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [1]),
        .I5(\rgf_selc0_rn_wb[1]_i_13_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hBBABAAAABBBBBBBB)) 
    \rgf_selc0_rn_wb[1]_i_9 
       (.I0(\badrx[15]_INST_0_i_5_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_14_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_15_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(\fch/ir0 [4]),
        .O(\rgf_selc0_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0040004000405555)) 
    \rgf_selc0_rn_wb[2]_i_1 
       (.I0(\ctl0/stat [2]),
        .I1(\fch/ir0 [10]),
        .I2(\ccmd[4]_INST_0_i_8_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I4(\ccmd[3]_INST_0_i_3_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_3_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080CC8000)) 
    \rgf_selc0_rn_wb[2]_i_10 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [8]),
        .I2(crdy),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [9]),
        .O(\rgf_selc0_rn_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_11 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .I2(brdy),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h7F5F7FFF7FFF7FFF)) 
    \rgf_selc0_rn_wb[2]_i_12 
       (.I0(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I5(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h5D00FFFF50005000)) 
    \rgf_selc0_rn_wb[2]_i_13 
       (.I0(\fch/ir0 [8]),
        .I1(crdy),
        .I2(\fch/ir0 [7]),
        .I3(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hA888888888888888)) 
    \rgf_selc0_rn_wb[2]_i_14 
       (.I0(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I1(crdy),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [6]),
        .O(\rgf_selc0_rn_wb[2]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hBFEFFFEF)) 
    \rgf_selc0_rn_wb[2]_i_15 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [6]),
        .O(\rgf_selc0_rn_wb[2]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc0_rn_wb[2]_i_16 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [11]),
        .O(\rgf_selc0_rn_wb[2]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \rgf_selc0_rn_wb[2]_i_2 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .O(\rgf_selc0_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFF4FF04FFF40F040)) 
    \rgf_selc0_rn_wb[2]_i_3 
       (.I0(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I2(\ctl0/stat [0]),
        .I3(\ctl0/stat [1]),
        .I4(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF88F800F000F0)) 
    \rgf_selc0_rn_wb[2]_i_4 
       (.I0(brdy),
        .I1(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I4(\stat[0]_i_29__0_n_0 ),
        .I5(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5515FFFFFFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_5 
       (.I0(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [3]),
        .I3(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\rgf_selc0_rn_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2022AAAAA8AA)) 
    \rgf_selc0_rn_wb[2]_i_6 
       (.I0(\rgf_selc0_rn_wb[2]_i_12_n_0 ),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [11]),
        .I5(crdy),
        .O(\rgf_selc0_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00BF00BF000000BF)) 
    \rgf_selc0_rn_wb[2]_i_7 
       (.I0(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I1(\fch/ir0 [2]),
        .I2(\stat[2]_i_10_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_13_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00000880)) 
    \rgf_selc0_rn_wb[2]_i_8 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [6]),
        .O(\rgf_selc0_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF47CF)) 
    \rgf_selc0_rn_wb[2]_i_9 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [2]),
        .I3(crdy),
        .I4(\fch/ir0 [11]),
        .I5(\rgf_selc0_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    rgf_selc0_stat_i_1
       (.I0(fch_term),
        .I1(rst_n),
        .O(rgf_selc0_stat_i_1_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc0_stat_i_2
       (.I0(ctl_selc0),
        .I1(\rgf_selc0_wb[0]_i_1_n_0 ),
        .O(rgf_selc0_stat_i_2_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc0_stat_i_3
       (.I0(fch_wrbufn0),
        .O(\rgf/rctl/p_2_in ));
  LUT5 #(
    .INIT(32'hFFFF8880)) 
    rgf_selc0_stat_i_4
       (.I0(\ir0_id_fl[20]_i_2_n_0 ),
        .I1(\fch/rst_n_fl ),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/ir0_id_fl [20]),
        .I4(\fch/fch_irq_req_fl ),
        .O(fch_wrbufn0));
  LUT6 #(
    .INIT(64'h4544454445444545)) 
    \rgf_selc0_wb[0]_i_1 
       (.I0(\ctl0/stat [2]),
        .I1(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_3_n_0 ),
        .I4(\rgf_selc0_wb[0]_i_4_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_5_n_0 ),
        .O(\rgf_selc0_wb[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0051515511515155)) 
    \rgf_selc0_wb[0]_i_10 
       (.I0(\rgf_selc0_wb[0]_i_15_n_0 ),
        .I1(\ccmd[4]_INST_0_i_14_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\ctl0/stat [0]),
        .I4(crdy),
        .I5(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\rgf_selc0_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7F7FAAAA3737AAFF)) 
    \rgf_selc0_wb[0]_i_11 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [8]),
        .I2(crdy),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [7]),
        .O(\rgf_selc0_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFF77BF76)) 
    \rgf_selc0_wb[0]_i_12 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [3]),
        .O(\rgf_selc0_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    \rgf_selc0_wb[0]_i_13 
       (.I0(\rgf_selc0_wb[0]_i_16_n_0 ),
        .I1(\ccmd[4]_INST_0_i_22_n_0 ),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [8]),
        .I4(brdy),
        .I5(\rgf_selc0_wb[0]_i_17_n_0 ),
        .O(\rgf_selc0_wb[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[0]_i_14 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .O(\rgf_selc0_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0140010000400000)) 
    \rgf_selc0_wb[0]_i_15 
       (.I0(\ccmd[4]_INST_0_i_16_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [6]),
        .I4(brdy),
        .I5(\fch/ir0 [7]),
        .O(\rgf_selc0_wb[0]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h01FF)) 
    \rgf_selc0_wb[0]_i_16 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [9]),
        .O(\rgf_selc0_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00550055C0550055)) 
    \rgf_selc0_wb[0]_i_17 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [4]),
        .O(\rgf_selc0_wb[0]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0010)) 
    \rgf_selc0_wb[0]_i_2 
       (.I0(\ccmd[4]_INST_0_i_12_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I4(\rgf_selc0_wb[0]_i_7_n_0 ),
        .O(\rgf_selc0_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h40400000404000FF)) 
    \rgf_selc0_wb[0]_i_3 
       (.I0(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I1(\stat[0]_i_18__0_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_9_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_10_n_0 ),
        .I4(\ctl0/stat [1]),
        .I5(\fch/ir0 [11]),
        .O(\rgf_selc0_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0002AAAA0000AAA0)) 
    \rgf_selc0_wb[0]_i_4 
       (.I0(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [9]),
        .I5(\ctl0/stat [0]),
        .O(\rgf_selc0_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBFFFFFFFB)) 
    \rgf_selc0_wb[0]_i_5 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [11]),
        .I2(\ccmd[4]_INST_0_i_16_n_0 ),
        .I3(\ctl0/stat [0]),
        .I4(\rgf_selc0_wb[0]_i_12_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_13_n_0 ),
        .O(\rgf_selc0_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc0_wb[0]_i_6 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .I3(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0100111110110111)) 
    \rgf_selc0_wb[0]_i_7 
       (.I0(\ccmd[3]_INST_0_i_8_n_0 ),
        .I1(\ctl0/stat [1]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [12]),
        .O(\rgf_selc0_wb[0]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc0_wb[0]_i_8 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [7]),
        .O(\rgf_selc0_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hCFCC1111)) 
    \rgf_selc0_wb[0]_i_9 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [6]),
        .I3(brdy),
        .I4(\fch/ir0 [11]),
        .O(\rgf_selc0_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF000D0F0D)) 
    \rgf_selc0_wb[1]_i_1 
       (.I0(\rgf_selc0_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I2(\ctl0/stat [2]),
        .I3(\ctl0/stat [1]),
        .I4(\rgf_selc0_wb[1]_i_4_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_5_n_0 ),
        .O(ctl_selc0));
  LUT6 #(
    .INIT(64'hEEEEEEEEEFEEEEEE)) 
    \rgf_selc0_wb[1]_i_10 
       (.I0(\rgf_selc0_wb[1]_i_26_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I2(\fch/ir0 [14]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir0 [11]),
        .I5(\ctl0/stat [0]),
        .O(\rgf_selc0_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBAABBAAAAAABAAA)) 
    \rgf_selc0_wb[1]_i_11 
       (.I0(\rgf_selc0_wb[1]_i_28_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_29_n_0 ),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [12]),
        .I4(\rgf_selc0_wb[1]_i_30_n_0 ),
        .I5(\fch/ir0 [15]),
        .O(\rgf_selc0_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000045FF000045)) 
    \rgf_selc0_wb[1]_i_12 
       (.I0(\bdatw[15]_INST_0_i_21_n_0 ),
        .I1(\ccmd[1]_INST_0_i_11_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_31_n_0 ),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [14]),
        .I5(\ctl0/stat [0]),
        .O(\rgf_selc0_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h77F7000077F777F7)) 
    \rgf_selc0_wb[1]_i_13 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [14]),
        .I2(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I3(\stat[0]_i_29__0_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_32_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .O(\rgf_selc0_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEFFFFFFFFF)) 
    \rgf_selc0_wb[1]_i_14 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .I4(brdy),
        .I5(\fch/ir0 [11]),
        .O(\rgf_selc0_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \rgf_selc0_wb[1]_i_15 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [12]),
        .I5(\ctl0/stat [0]),
        .O(\rgf_selc0_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \rgf_selc0_wb[1]_i_16 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\ctl0/stat [2]),
        .I3(\ccmd[4]_INST_0_i_18_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [0]),
        .O(\rgf_selc0_wb[1]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc0_wb[1]_i_17 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [12]),
        .O(\rgf_selc0_wb[1]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc0_wb[1]_i_18 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [4]),
        .O(\rgf_selc0_wb[1]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_wb[1]_i_19 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAAAABABABAB)) 
    \rgf_selc0_wb[1]_i_2 
       (.I0(\ccmd[3]_INST_0_i_3_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_7_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_8_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_9_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\rgf_selc0_wb[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h80008080)) 
    \rgf_selc0_wb[1]_i_20 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .O(\rgf_selc0_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h222200000000FF0F)) 
    \rgf_selc0_wb[1]_i_21 
       (.I0(brdy),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(crdy),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [8]),
        .O(\rgf_selc0_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAA0A2A2A0E0A0A0B)) 
    \rgf_selc0_wb[1]_i_22 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [4]),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [3]),
        .O(\rgf_selc0_wb[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[1]_i_23 
       (.I0(brdy),
        .I1(\fch/ir0 [6]),
        .O(\rgf_selc0_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h05C5C5C505C50505)) 
    \rgf_selc0_wb[1]_i_24 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [7]),
        .I2(\ctl0/stat [0]),
        .I3(brdy),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [6]),
        .O(\rgf_selc0_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h4440000444400000)) 
    \rgf_selc0_wb[1]_i_25 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [3]),
        .O(\rgf_selc0_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AFBFFFAF)) 
    \rgf_selc0_wb[1]_i_26 
       (.I0(\rgf_selc0_wb[1]_i_33_n_0 ),
        .I1(\rgf/sreg/sr [4]),
        .I2(\ccmd[1]_INST_0_i_21_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .I5(\rgf_selc0_wb[1]_i_34_n_0 ),
        .O(\rgf_selc0_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000101)) 
    \rgf_selc0_wb[1]_i_27 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(\ccmd[0]_INST_0_i_23_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [3]),
        .I5(\rgf_selc0_wb[1]_i_35_n_0 ),
        .O(\rgf_selc0_wb[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4444104544441044)) 
    \rgf_selc0_wb[1]_i_28 
       (.I0(\rgf_selc0_wb[1]_i_36_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [13]),
        .O(\rgf_selc0_wb[1]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_29 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [14]),
        .O(\rgf_selc0_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55450000)) 
    \rgf_selc0_wb[1]_i_3 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [2]),
        .I2(\ctl0/stat [0]),
        .I3(brdy),
        .I4(\rgf_selc0_wb[1]_i_10_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_11_n_0 ),
        .O(\rgf_selc0_wb[1]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_selc0_wb[1]_i_30 
       (.I0(\fch/ir0 [11]),
        .I1(\rgf/sreg/sr [7]),
        .O(\rgf_selc0_wb[1]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h8FAF)) 
    \rgf_selc0_wb[1]_i_31 
       (.I0(\fch/ir0 [1]),
        .I1(\ctl0/stat [0]),
        .I2(\fch/ir0 [0]),
        .I3(brdy),
        .O(\rgf_selc0_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \rgf_selc0_wb[1]_i_32 
       (.I0(\ccmd[0]_INST_0_i_23_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [3]),
        .I5(\rgf_selc0_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_wb[1]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_selc0_wb[1]_i_33 
       (.I0(\ccmd[1]_INST_0_i_11_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_37_n_0 ),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [12]),
        .I5(\rgf_selc0_wb[1]_i_38_n_0 ),
        .O(\rgf_selc0_wb[1]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hBAABABBAABBAABBA)) 
    \rgf_selc0_wb[1]_i_34 
       (.I0(\ctl0/stat [0]),
        .I1(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir0 [11]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\fch/ir0 [12]),
        .O(\rgf_selc0_wb[1]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFDFDFFF)) 
    \rgf_selc0_wb[1]_i_35 
       (.I0(\stat[2]_i_14_n_0 ),
        .I1(\bdatw[15]_INST_0_i_21_n_0 ),
        .I2(\ctl0/stat [0]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [1]),
        .I5(\rgf_selc0_wb[1]_i_39_n_0 ),
        .O(\rgf_selc0_wb[1]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_36 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [12]),
        .O(\rgf_selc0_wb[1]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc0_wb[1]_i_37 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[1]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_selc0_wb[1]_i_38 
       (.I0(\fch/ir0 [8]),
        .I1(crdy),
        .I2(\fch/ir0 [9]),
        .O(\rgf_selc0_wb[1]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc0_wb[1]_i_39 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [12]),
        .O(\rgf_selc0_wb[1]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFEF0000FFEFFFEF)) 
    \rgf_selc0_wb[1]_i_4 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [15]),
        .I2(\rgf_selc0_wb[1]_i_12_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_13_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_15_n_0 ),
        .O(\rgf_selc0_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000002000000000)) 
    \rgf_selc0_wb[1]_i_5 
       (.I0(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\ctl0/stat [1]),
        .I5(\bdatw[8]_INST_0_i_15_n_0 ),
        .O(\rgf_selc0_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0004550400040004)) 
    \rgf_selc0_wb[1]_i_6 
       (.I0(\rgf_selc0_wb[1]_i_19_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_20_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\ctl0/stat [0]),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_21_n_0 ),
        .O(\rgf_selc0_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAA0CAA0000000000)) 
    \rgf_selc0_wb[1]_i_7 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(\bcmd[0]_INST_0_i_26_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [10]),
        .I5(crdy),
        .O(\rgf_selc0_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0001C07F0001403F)) 
    \rgf_selc0_wb[1]_i_8 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [9]),
        .I5(crdy),
        .O(\rgf_selc0_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF773F)) 
    \rgf_selc0_wb[1]_i_9 
       (.I0(\rgf_selc0_wb[1]_i_22_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(\rgf_selc0_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_25_n_0 ),
        .O(\rgf_selc0_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF04)) 
    \rgf_selc1_rn_wb[0]_i_1 
       (.I0(\rgf_selc1_rn_wb[0]_i_2_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_4_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(ctl_selc1_rn[0]));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[0]_i_10 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h40F0000000000000)) 
    \rgf_selc1_rn_wb[0]_i_11 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .I1(brdy),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [1]),
        .I4(\bdatw[8]_INST_0_i_59_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \rgf_selc1_rn_wb[0]_i_12 
       (.I0(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h3FFFFFFFFFFFAAFF)) 
    \rgf_selc1_rn_wb[0]_i_13 
       (.I0(\fch/ir1 [4]),
        .I1(\stat[0]_i_7__0_n_0 ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [6]),
        .O(\rgf_selc1_rn_wb[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_14 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF4FFFFFFFFFFF4FF)) 
    \rgf_selc1_rn_wb[0]_i_15 
       (.I0(\rgf_selc1_rn_wb[0]_i_21_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_22_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h3F2A3F3F3F2A3F00)) 
    \rgf_selc1_rn_wb[0]_i_16 
       (.I0(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [14]),
        .I5(\stat[0]_i_22_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h08000800C8000800)) 
    \rgf_selc1_rn_wb[0]_i_17 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_24_n_0 ),
        .I2(\stat[0]_i_7__0_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_26_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF08008088)) 
    \rgf_selc1_rn_wb[0]_i_18 
       (.I0(\stat[2]_i_5__0_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [13]),
        .I5(\rgf_selc1_rn_wb[0]_i_28_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[0]_i_19 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .O(\rgf_selc1_rn_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000D5DD)) 
    \rgf_selc1_rn_wb[0]_i_2 
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_11_n_0 ),
        .I5(\ctl1/stat [0]),
        .O(\rgf_selc1_rn_wb[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc1_rn_wb[0]_i_20 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [6]),
        .O(\rgf_selc1_rn_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_21 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[0]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_rn_wb[0]_i_22 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [3]),
        .O(\rgf_selc1_rn_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA200A2A2)) 
    \rgf_selc1_rn_wb[0]_i_23 
       (.I0(\badr[15]_INST_0_i_238_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_29_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_30_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_30_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_selc1_rn_wb[0]_i_24 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [1]),
        .O(\rgf_selc1_rn_wb[0]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h54)) 
    \rgf_selc1_rn_wb[0]_i_25 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [3]),
        .O(\rgf_selc1_rn_wb[0]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_selc1_rn_wb[0]_i_26 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [2]),
        .O(\rgf_selc1_rn_wb[0]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_27 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat [0]),
        .O(\rgf_selc1_rn_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \rgf_selc1_rn_wb[0]_i_28 
       (.I0(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .I1(\stat[0]_i_32__0_n_0 ),
        .I2(\ctl1/stat [1]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [11]),
        .I5(\badr[15]_INST_0_i_245_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF3F2BFFEFFFEFFFF)) 
    \rgf_selc1_rn_wb[0]_i_29 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [0]),
        .O(\rgf_selc1_rn_wb[0]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_3 
       (.I0(\ctl1/stat [1]),
        .I1(\fch/ir1 [15]),
        .O(\rgf_selc1_rn_wb[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_selc1_rn_wb[0]_i_30 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[0]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \rgf_selc1_rn_wb[0]_i_31 
       (.I0(\fch/ir1 [2]),
        .I1(\ctl1/stat [2]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [3]),
        .I4(\fadr[15]_INST_0_i_18_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_rn_wb[0]_i_32 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAAA882AAAAAAAAAA)) 
    \rgf_selc1_rn_wb[0]_i_4 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [0]),
        .I5(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h02AAAAAA02AA02AA)) 
    \rgf_selc1_rn_wb[0]_i_5 
       (.I0(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_13_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I5(\fch/ir1 [3]),
        .O(\rgf_selc1_rn_wb[0]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF01)) 
    \rgf_selc1_rn_wb[0]_i_6 
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [0]),
        .I2(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .I3(\ctl1/stat [2]),
        .I4(\rgf_selc1_rn_wb[0]_i_17_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[0]_i_7 
       (.I0(\ctl1/stat [2]),
        .I1(\rgf_selc1_rn_wb[0]_i_18_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF7FFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_8 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [0]),
        .O(\rgf_selc1_rn_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5C5FFFFF5F5FFFFF)) 
    \rgf_selc1_rn_wb[0]_i_9 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [7]),
        .I5(\stat[0]_i_7__0_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5454545444544444)) 
    \rgf_selc1_rn_wb[1]_i_1 
       (.I0(\ctl1/stat [2]),
        .I1(\rgf_selc1_rn_wb[1]_i_2_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I4(\fch/ir1 [4]),
        .I5(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0E0F0F0F0F0F0F0F)) 
    \rgf_selc1_rn_wb[1]_i_10 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [12]),
        .O(\rgf_selc1_rn_wb[1]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_11 
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [0]),
        .O(\rgf_selc1_rn_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8A88AAAAAAAAAAAA)) 
    \rgf_selc1_rn_wb[1]_i_12 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0080AAAA00800080)) 
    \rgf_selc1_rn_wb[1]_i_13 
       (.I0(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I2(\bcmd[0]_INST_0_i_23_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I5(\fch/ir1 [4]),
        .O(\rgf_selc1_rn_wb[1]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00002800)) 
    \rgf_selc1_rn_wb[1]_i_14 
       (.I0(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [0]),
        .O(\rgf_selc1_rn_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5FFFFFF7EFFFF)) 
    \rgf_selc1_rn_wb[1]_i_15 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0FF7CFC00FFFF)) 
    \rgf_selc1_rn_wb[1]_i_16 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45444444)) 
    \rgf_selc1_rn_wb[1]_i_2 
       (.I0(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I2(\fch/ir1 [6]),
        .I3(\stat[0]_i_7__0_n_0 ),
        .I4(\fch/ir1 [4]),
        .I5(\rgf_selc1_rn_wb[1]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_selc1_rn_wb[1]_i_3 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat [1]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [15]),
        .O(\rgf_selc1_rn_wb[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h54555555)) 
    \rgf_selc1_rn_wb[1]_i_4 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .I3(brdy),
        .I4(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h3000FFFF3000BA00)) 
    \rgf_selc1_rn_wb[1]_i_5 
       (.I0(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_8_n_0 ),
        .I2(\stat[0]_i_7__0_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\rgf_selc1_rn_wb[1]_i_9_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0FFFFFF)) 
    \rgf_selc1_rn_wb[1]_i_6 
       (.I0(\fch/ir1 [1]),
        .I1(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_10_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_11_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_12_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF800F800F800)) 
    \rgf_selc1_rn_wb[1]_i_7 
       (.I0(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_144_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_14_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[1]_i_8 
       (.I0(ctl_fetch1_fl_i_11_n_0),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [8]),
        .I5(\bdatw[11]_INST_0_i_27_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_selc1_rn_wb[1]_i_9 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF0D0000)) 
    \rgf_selc1_rn_wb[2]_i_1 
       (.I0(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_3_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_5_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_7_n_0 ),
        .O(ctl_selc1_rn[2]));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[2]_i_10 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_11 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [2]),
        .I2(ctl_fetch1_fl_i_11_n_0),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [6]),
        .I5(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_selc1_rn_wb[2]_i_12 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [2]),
        .O(\rgf_selc1_rn_wb[2]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc1_rn_wb[2]_i_13 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[2]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_rn_wb[2]_i_14 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[2]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF000D)) 
    \rgf_selc1_rn_wb[2]_i_15 
       (.I0(\fch/ir1 [2]),
        .I1(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[2]_i_16 
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [2]),
        .O(\rgf_selc1_rn_wb[2]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h28AA2AAA)) 
    \rgf_selc1_rn_wb[2]_i_17 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h8808CCCC08080CCC)) 
    \rgf_selc1_rn_wb[2]_i_18 
       (.I0(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_23_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[2]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[2]_i_19 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFF7FFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_2 
       (.I0(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I1(brdy),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\fch/ir1 [5]),
        .O(\rgf_selc1_rn_wb[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \rgf_selc1_rn_wb[2]_i_20 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F2F2F200F2F2)) 
    \rgf_selc1_rn_wb[2]_i_21 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [2]),
        .I2(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\ctl1/stat [1]),
        .I5(\ctl1/stat [0]),
        .O(\rgf_selc1_rn_wb[2]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFBEFD55FFFEFD55)) 
    \rgf_selc1_rn_wb[2]_i_22 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [6]),
        .O(\rgf_selc1_rn_wb[2]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_23 
       (.I0(\rgf_selc1_rn_wb[2]_i_24_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [2]),
        .O(\rgf_selc1_rn_wb[2]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFF77BF76)) 
    \rgf_selc1_rn_wb[2]_i_24 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [3]),
        .O(\rgf_selc1_rn_wb[2]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h3000FFFF3000BA00)) 
    \rgf_selc1_rn_wb[2]_i_3 
       (.I0(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I2(\stat[0]_i_7__0_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\rgf_selc1_rn_wb[2]_i_12_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_rn_wb[2]_i_4 
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [0]),
        .O(\rgf_selc1_rn_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0008)) 
    \rgf_selc1_rn_wb[2]_i_5 
       (.I0(\fch/ir1 [5]),
        .I1(brdy),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \rgf_selc1_rn_wb[2]_i_6 
       (.I0(\ctl1/stat [2]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [15]),
        .O(\rgf_selc1_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h8080808080FF8080)) 
    \rgf_selc1_rn_wb[2]_i_7 
       (.I0(\fch/ir1 [10]),
        .I1(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I4(\bcmd[2]_INST_0_i_4_n_0 ),
        .I5(\ctl1/stat [0]),
        .O(\rgf_selc1_rn_wb[2]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h6000)) 
    \rgf_selc1_rn_wb[2]_i_8 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \rgf_selc1_rn_wb[2]_i_9 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc1_stat_i_1
       (.I0(ctl_selc1),
        .I1(\rgf_selc1_wb[0]_i_1_n_0 ),
        .O(rgf_selc1_stat_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc1_stat_i_2
       (.I0(fch_wrbufn1),
        .O(rgf_selc1_stat_i_2_n_0));
  LUT5 #(
    .INIT(32'h54554444)) 
    \rgf_selc1_wb[0]_i_1 
       (.I0(\ctl1/stat [2]),
        .I1(\rgf_selc1_wb[0]_i_2_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_5_n_0 ),
        .O(\rgf_selc1_wb[0]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hDDD0DDDDEEEEEEEE)) 
    \rgf_selc1_wb[0]_i_10 
       (.I0(\fch/ir1 [8]),
        .I1(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I2(\fch/ir1 [6]),
        .I3(\bcmd[2]_INST_0_i_1_n_0 ),
        .I4(brdy),
        .I5(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[0]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFBFFF)) 
    \rgf_selc1_wb[0]_i_11 
       (.I0(\ctl1/stat [0]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .O(\rgf_selc1_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AABA0000)) 
    \rgf_selc1_wb[0]_i_12 
       (.I0(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(brdy),
        .I3(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_18_n_0 ),
        .O(\rgf_selc1_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBFF0FF5FBFF0FFF0)) 
    \rgf_selc1_wb[0]_i_13 
       (.I0(\fch/ir1 [6]),
        .I1(\stat[0]_i_7__0_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_wb[0]_i_14 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [14]),
        .O(\rgf_selc1_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h333F333333337777)) 
    \rgf_selc1_wb[0]_i_15 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [9]),
        .I2(\rgf_selc1_rn_wb[2]_i_24_n_0 ),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [10]),
        .O(\rgf_selc1_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h77777777FFFF7FFF)) 
    \rgf_selc1_wb[0]_i_16 
       (.I0(\fch/ir1 [8]),
        .I1(\ctl1/stat [0]),
        .I2(\rgf_selc1_wb[0]_i_19_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_20_n_0 ),
        .I4(\fch/ir1 [4]),
        .I5(\rgf_selc1_wb[0]_i_21_n_0 ),
        .O(\rgf_selc1_wb[0]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[0]_i_17 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat [1]),
        .O(\rgf_selc1_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h030F033F0C0C0100)) 
    \rgf_selc1_wb[0]_i_18 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [7]),
        .I5(\ctl1/stat [0]),
        .O(\rgf_selc1_wb[0]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc1_wb[0]_i_19 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF8F8F8F8FFF8F8F8)) 
    \rgf_selc1_wb[0]_i_2 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_7_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_9_n_0 ),
        .I4(\fch/ir1 [14]),
        .I5(\ctl1/stat [1]),
        .O(\rgf_selc1_wb[0]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_wb[0]_i_20 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[0]_i_21 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1111F111)) 
    \rgf_selc1_wb[0]_i_3 
       (.I0(\rgf_selc1_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I3(\ctl1/stat [0]),
        .I4(\ctl1/stat [1]),
        .I5(\rgf_selc1_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_wb[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFFFB)) 
    \rgf_selc1_wb[0]_i_4 
       (.I0(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\ctl1/stat [1]),
        .I3(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[0]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \rgf_selc1_wb[0]_i_5 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [15]),
        .O(\rgf_selc1_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0440)) 
    \rgf_selc1_wb[0]_i_6 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [1]),
        .O(\rgf_selc1_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_selc1_wb[0]_i_7 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [15]),
        .I4(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0808880800080808)) 
    \rgf_selc1_wb[0]_i_8 
       (.I0(\fch/ir1 [15]),
        .I1(\badr[15]_INST_0_i_144_n_0 ),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [12]),
        .O(\rgf_selc1_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h10001100)) 
    \rgf_selc1_wb[0]_i_9 
       (.I0(\fch/ir1 [12]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0F0FDF0FFF0FD)) 
    \rgf_selc1_wb[1]_i_1 
       (.I0(\rgf_selc1_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_4_n_0 ),
        .I3(\ctl1/stat [2]),
        .I4(\ctl1/stat [1]),
        .I5(\rgf_selc1_wb[1]_i_5_n_0 ),
        .O(ctl_selc1));
  LUT6 #(
    .INIT(64'hEFECEFEFEFEFEFEC)) 
    \rgf_selc1_wb[1]_i_10 
       (.I0(\fch/ir1 [15]),
        .I1(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [11]),
        .I5(\rgf/sreg/sr [7]),
        .O(\rgf_selc1_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000E00000F0F)) 
    \rgf_selc1_wb[1]_i_11 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\rgf_selc1_wb[1]_i_31_n_0 ),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [13]),
        .I5(\ctl1/stat [0]),
        .O(\rgf_selc1_wb[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h3C333F31)) 
    \rgf_selc1_wb[1]_i_12 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [11]),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_selc1_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_selc1_wb[1]_i_13 
       (.I0(\rgf_selc1_wb[1]_i_32_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [4]),
        .I5(\fadr[15]_INST_0_i_19_n_0 ),
        .O(\rgf_selc1_wb[1]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFBFF)) 
    \rgf_selc1_wb[1]_i_14 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [3]),
        .I3(\ctl1/stat [0]),
        .O(\rgf_selc1_wb[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc1_wb[1]_i_15 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [12]),
        .O(\rgf_selc1_wb[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_wb[1]_i_16 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [15]),
        .O(\rgf_selc1_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFE0FFE)) 
    \rgf_selc1_wb[1]_i_17 
       (.I0(\bdatw[15]_INST_0_i_42_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [12]),
        .I4(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .O(\rgf_selc1_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h2FFF2F2F28282828)) 
    \rgf_selc1_wb[1]_i_18 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [1]),
        .I3(\ctl1/stat [0]),
        .I4(\stat[0]_i_7__0_n_0 ),
        .I5(\fch/ir1 [0]),
        .O(\rgf_selc1_wb[1]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFF8)) 
    \rgf_selc1_wb[1]_i_19 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [13]),
        .O(\rgf_selc1_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF11105555)) 
    \rgf_selc1_wb[1]_i_2 
       (.I0(\rgf_selc1_wb[1]_i_6_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_7_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_8_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_9_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\rgf_selc1_wb[1]_i_10_n_0 ),
        .O(\rgf_selc1_wb[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_wb[1]_i_20 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [13]),
        .O(\rgf_selc1_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000F20000)) 
    \rgf_selc1_wb[1]_i_21 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [15]),
        .I4(\rgf_selc1_wb[1]_i_34_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_35_n_0 ),
        .O(\rgf_selc1_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFAAAAFFEF)) 
    \rgf_selc1_wb[1]_i_22 
       (.I0(\rgf_selc1_wb[1]_i_36_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\ctl1/stat [0]),
        .I5(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .O(\rgf_selc1_wb[1]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_selc1_wb[1]_i_23 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[1]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h13)) 
    \rgf_selc1_wb[1]_i_24 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .O(\rgf_selc1_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA0A3A0A0)) 
    \rgf_selc1_wb[1]_i_25 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [7]),
        .I4(\stat[0]_i_13__0_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_38_n_0 ),
        .O(\rgf_selc1_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h88880000AAFB0000)) 
    \rgf_selc1_wb[1]_i_26 
       (.I0(\rgf_selc1_wb[1]_i_39_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [10]),
        .I5(\ctl1/stat [0]),
        .O(\rgf_selc1_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF7FBBBF7F)) 
    \rgf_selc1_wb[1]_i_27 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [3]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [4]),
        .O(\rgf_selc1_wb[1]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hFF7E)) 
    \rgf_selc1_wb[1]_i_28 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .O(\rgf_selc1_wb[1]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_wb[1]_i_29 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .O(\rgf_selc1_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAEAFAAABAAAB)) 
    \rgf_selc1_wb[1]_i_3 
       (.I0(\rgf_selc1_wb[1]_i_11_n_0 ),
        .I1(\fch/ir1 [12]),
        .I2(\ctl1/stat [0]),
        .I3(\rgf_selc1_wb[1]_i_12_n_0 ),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [15]),
        .O(\rgf_selc1_wb[1]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_wb[1]_i_30 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .O(\rgf_selc1_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAAFB)) 
    \rgf_selc1_wb[1]_i_31 
       (.I0(\rgf_selc1_wb[1]_i_40_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\rgf_selc1_wb[1]_i_41_n_0 ),
        .O(\rgf_selc1_wb[1]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[1]_i_32 
       (.I0(\ctl1/stat [1]),
        .I1(\fch/ir1 [15]),
        .O(\rgf_selc1_wb[1]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc1_wb[1]_i_33 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [7]),
        .I5(\fadr[15]_INST_0_i_21_n_0 ),
        .O(\rgf_selc1_wb[1]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_34 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .O(\rgf_selc1_wb[1]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFFFFFFFFFFFF)) 
    \rgf_selc1_wb[1]_i_35 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[1]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_wb[1]_i_36 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [10]),
        .O(\rgf_selc1_wb[1]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_wb[1]_i_37 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[1]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h1001)) 
    \rgf_selc1_wb[1]_i_38 
       (.I0(\fch/ir1 [14]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [11]),
        .I3(\rgf/sreg/sr [7]),
        .O(\rgf_selc1_wb[1]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc1_wb[1]_i_39 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [5]),
        .O(\rgf_selc1_wb[1]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \rgf_selc1_wb[1]_i_4 
       (.I0(\rgf_selc1_wb[1]_i_13_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_14_n_0 ),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [7]),
        .I5(\rgf_selc1_wb[1]_i_15_n_0 ),
        .O(\rgf_selc1_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB8B8B888)) 
    \rgf_selc1_wb[1]_i_40 
       (.I0(\rgf_selc1_wb[1]_i_42_n_0 ),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [11]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\ctl1/stat [0]),
        .O(\rgf_selc1_wb[1]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FF0040)) 
    \rgf_selc1_wb[1]_i_41 
       (.I0(\fch/ir1 [14]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [11]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [15]),
        .I5(\rgf_selc1_wb[1]_i_43_n_0 ),
        .O(\rgf_selc1_wb[1]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h9666)) 
    \rgf_selc1_wb[1]_i_42 
       (.I0(\fch/ir1 [11]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [7]),
        .O(\rgf_selc1_wb[1]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \rgf_selc1_wb[1]_i_43 
       (.I0(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I1(\bdatw[9]_INST_0_i_20_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_44_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_45_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_46_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_47_n_0 ),
        .O(\rgf_selc1_wb[1]_i_43_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_wb[1]_i_44 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [0]),
        .O(\rgf_selc1_wb[1]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_45 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [10]),
        .O(\rgf_selc1_wb[1]_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_selc1_wb[1]_i_46 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [1]),
        .O(\rgf_selc1_wb[1]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc1_wb[1]_i_47 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .I4(\badr[15]_INST_0_i_296_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[1]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEEFFEF)) 
    \rgf_selc1_wb[1]_i_5 
       (.I0(\rgf_selc1_wb[1]_i_16_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_17_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_20_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_21_n_0 ),
        .O(\rgf_selc1_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55550040)) 
    \rgf_selc1_wb[1]_i_6 
       (.I0(\rgf_selc1_wb[1]_i_22_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I2(brdy),
        .I3(\bcmd[2]_INST_0_i_1_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_25_n_0 ),
        .O(\rgf_selc1_wb[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h41115113)) 
    \rgf_selc1_wb[1]_i_7 
       (.I0(\fch/ir1 [9]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h3323333300003000)) 
    \rgf_selc1_wb[1]_i_8 
       (.I0(\fch/ir1 [10]),
        .I1(\rgf_selc1_wb[1]_i_26_n_0 ),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [6]),
        .I4(\stat[0]_i_7__0_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_27_n_0 ),
        .O(\rgf_selc1_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h40004040FFFFFFFF)) 
    \rgf_selc1_wb[1]_i_9 
       (.I0(\fch/ir1 [7]),
        .I1(\rgf_selc1_wb[1]_i_28_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [3]),
        .I4(\ctl1/stat [0]),
        .I5(\rgf_selc1_wb[1]_i_29_n_0 ),
        .O(\rgf_selc1_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[0]_i_1 
       (.I0(\sp[0]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [0]),
        .I4(\rgf/rgf_c1bus_0 [0]),
        .O(\sp[0]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFD08)) 
    \sp[0]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [0]),
        .I2(\sp[15]_i_6_n_0 ),
        .I3(\rgf/sptr/sp [0]),
        .O(\sp[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[10]_i_1 
       (.I0(\sp[10]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [10]),
        .I4(\rgf/rgf_c1bus_0 [10]),
        .O(\sp[10]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[10]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/sptr/sp [10]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [10]),
        .O(\sp[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[11]_i_1 
       (.I0(\sp[11]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [11]),
        .I4(\rgf/rgf_c1bus_0 [11]),
        .O(\sp[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[11]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/sptr/sp [11]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [11]),
        .O(\sp[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[12]_i_1 
       (.I0(\sp[12]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [12]),
        .I4(\rgf/rgf_c1bus_0 [12]),
        .O(\sp[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[12]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/sptr/sp [12]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [12]),
        .O(\sp[12]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[13]_i_1 
       (.I0(\sp[13]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [13]),
        .I4(\rgf/rgf_c1bus_0 [13]),
        .O(\sp[13]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[13]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/sptr/sp [13]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [13]),
        .O(\sp[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[14]_i_1 
       (.I0(\sp[14]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [14]),
        .I4(\rgf/rgf_c1bus_0 [14]),
        .O(\sp[14]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[14]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/sptr/sp [14]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [14]),
        .O(\sp[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[15]_i_1 
       (.I0(\sp[15]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [15]),
        .I4(\rgf/rgf_c1bus_0 [15]),
        .O(\sp[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00FFFF0200FFFFFF)) 
    \sp[15]_i_10 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [1]),
        .O(\sp[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h7E7EFFFFFFFFFF7E)) 
    \sp[15]_i_11 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [5]),
        .O(\sp[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF3E3EFFFF3E)) 
    \sp[15]_i_12 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .I5(\ctl0/stat [0]),
        .O(\sp[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \sp[15]_i_13 
       (.I0(\bcmd[1]_INST_0_i_3_n_0 ),
        .I1(brdy),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .I3(\bcmd[1]_INST_0_i_19_n_0 ),
        .I4(\sp[15]_i_21_n_0 ),
        .I5(\sp[15]_i_22_n_0 ),
        .O(ctl_sp_inc1));
  LUT5 #(
    .INIT(32'hF2F3DEDF)) 
    \sp[15]_i_14 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [6]),
        .O(\sp[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFF2FFF2FFF2FFFF)) 
    \sp[15]_i_15 
       (.I0(\fch/ir0 [10]),
        .I1(\sp[15]_i_23_n_0 ),
        .I2(\sp[15]_i_24_n_0 ),
        .I3(\stat[0]_i_10__0_n_0 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .O(\sp[15]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h44FFFFFC)) 
    \sp[15]_i_16 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .O(\sp[15]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00000004)) 
    \sp[15]_i_17 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .I1(brdy),
        .I2(\ctl1/stat [2]),
        .I3(\fch/ir1 [15]),
        .I4(\ctl1/stat [1]),
        .O(\sp[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFCFE6CFF7)) 
    \sp[15]_i_18 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [0]),
        .I5(\sp[15]_i_25_n_0 ),
        .O(\sp[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFF7FFFF00)) 
    \sp[15]_i_19 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [11]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [6]),
        .O(\sp[15]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[15]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/sptr/sp [15]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [15]),
        .O(\sp[15]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h1011)) 
    \sp[15]_i_20 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [12]),
        .I2(\ctl1/stat [0]),
        .I3(\pc0[15]_i_3_n_0 ),
        .O(\sp[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hE6E6FFFFFFFFFFE6)) 
    \sp[15]_i_21 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [11]),
        .I2(\ctl1/stat [0]),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [5]),
        .O(\sp[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF88FFFFF8)) 
    \sp[15]_i_22 
       (.I0(\ctl1/stat [0]),
        .I1(\bdatw[10]_INST_0_i_53_n_0 ),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [6]),
        .I5(\sp[15]_i_26_n_0 ),
        .O(\sp[15]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sp[15]_i_23 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [12]),
        .I2(\ctl0/stat [0]),
        .O(\sp[15]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h3E)) 
    \sp[15]_i_24 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .O(\sp[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7EFF7E7E7E7E)) 
    \sp[15]_i_25 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [8]),
        .I4(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I5(\fch/ir1 [4]),
        .O(\sp[15]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h7EFF7EFFFF7EFFFF)) 
    \sp[15]_i_26 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [5]),
        .O(\sp[15]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFF44445545)) 
    \sp[15]_i_5 
       (.I0(\sp[15]_i_8_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\pc0[15]_i_3_n_0 ),
        .I3(\ctl0/stat [0]),
        .I4(\fadr[15]_INST_0_i_11_n_0 ),
        .I5(ctl_sp_dec1),
        .O(\sp[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000001)) 
    \sp[15]_i_6 
       (.I0(\bcmd[1]_INST_0_i_14_n_0 ),
        .I1(\sp[15]_i_10_n_0 ),
        .I2(\sp[15]_i_11_n_0 ),
        .I3(\stat[0]_i_10__0_n_0 ),
        .I4(\sp[15]_i_12_n_0 ),
        .I5(ctl_sp_inc1),
        .O(\sp[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFFFFFFFFE)) 
    \sp[15]_i_8 
       (.I0(\sp[15]_i_14_n_0 ),
        .I1(\sp[15]_i_15_n_0 ),
        .I2(\sp[15]_i_16_n_0 ),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [10]),
        .O(\sp[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    \sp[15]_i_9 
       (.I0(\sp[15]_i_17_n_0 ),
        .I1(\sp[15]_i_18_n_0 ),
        .I2(\sp[15]_i_19_n_0 ),
        .I3(\bcmd[1]_INST_0_i_18_n_0 ),
        .I4(\fch/ir1 [10]),
        .I5(\sp[15]_i_20_n_0 ),
        .O(ctl_sp_dec1));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[1]_i_1 
       (.I0(\sp[1]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [1]),
        .I4(\rgf/rgf_c1bus_0 [1]),
        .O(\sp[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[1]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/sptr/sp [1]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [1]),
        .O(\sp[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[2]_i_1 
       (.I0(\sp[2]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .O(\sp[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[2]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/sptr/sp [2]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [2]),
        .O(\sp[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[3]_i_1 
       (.I0(\sp[3]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\rgf/rgf_c1bus_0 [3]),
        .O(\sp[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[3]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/sptr/sp [3]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [3]),
        .O(\sp[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[4]_i_1 
       (.I0(\sp[4]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [4]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .O(\sp[4]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[4]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/sptr/sp [4]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [4]),
        .O(\sp[4]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[5]_i_1 
       (.I0(\sp[5]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [5]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .O(\sp[5]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[5]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/sptr/sp [5]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [5]),
        .O(\sp[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[6]_i_1 
       (.I0(\sp[6]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [6]),
        .I4(\rgf/rgf_c1bus_0 [6]),
        .O(\sp[6]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[6]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/sptr/sp [6]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [6]),
        .O(\sp[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[7]_i_1 
       (.I0(\sp[7]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [7]),
        .I4(\rgf/rgf_c1bus_0 [7]),
        .O(\sp[7]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[7]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/sptr/sp [7]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [7]),
        .O(\sp[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[8]_i_1 
       (.I0(\sp[8]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [8]),
        .I4(\rgf/rgf_c1bus_0 [8]),
        .O(\sp[8]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[8]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/sptr/sp [8]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [8]),
        .O(\sp[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[9]_i_1 
       (.I0(\sp[9]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [9]),
        .I4(\rgf/rgf_c1bus_0 [9]),
        .O(\sp[9]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[9]_i_2 
       (.I0(\sp[15]_i_5_n_0 ),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/sptr/sp [9]),
        .I3(\sp[15]_i_6_n_0 ),
        .I4(\rgf/sptr/data2 [9]),
        .O(\sp[9]_i_2_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [11:8]),
        .S(\rgf/sptr/sp [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_7 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_7_n_1 ,\sp_reg[15]_i_7_n_2 ,\sp_reg[15]_i_7_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [15:12]),
        .S(\rgf/sptr/sp [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\badr[0]_INST_0_i_29_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [7:4]),
        .S(\rgf/sptr/sp [7:4]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[0]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [0]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[0]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [0]),
        .O(\rgf/rgf_c1bus_0 [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[0]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [0]),
        .O(\rgf/rgf_c0bus_0 [0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[10]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [10]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[10]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [10]),
        .O(\rgf/rgf_c1bus_0 [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[10]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [10]),
        .O(\rgf/rgf_c0bus_0 [10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[11]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [11]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in [11]));
  LUT6 #(
    .INIT(64'h444E000E000A000E)) 
    \sr[11]_i_10 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(\sr[11]_i_11_n_0 ),
        .I3(\ctl1/stat [2]),
        .I4(\rgf/rctl/rgf_selc1_stat ),
        .I5(\rgf/rctl/rgf_selc1_wb [0]),
        .O(\rgf/rctl/rgf_selc1 [0]));
  LUT6 #(
    .INIT(64'h00000000555555FD)) 
    \sr[11]_i_11 
       (.I0(\rgf_selc1_wb[0]_i_5_n_0 ),
        .I1(\sr[11]_i_12_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I3(\sr[11]_i_13_n_0 ),
        .I4(\sr[11]_i_14_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_2_n_0 ),
        .O(\sr[11]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \sr[11]_i_12 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [10]),
        .O(\sr[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF44440400)) 
    \sr[11]_i_13 
       (.I0(\rgf_selc1_wb[0]_i_18_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I2(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I3(\stat[0]_i_7__0_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_15_n_0 ),
        .I5(\sr[11]_i_15_n_0 ),
        .O(\sr[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0040444400401151)) 
    \sr[11]_i_14 
       (.I0(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\stat[0]_i_7__0_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\fch/ir1 [8]),
        .O(\sr[11]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[11]_i_15 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [1]),
        .O(\sr[11]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \sr[11]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(rst_n),
        .O(\sr[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[11]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [11]),
        .O(\rgf/rgf_c1bus_0 [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_4 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[11]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [11]),
        .O(\rgf/rgf_c0bus_0 [11]));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[11]_i_5 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\sr[15]_i_4_n_0 ),
        .I2(ctl_sr_ldie1),
        .I3(\sr[15]_i_6_n_0 ),
        .O(\sr[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_6 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(ctl_selc1_rn[2]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_rn_wb [2]),
        .O(\rgf/rctl/rgf_selc1_rn [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_7 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(ctl_selc1_rn[0]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_rn_wb [0]),
        .O(\rgf/rctl/rgf_selc1_rn [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_8 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(\rgf_selc1_rn_wb[1]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_rn_wb [1]),
        .O(\rgf/rctl/rgf_selc1_rn [1]));
  LUT6 #(
    .INIT(64'hAAFFAAFFBABFFFFF)) 
    \sr[11]_i_9 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1_wb [1]),
        .I2(\rgf/rctl/rgf_selc1_stat ),
        .I3(ctl_selc1),
        .I4(fch_term),
        .I5(fch_wrbufn1),
        .O(\sr[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFE00FE00FE00)) 
    \sr[12]_i_1 
       (.I0(ctl_sr_ldie0),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr[13]_i_4_n_0 ),
        .I3(cpuid[0]),
        .I4(\rgf/sreg/sr [12]),
        .I5(\sr[15]_i_2_n_0 ),
        .O(\rgf/sreg/p_0_in [12]));
  LUT6 #(
    .INIT(64'hFFFFFE00FE00FE00)) 
    \sr[13]_i_1 
       (.I0(ctl_sr_ldie0),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr[13]_i_4_n_0 ),
        .I3(cpuid[1]),
        .I4(\rgf/sreg/sr [13]),
        .I5(\sr[15]_i_2_n_0 ),
        .O(\rgf/sreg/p_0_in [13]));
  LUT4 #(
    .INIT(16'h0008)) 
    \sr[13]_i_10 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFF51BB0000)) 
    \sr[13]_i_11 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [15]),
        .I5(\sr[13]_i_12_n_0 ),
        .O(\sr[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000E222)) 
    \sr[13]_i_12 
       (.I0(\sr[13]_i_13_n_0 ),
        .I1(\sr[13]_i_14_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\sr[13]_i_15_n_0 ),
        .I4(\fch/ir0 [15]),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\sr[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AA040004)) 
    \sr[13]_i_13 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [6]),
        .I2(\bcmd[1]_INST_0_i_11_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [10]),
        .I5(\sr[13]_i_16_n_0 ),
        .O(\sr[13]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h37)) 
    \sr[13]_i_14 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .O(\sr[13]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h37)) 
    \sr[13]_i_15 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .O(\sr[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hC0BFFFFFC0FFFFC0)) 
    \sr[13]_i_16 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [4]),
        .O(\sr[13]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \sr[13]_i_2 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\sr[13]_i_5_n_0 ),
        .I3(\sr[13]_i_6_n_0 ),
        .I4(\sr[13]_i_7_n_0 ),
        .I5(\sr[13]_i_8_n_0 ),
        .O(ctl_sr_ldie0));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[13]_i_3 
       (.I0(ctl_sr_upd0),
        .I1(\rgf/c0bus_sel_cr [5]),
        .O(\sr[13]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_4 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\sr[15]_i_6_n_0 ),
        .I2(ctl_sr_ldie1),
        .I3(\sr[15]_i_4_n_0 ),
        .O(\sr[13]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_5 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .O(\sr[13]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_6 
       (.I0(\fch/ir0 [9]),
        .I1(\ctl0/stat [1]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [1]),
        .O(\sr[13]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[13]_i_7 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [3]),
        .O(\sr[13]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBF)) 
    \sr[13]_i_8 
       (.I0(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I1(\fch/ir0 [0]),
        .I2(brdy),
        .I3(\ctl0/stat [2]),
        .I4(\fch/ir0 [11]),
        .O(\sr[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    \sr[13]_i_9 
       (.I0(\sr[13]_i_11_n_0 ),
        .I1(\ctl0/stat [0]),
        .I2(\ctl0/stat [1]),
        .I3(\ctl0/stat [2]),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [15]),
        .O(ctl_sr_upd0));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[14]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [14]),
        .O(\rgf/sreg/p_0_in [14]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[15]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [15]),
        .O(\rgf/sreg/p_0_in [15]));
  LUT4 #(
    .INIT(16'h00FD)) 
    \sr[15]_i_2 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\sr[15]_i_4_n_0 ),
        .I2(ctl_sr_ldie1),
        .I3(\sr[15]_i_6_n_0 ),
        .O(\sr[15]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \sr[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [0]));
  LUT5 #(
    .INIT(32'hABAAAAAA)) 
    \sr[15]_i_4 
       (.I0(ctl_sr_upd1),
        .I1(\sr[11]_i_9_n_0 ),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\sr[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \sr[15]_i_5 
       (.I0(\sr[15]_i_7_n_0 ),
        .I1(\sr[15]_i_8_n_0 ),
        .I2(\bdatw[9]_INST_0_i_20_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I4(\bcmd[1]_INST_0_i_3_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_33_n_0 ),
        .O(ctl_sr_ldie1));
  LUT5 #(
    .INIT(32'h0001FFFF)) 
    \sr[15]_i_6 
       (.I0(\sr[11]_i_9_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(rst_n),
        .O(\sr[15]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \sr[15]_i_7 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .I1(brdy),
        .I2(\fch/ir1 [0]),
        .O(\sr[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[15]_i_8 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [3]),
        .O(\sr[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[1]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [1]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[1]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [1]),
        .O(\rgf/rgf_c1bus_0 [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[1]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [1]),
        .O(\rgf/rgf_c0bus_0 [1]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[2]_i_1 
       (.I0(\sr[2]_i_2_n_0 ),
        .I1(\sr[11]_i_2_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\sr[11]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in [2]));
  LUT5 #(
    .INIT(32'h8888F888)) 
    \sr[2]_i_2 
       (.I0(\rgf/sreg/sr [2]),
        .I1(\sr[3]_i_5_n_0 ),
        .I2(\sr[3]_i_6_n_0 ),
        .I3(fch_irq_lev[0]),
        .I4(\sr[15]_i_4_n_0 ),
        .O(\sr[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[2]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [2]),
        .O(\rgf/rgf_c1bus_0 [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[2]_i_4 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[2]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [2]),
        .O(\rgf/rgf_c0bus_0 [2]));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[3]_i_1 
       (.I0(\sr[3]_i_2_n_0 ),
        .I1(\sr[11]_i_2_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\sr[11]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in [3]));
  LUT5 #(
    .INIT(32'h8888F888)) 
    \sr[3]_i_2 
       (.I0(\rgf/sreg/sr [3]),
        .I1(\sr[3]_i_5_n_0 ),
        .I2(\sr[3]_i_6_n_0 ),
        .I3(fch_irq_lev[1]),
        .I4(\sr[15]_i_4_n_0 ),
        .O(\sr[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[3]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[3]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [3]),
        .O(\rgf/rgf_c1bus_0 [3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[3]_i_4 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[3]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [3]),
        .O(\rgf/rgf_c0bus_0 [3]));
  LUT6 #(
    .INIT(64'h0000FFFF0000000B)) 
    \sr[3]_i_5 
       (.I0(\sr[13]_i_3_n_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\rgf/c0bus_sel_cr [0]),
        .I3(ctl_sr_ldie1),
        .I4(\sr[15]_i_6_n_0 ),
        .I5(\sr[15]_i_4_n_0 ),
        .O(\sr[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00FF0004)) 
    \sr[3]_i_6 
       (.I0(\sr[13]_i_3_n_0 ),
        .I1(ctl_sr_ldie0),
        .I2(\rgf/c0bus_sel_cr [0]),
        .I3(\sr[15]_i_6_n_0 ),
        .I4(ctl_sr_ldie1),
        .O(\sr[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \sr[4]_i_1 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr[4]_i_3_n_0 ),
        .I2(\sr[4]_i_4_n_0 ),
        .I3(\sr[4]_i_5_n_0 ),
        .I4(alu_sr_flag1),
        .I5(\sr[4]_i_7_n_0 ),
        .O(\rgf/sreg/p_0_in [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_10 
       (.I0(\rgf_c0bus_wb[11]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .I4(\sr[4]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .O(\sr[4]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_11 
       (.I0(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .O(\sr[4]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_12 
       (.I0(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \sr[4]_i_13 
       (.I0(\sr[4]_i_26_n_0 ),
        .I1(\sr[4]_i_27_n_0 ),
        .I2(\sr[4]_i_28_n_0 ),
        .I3(\sr[4]_i_29_n_0 ),
        .I4(\sr[4]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .O(\sr[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_14 
       (.I0(\rgf_c1bus_wb[13]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_2_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .O(\sr[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDFFCF)) 
    \sr[4]_i_15 
       (.I0(\rgf_c1bus_wb[6]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_16 
       (.I0(\rgf_c1bus_wb[11]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .O(\sr[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \sr[4]_i_17 
       (.I0(\sr[4]_i_31_n_0 ),
        .I1(\sr[4]_i_32_n_0 ),
        .I2(\sr[4]_i_33_n_0 ),
        .I3(\sr[4]_i_34_n_0 ),
        .I4(\sr[4]_i_35_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_2_n_0 ),
        .O(\sr[4]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hAAABAAAA)) 
    \sr[4]_i_18 
       (.I0(\sr[4]_i_36_n_0 ),
        .I1(\sr[4]_i_37_n_0 ),
        .I2(\sr[4]_i_38_n_0 ),
        .I3(\sr[4]_i_39_n_0 ),
        .I4(\sr[4]_i_40_n_0 ),
        .O(\sr[4]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE000000)) 
    \sr[4]_i_19 
       (.I0(\sr[4]_i_41_n_0 ),
        .I1(\sr[4]_i_42_n_0 ),
        .I2(\sr[4]_i_43_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [15]),
        .O(ctl_sr_upd1));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\rgf/sreg/sr [4]),
        .O(\sr[4]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_20 
       (.I0(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[8]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb_reg[9]_i_3_n_0 ),
        .O(\sr[4]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_21 
       (.I0(\rgf_c0bus_wb_reg[0]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .O(\sr[4]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_22 
       (.I0(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb_reg[10]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .O(\sr[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \sr[4]_i_23 
       (.I0(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_8_n_0 ),
        .I2(\sr[4]_i_44_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .I5(\sr[4]_i_45_n_0 ),
        .O(\sr[4]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF07)) 
    \sr[4]_i_24 
       (.I0(tout__1_carry_i_12__0_n_0),
        .I1(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I2(\sr[4]_i_46_n_0 ),
        .I3(\rgf/sreg/sr [4]),
        .I4(\sr[4]_i_47_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .O(\sr[4]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h54FF54FFFFFF54FF)) 
    \sr[4]_i_25 
       (.I0(\sr[4]_i_48_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\sr[4]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I4(\sr[4]_i_50_n_0 ),
        .I5(\sr[4]_i_51_n_0 ),
        .O(\sr[4]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAAAA)) 
    \sr[4]_i_26 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_8_n_0 ),
        .I2(\bdatw[11]_INST_0_i_16_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .I5(\sr[4]_i_52_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hABABABABABABABAA)) 
    \sr[4]_i_27 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\sr[4]_i_53_n_0 ),
        .I2(\sr[4]_i_54_n_0 ),
        .I3(\sr[4]_i_55_n_0 ),
        .I4(\sr[4]_i_56_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\sr[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEFAAAA)) 
    \sr[4]_i_28 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\sr[4]_i_57_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .I4(\sr[4]_i_58_n_0 ),
        .I5(\sr[4]_i_59_n_0 ),
        .O(\sr[4]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEAAAEF)) 
    \sr[4]_i_29 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\sr[4]_i_60_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_6_n_0 ),
        .O(\sr[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[4]_i_3 
       (.I0(\sr[7]_i_3_n_0 ),
        .I1(\rgf/rctl/rgf_c1bus_wb [4]),
        .I2(\rgf/rctl/rgf_selc1_stat ),
        .I3(c1bus[4]),
        .I4(fch_term),
        .I5(fch_wrbufn1),
        .O(\sr[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBABBBABBBABA)) 
    \sr[4]_i_30 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .I2(\sr[4]_i_61_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I5(\sr[4]_i_62_n_0 ),
        .O(\sr[4]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBABABBBABBBABBBA)) 
    \sr[4]_i_31 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\sr[4]_i_63_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .O(\sr[4]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFCFCCCCCCCC)) 
    \sr[4]_i_32 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\sr[4]_i_64_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_10_n_0 ),
        .O(\sr[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hABABABABABABABAA)) 
    \sr[4]_i_33 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_11_n_0 ),
        .I2(\sr[4]_i_65_n_0 ),
        .I3(\sr[4]_i_66_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_15_n_0 ),
        .I5(\sr[4]_i_67_n_0 ),
        .O(\sr[4]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_34 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\sr[4]_i_68_n_0 ),
        .I2(\sr[4]_i_69_n_0 ),
        .O(\sr[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBABABBBA)) 
    \sr[4]_i_35 
       (.I0(\bdatw[12]_INST_0_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .I3(\sr[4]_i_70_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I5(\sr[4]_i_71_n_0 ),
        .O(\sr[4]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055551150)) 
    \sr[4]_i_36 
       (.I0(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I1(tout__1_carry_i_9__0_n_0),
        .I2(tout__1_carry_i_11__0_n_0),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\rgf/sreg/sr [4]),
        .I5(\sr[4]_i_72_n_0 ),
        .O(\sr[4]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_37 
       (.I0(\rgf_c1bus_wb[1]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .O(\sr[4]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_38 
       (.I0(\rgf_c1bus_wb[5]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_2_n_0 ),
        .I4(\sr[4]_i_73_n_0 ),
        .O(\sr[4]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_39 
       (.I0(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .O(\sr[4]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h88888888888888A8)) 
    \sr[4]_i_4 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr[4]_i_8_n_0 ),
        .I2(\sr[4]_i_9_n_0 ),
        .I3(\sr[4]_i_10_n_0 ),
        .I4(\sr[4]_i_11_n_0 ),
        .I5(\sr[4]_i_12_n_0 ),
        .O(\sr[4]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[4]_i_40 
       (.I0(\rgf_c1bus_wb_reg[0]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .O(\sr[4]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'h0FD50000)) 
    \sr[4]_i_41 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [15]),
        .O(\sr[4]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h755F755F557F555F)) 
    \sr[4]_i_42 
       (.I0(\fch/ir1 [8]),
        .I1(\sr[4]_i_74_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [11]),
        .O(\sr[4]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABABFFFBBBBB)) 
    \sr[4]_i_43 
       (.I0(\sr[4]_i_75_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(\sr[4]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'h80288088)) 
    \sr[4]_i_44 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\sr[4]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \sr[4]_i_45 
       (.I0(\sr[4]_i_76_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_45_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \sr[4]_i_46 
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .O(\sr[4]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_47 
       (.I0(\sr[4]_i_77_n_0 ),
        .I1(\alu0/art/add/tout__1_carry__2_n_6 ),
        .I2(\alu0/art/add/tout__1_carry__2_n_5 ),
        .I3(\alu0/art/add/tout__1_carry__2_n_7 ),
        .I4(\alu0/art/p_0_in ),
        .I5(\sr[4]_i_78_n_0 ),
        .O(\sr[4]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7020FFFF)) 
    \sr[4]_i_48 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\sr[4]_i_79_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I5(\sr[5]_i_12_n_0 ),
        .O(\sr[4]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hAA20AAAAAA20AA20)) 
    \sr[4]_i_49 
       (.I0(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .O(\sr[4]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[4]_i_5 
       (.I0(\sr[5]_i_5_n_0 ),
        .I1(\rgf/rctl/rgf_c0bus_wb [4]),
        .I2(\rgf/rctl/rgf_selc0_stat ),
        .I3(c0bus[4]),
        .I4(fch_term),
        .I5(fch_wrbufn0),
        .O(\sr[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB800B8FF)) 
    \sr[4]_i_50 
       (.I0(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0E000E000E000000)) 
    \sr[4]_i_51 
       (.I0(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .I2(\sr[4]_i_80_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_23_n_0 ),
        .I5(\sr[4]_i_81_n_0 ),
        .O(\sr[4]_i_51_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_52 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_6_n_0 ),
        .O(\sr[4]_i_52_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \sr[4]_i_53 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\sr[4]_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_54 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0C440C440C000CCC)) 
    \sr[4]_i_55 
       (.I0(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\sr[4]_i_55_n_0 ));
  LUT4 #(
    .INIT(16'h028A)) 
    \sr[4]_i_56 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .O(\sr[4]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \sr[4]_i_57 
       (.I0(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\sr[4]_i_82_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_57_n_0 ));
  LUT5 #(
    .INIT(32'h00400545)) 
    \sr[4]_i_58 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .O(\sr[4]_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hBABFAAAA)) 
    \sr[4]_i_59 
       (.I0(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000010)) 
    \sr[4]_i_6 
       (.I0(\sr[4]_i_13_n_0 ),
        .I1(\sr[4]_i_14_n_0 ),
        .I2(\sr[4]_i_15_n_0 ),
        .I3(\sr[4]_i_16_n_0 ),
        .I4(\sr[4]_i_17_n_0 ),
        .I5(\sr[4]_i_18_n_0 ),
        .O(alu_sr_flag1));
  LUT5 #(
    .INIT(32'h0400FFFF)) 
    \sr[4]_i_60 
       (.I0(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_60_n_0 ));
  LUT4 #(
    .INIT(16'h028A)) 
    \sr[4]_i_61 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .O(\sr[4]_i_61_n_0 ));
  LUT4 #(
    .INIT(16'hA202)) 
    \sr[4]_i_62 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .O(\sr[4]_i_62_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[4]_i_63 
       (.I0(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I3(\bdatw[11]_INST_0_i_16_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_63_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_64 
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .O(\sr[4]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \sr[4]_i_65 
       (.I0(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I1(a1bus_0[9]),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .O(\sr[4]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCEEECCCCCCCC)) 
    \sr[4]_i_66 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(\sr[4]_i_66_n_0 ));
  LUT5 #(
    .INIT(32'h00022202)) 
    \sr[4]_i_67 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .O(\sr[4]_i_67_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[4]_i_68 
       (.I0(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\sr[4]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBABABBBABAB)) 
    \sr[4]_i_69 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .O(\sr[4]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFF70000)) 
    \sr[4]_i_7 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(ctl_sr_upd1),
        .I5(\sr[15]_i_6_n_0 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h4)) 
    \sr[4]_i_70 
       (.I0(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .O(\sr[4]_i_70_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[4]_i_71 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .O(\sr[4]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_72 
       (.I0(\sr[4]_i_83_n_0 ),
        .I1(\alu1/art/add/tout__1_carry_n_4 ),
        .I2(\alu1/art/add/tout__1_carry__2_n_5 ),
        .I3(\alu1/art/add/tout__1_carry__1_n_4 ),
        .I4(\alu1/art/add/tout__1_carry__2_n_6 ),
        .I5(\sr[4]_i_84_n_0 ),
        .O(\sr[4]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFEAFF00FFEAFF11)) 
    \sr[4]_i_73 
       (.I0(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_25_n_0 ),
        .I3(\sr[4]_i_85_n_0 ),
        .I4(tout__1_carry_i_12_n_0),
        .I5(\ctl1/stat [2]),
        .O(\sr[4]_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hFFBF767676767676)) 
    \sr[4]_i_74 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [5]),
        .O(\sr[4]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \sr[4]_i_75 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [12]),
        .O(\sr[4]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0A05FFFFFEC00)) 
    \sr[4]_i_76 
       (.I0(\ccmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .I2(\ccmd[2]_INST_0_i_8_n_0 ),
        .I3(\ccmd[3]_INST_0_i_1_n_0 ),
        .I4(\ctl0/stat [2]),
        .I5(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_76_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_77 
       (.I0(\alu0/art/add/tout__1_carry__1_n_7 ),
        .I1(\alu0/art/add/tout__1_carry__1_n_6 ),
        .I2(\alu0/art/add/tout__1_carry__1_n_5 ),
        .I3(\alu0/art/add/tout__1_carry__1_n_4 ),
        .O(\sr[4]_i_77_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_78 
       (.I0(\alu0/art/add/tout__1_carry__0_n_4 ),
        .I1(\alu0/art/add/tout__1_carry__0_n_5 ),
        .I2(\alu0/art/add/tout__1_carry__0_n_6 ),
        .I3(\alu0/art/add/tout__1_carry__0_n_7 ),
        .I4(\sr[4]_i_86_n_0 ),
        .O(\sr[4]_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h000FFF0F33AA33AA)) 
    \sr[4]_i_79 
       (.I0(\rgf_c0bus_wb[15]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\sr[4]_i_79_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0100)) 
    \sr[4]_i_8 
       (.I0(\sr[4]_i_20_n_0 ),
        .I1(\sr[4]_i_21_n_0 ),
        .I2(\sr[4]_i_22_n_0 ),
        .I3(\sr[4]_i_23_n_0 ),
        .I4(\sr[4]_i_24_n_0 ),
        .O(\sr[4]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \sr[4]_i_80 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I2(a0bus_0[0]),
        .I3(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .O(\sr[4]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h30303F3F505F505F)) 
    \sr[4]_i_81 
       (.I0(\rgf_c0bus_wb[15]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_40_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\sr[4]_i_81_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_82 
       (.I0(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I1(a1bus_0[15]),
        .O(\sr[4]_i_82_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_83 
       (.I0(\alu1/art/add/tout__1_carry_n_6 ),
        .I1(\alu1/art/add/tout__1_carry_n_5 ),
        .I2(\alu1/art/add/tout__1_carry__0_n_7 ),
        .I3(\alu1/art/add/tout__1_carry__0_n_6 ),
        .O(\sr[4]_i_83_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_84 
       (.I0(\alu1/art/add/tout__1_carry__1_n_7 ),
        .I1(\alu1/art/add/tout__1_carry__0_n_5 ),
        .I2(\alu1/art/p_0_in ),
        .I3(\alu1/art/add/tout__1_carry__1_n_5 ),
        .I4(\sr[4]_i_87_n_0 ),
        .O(\sr[4]_i_84_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_85 
       (.I0(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_22_n_0 ),
        .O(\sr[4]_i_85_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_86 
       (.I0(\alu0/art/add/tout__1_carry_n_6 ),
        .I1(\alu0/art/add/tout__1_carry_n_5 ),
        .I2(\alu0/art/add/tout__1_carry_n_7 ),
        .I3(\alu0/art/add/tout__1_carry_n_4 ),
        .O(\sr[4]_i_86_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_87 
       (.I0(\alu1/art/add/tout__1_carry__0_n_4 ),
        .I1(\alu1/art/add/tout__1_carry__2_n_7 ),
        .I2(\alu1/art/add/tout__1_carry_n_7 ),
        .I3(\alu1/art/add/tout__1_carry__1_n_6 ),
        .O(\sr[4]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000BBBF)) 
    \sr[4]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .O(\sr[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \sr[5]_i_1 
       (.I0(\sr[5]_i_2_n_0 ),
        .I1(\sr[5]_i_3_n_0 ),
        .I2(\sr[5]_i_4_n_0 ),
        .I3(\sr[5]_i_5_n_0 ),
        .I4(\rgf/rgf_c0bus_0 [5]),
        .I5(\sr[5]_i_7_n_0 ),
        .O(\rgf/sreg/p_0_in [5]));
  LUT5 #(
    .INIT(32'h00090600)) 
    \sr[5]_i_10 
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[15]_INST_0_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I3(\alu1/art/p_0_in ),
        .I4(a1bus_0[15]),
        .O(\sr[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFBAAAAAAFBFBFBFB)) 
    \sr[5]_i_11 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(a0bus_0[14]),
        .I5(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .O(\sr[5]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hD0)) 
    \sr[5]_i_12 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_30_n_0 ),
        .O(\sr[5]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[5]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\rgf/sreg/sr [5]),
        .O(\sr[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[5]_i_3 
       (.I0(\sr[7]_i_3_n_0 ),
        .I1(\rgf/rctl/rgf_c1bus_wb [5]),
        .I2(\rgf/rctl/rgf_selc1_stat ),
        .I3(c1bus[5]),
        .I4(fch_term),
        .I5(fch_wrbufn1),
        .O(\sr[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA20000020)) 
    \sr[5]_i_4 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_7_n_0 ),
        .I4(\sr[5]_i_8_n_0 ),
        .I5(\sr[5]_i_9_n_0 ),
        .O(\sr[5]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00001110)) 
    \sr[5]_i_5 
       (.I0(ctl_sr_ldie1),
        .I1(\sr[15]_i_4_n_0 ),
        .I2(\rgf/c0bus_sel_cr [0]),
        .I3(\rgf/c0bus_sel_cr [5]),
        .I4(\sr[15]_i_6_n_0 ),
        .O(\sr[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[5]_i_6 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[5]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [5]),
        .O(\rgf/rgf_c0bus_0 [5]));
  LUT6 #(
    .INIT(64'hAAAAAAAA00002800)) 
    \sr[5]_i_7 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(\sr[6]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I5(\sr[5]_i_10_n_0 ),
        .O(\sr[5]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \sr[5]_i_8 
       (.I0(\sr[5]_i_11_n_0 ),
        .I1(\sr[5]_i_12_n_0 ),
        .I2(\sr[6]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .O(\sr[5]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00060900)) 
    \sr[5]_i_9 
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[15]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I3(\alu0/art/p_0_in ),
        .I4(a0bus_0[15]),
        .O(\sr[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \sr[6]_i_1 
       (.I0(\sr[6]_i_2_n_0 ),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\sr[6]_i_4_n_0 ),
        .I4(\sr[6]_i_5_n_0 ),
        .I5(\sr[6]_i_6_n_0 ),
        .O(\rgf/sreg/p_0_in [6]));
  LUT6 #(
    .INIT(64'h55CF550055C05500)) 
    \sr[6]_i_10 
       (.I0(\sr[6]_i_17_n_0 ),
        .I1(\sr[6]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .O(\sr[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAFEAE)) 
    \sr[6]_i_11 
       (.I0(\sr[6]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_17_n_0 ),
        .O(\sr[6]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[6]_i_12 
       (.I0(\rgf_c0bus_wb[15]_i_31_n_0 ),
        .I1(a0bus_0[15]),
        .O(\sr[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h1FFF11BB1FFF1FFF)) 
    \sr[6]_i_13 
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I3(\ccmd[2]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .O(\sr[6]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_14 
       (.I0(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .O(\sr[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAA0AA8800000000)) 
    \sr[6]_i_15 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I2(\sr[6]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I5(\sr[6]_i_21_n_0 ),
        .O(\sr[6]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0003005300F300F3)) 
    \sr[6]_i_16 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .I3(\bdatw[12]_INST_0_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .I5(\sr[6]_i_22_n_0 ),
        .O(\sr[6]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \sr[6]_i_17 
       (.I0(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .O(\sr[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00F0DDFD00F000F0)) 
    \sr[6]_i_18 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .O(\sr[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFF400F4)) 
    \sr[6]_i_19 
       (.I0(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I2(\sr[6]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_33_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .O(\sr[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h3F3050503F3F5F5F)) 
    \sr[6]_i_20 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I4(\bdatw[8]_INST_0_i_14_n_0 ),
        .I5(a1bus_0[15]),
        .O(\sr[6]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[6]_i_21 
       (.I0(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .O(\sr[6]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h5555DF55FFFFDF55)) 
    \sr[6]_i_22 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .I3(\sr[6]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .O(\sr[6]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h3F002A0000002A00)) 
    \sr[6]_i_23 
       (.I0(\rgf_c0bus_wb[12]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_30_n_0 ),
        .O(\sr[6]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h30FF75FFFFFF75FF)) 
    \sr[6]_i_24 
       (.I0(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .O(\sr[6]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[6]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[6]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [6]),
        .O(\rgf/rgf_c1bus_0 [6]));
  LUT5 #(
    .INIT(32'h8A88888A)) 
    \sr[6]_i_4 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr[6]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I3(tout__1_carry_i_8__0_n_0),
        .I4(\alu0/art/add/tout ),
        .O(\sr[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[6]_i_5 
       (.I0(\sr[5]_i_5_n_0 ),
        .I1(\rgf/rctl/rgf_c0bus_wb [6]),
        .I2(\rgf/rctl/rgf_selc0_stat ),
        .I3(c0bus[6]),
        .I4(fch_term),
        .I5(fch_wrbufn0),
        .O(\sr[6]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA8A80)) 
    \sr[6]_i_6 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(tout__1_carry_i_10__0_n_0),
        .I2(\alu1/art/add/tout ),
        .I3(tout__1_carry_i_8_n_0),
        .I4(\sr[6]_i_8_n_0 ),
        .O(\sr[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022220FFF)) 
    \sr[6]_i_7 
       (.I0(\sr[6]_i_9_n_0 ),
        .I1(\sr[6]_i_10_n_0 ),
        .I2(\sr[6]_i_11_n_0 ),
        .I3(\sr[6]_i_12_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\sr[6]_i_13_n_0 ),
        .O(\sr[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000033BF)) 
    \sr[6]_i_8 
       (.I0(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(\sr[6]_i_15_n_0 ),
        .I4(\sr[6]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .O(\sr[6]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h47FF)) 
    \sr[6]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\sr[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \sr[7]_i_1 
       (.I0(\sr[7]_i_2_n_0 ),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\sr[7]_i_5_n_0 ),
        .I4(\sr[7]_i_6_n_0 ),
        .I5(\sr[7]_i_7_n_0 ),
        .O(\rgf/sreg/p_0_in [7]));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[7]_i_2 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(\rgf/sreg/sr [7]),
        .O(\sr[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00090000)) 
    \sr[7]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\sr[11]_i_9_n_0 ),
        .I4(rst_n),
        .O(\sr[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[7]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[7]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [7]),
        .O(\rgf/rgf_c1bus_0 [7]));
  LUT5 #(
    .INIT(32'hEEFE0000)) 
    \sr[7]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .I2(\alu0/art/p_0_in ),
        .I3(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I4(\sr[7]_i_9_n_0 ),
        .O(\sr[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAA00AA008A800000)) 
    \sr[7]_i_6 
       (.I0(\sr[5]_i_5_n_0 ),
        .I1(\rgf/rctl/rgf_c0bus_wb [7]),
        .I2(\rgf/rctl/rgf_selc0_stat ),
        .I3(c0bus[7]),
        .I4(fch_term),
        .I5(fch_wrbufn0),
        .O(\sr[7]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEEFE0000)) 
    \sr[7]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\alu1/art/p_0_in ),
        .I3(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I4(\sr[4]_i_7_n_0 ),
        .O(\sr[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055550001)) 
    \sr[7]_i_8 
       (.I0(\sr[15]_i_4_n_0 ),
        .I1(ctl_sr_upd0),
        .I2(\rgf/c0bus_sel_cr [5]),
        .I3(\rgf/c0bus_sel_cr [0]),
        .I4(ctl_sr_ldie1),
        .I5(\sr[15]_i_6_n_0 ),
        .O(\sr[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \sr[7]_i_9 
       (.I0(\rgf/c0bus_sel_cr [5]),
        .I1(ctl_sr_upd0),
        .I2(\sr[15]_i_4_n_0 ),
        .I3(ctl_sr_ldie1),
        .I4(\sr[15]_i_6_n_0 ),
        .I5(\rgf/c0bus_sel_cr [0]),
        .O(\sr[7]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[8]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf/sreg/p_0_in [8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \sr[9]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [9]),
        .I2(\sr[11]_i_2_n_0 ),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\sr[11]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[9]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [9]),
        .O(\rgf/rgf_c1bus_0 [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[9]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [9]),
        .O(\rgf/rgf_c0bus_0 [9]));
  LUT6 #(
    .INIT(64'h000000000000EAEE)) 
    \stat[0]_i_1 
       (.I0(\stat[0]_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_2_n_0 ),
        .I2(\stat[0]_i_3_n_0 ),
        .I3(\stat[0]_i_4_n_0 ),
        .I4(\stat[0]_i_5_n_0 ),
        .I5(\fch/ir0 [15]),
        .O(\ctl0/stat_nx [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000012)) 
    \stat[0]_i_10 
       (.I0(\stat[0]_i_22__0_n_0 ),
        .I1(\ctl0/stat [1]),
        .I2(\fch/ir0 [11]),
        .I3(\ctl0/stat [2]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [13]),
        .O(\stat[0]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \stat[0]_i_10__0 
       (.I0(\fch/ir0 [15]),
        .I1(\ctl0/stat [1]),
        .I2(\ctl0/stat [2]),
        .I3(brdy),
        .O(\stat[0]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'h01000001)) 
    \stat[0]_i_10__1 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\rgf/sreg/sr [5]),
        .O(\stat[0]_i_10__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFEEEE)) 
    \stat[0]_i_11 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(\fch/ir0 [14]),
        .I2(\ccmd[4]_INST_0_i_8_n_0 ),
        .I3(\ctl0/stat [2]),
        .I4(\fch/ir0 [13]),
        .I5(\stat[0]_i_24_n_0 ),
        .O(\stat[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF40FF40404040)) 
    \stat[0]_i_11__0 
       (.I0(\stat[0]_i_22_n_0 ),
        .I1(\stat[2]_i_5__0_n_0 ),
        .I2(\stat[0]_i_23__0_n_0 ),
        .I3(\stat[0]_i_24__0_n_0 ),
        .I4(\stat[0]_i_25__0_n_0 ),
        .I5(\stat[0]_i_26__0_n_0 ),
        .O(\stat[0]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF040404FF)) 
    \stat[0]_i_11__1 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [8]),
        .I3(\mem/bctl/fch_term_fl ),
        .I4(\mem/bctl/ctl/p_0_in [5]),
        .I5(\stat[0]_i_14__1_n_0 ),
        .O(\stat[0]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004400444)) 
    \stat[0]_i_12 
       (.I0(\fch/ir0 [4]),
        .I1(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I2(\fch/ir0 [0]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [1]),
        .I5(\ccmd[2]_INST_0_i_5_n_0 ),
        .O(\stat[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBBAABBAAFFAAF0AA)) 
    \stat[0]_i_12__0 
       (.I0(\stat[0]_i_27_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\rgf/ivec/iv [0]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [1]),
        .O(\stat[0]_i_12__0_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \stat[0]_i_12__1 
       (.I0(\fch/ir0 [12]),
        .I1(\ctl0/stat [1]),
        .I2(\fch/ir0 [13]),
        .O(\stat[0]_i_12__1_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFEFF0000)) 
    \stat[0]_i_13 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [6]),
        .I2(brdy),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [11]),
        .I5(\stat[0]_i_25_n_0 ),
        .O(\stat[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_13__0 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .O(\stat[0]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_13__1 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [6]),
        .O(\stat[0]_i_13__1_n_0 ));
  LUT6 #(
    .INIT(64'h0E0EEEEE0EFFEEEE)) 
    \stat[0]_i_14 
       (.I0(crdy),
        .I1(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\stat[0]_i_26_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\stat[0]_i_27__0_n_0 ),
        .O(\stat[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDD101C)) 
    \stat[0]_i_14__0 
       (.I0(\stat[0]_i_28__0_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .I5(\stat[0]_i_29_n_0 ),
        .O(\stat[0]_i_14__0_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[0]_i_14__1 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .O(\stat[0]_i_14__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF1F001F001F00)) 
    \stat[0]_i_15 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\stat[0]_i_28__0_n_0 ),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA88AA8AAA8)) 
    \stat[0]_i_15__0 
       (.I0(\ctl0/stat [0]),
        .I1(\stat[0]_i_28_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(brdy),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [5]),
        .O(\stat[0]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFB00000B0B0)) 
    \stat[0]_i_16 
       (.I0(\bcmd[0]_INST_0_i_26_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\stat[0]_i_29__0_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [10]),
        .I5(\stat[0]_i_30_n_0 ),
        .O(\stat[0]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[0]_i_16__0 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir1 [11]),
        .O(\stat[0]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'hA888A8888888A888)) 
    \stat[0]_i_17 
       (.I0(\fch/ir0 [10]),
        .I1(\stat[0]_i_31_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .I4(\stat[0]_i_32_n_0 ),
        .I5(\stat[0]_i_33_n_0 ),
        .O(\stat[0]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h01555555)) 
    \stat[0]_i_17__0 
       (.I0(\fch/fch_irq_req_fl ),
        .I1(\fch/ir0_id_fl [21]),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/rst_n_fl ),
        .I4(\ir0_id_fl[21]_i_2_n_0 ),
        .O(\stat[0]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h8000804000000000)) 
    \stat[0]_i_18 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\stat[0]_i_30__0_n_0 ),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [3]),
        .O(\stat[0]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_18__0 
       (.I0(\ctl0/stat [0]),
        .I1(\fch/ir0 [9]),
        .O(\stat[0]_i_18__0_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_19 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [11]),
        .I3(\ctl0/stat [2]),
        .O(\stat[0]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_19__0 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [9]),
        .O(\stat[0]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h000044444F444444)) 
    \stat[0]_i_1__0 
       (.I0(\stat[0]_i_2__1_n_0 ),
        .I1(\rgf/pcnt/pc [1]),
        .I2(\stat[2]_i_3__1_n_0 ),
        .I3(\fadr[15]_INST_0_i_4_n_0 ),
        .I4(\fch/stat [0]),
        .I5(\stat[0]_i_3__1_n_0 ),
        .O(\fch/fctl/stat_nx [0]));
  LUT6 #(
    .INIT(64'h000B0000FFFFFFFF)) 
    \stat[0]_i_1__1 
       (.I0(\stat[0]_i_2__2_n_0 ),
        .I1(\stat[0]_i_3__2_n_0 ),
        .I2(\stat[0]_i_4__0_n_0 ),
        .I3(\stat[0]_i_5__0_n_0 ),
        .I4(\stat[0]_i_6__0_n_0 ),
        .I5(\bcmd[2]_INST_0_i_1_n_0 ),
        .O(\mem/bctl/ctl/stat_nx [0]));
  LUT6 #(
    .INIT(64'h000000000000FF08)) 
    \stat[0]_i_1__2 
       (.I0(\stat[0]_i_2__0_n_0 ),
        .I1(\stat[0]_i_3__0_n_0 ),
        .I2(\stat[2]_i_3__0_n_0 ),
        .I3(\stat[0]_i_4__1_n_0 ),
        .I4(\stat[0]_i_5__1_n_0 ),
        .I5(\fch/ir1 [15]),
        .O(\ctl1/stat_nx [0]));
  LUT6 #(
    .INIT(64'h00000000FFFF08AA)) 
    \stat[0]_i_2 
       (.I0(\stat[0]_i_6__1_n_0 ),
        .I1(\stat[0]_i_7_n_0 ),
        .I2(\stat[0]_i_8_n_0 ),
        .I3(\stat[0]_i_9__0_n_0 ),
        .I4(\stat[0]_i_10_n_0 ),
        .I5(\stat[0]_i_11_n_0 ),
        .O(\stat[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_20 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [10]),
        .O(\stat[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_20__0 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [11]),
        .O(\stat[0]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBABBBABBBABABAB)) 
    \stat[0]_i_21 
       (.I0(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I1(\stat[0]_i_34__0_n_0 ),
        .I2(ctl_fetch0_fl_i_12_n_0),
        .I3(\ctl0/stat [2]),
        .I4(\ctl0/stat [1]),
        .I5(\fch/ir0 [1]),
        .O(\stat[0]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_21__0 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [5]),
        .O(\stat[0]_i_21__0_n_0 ));
  LUT6 #(
    .INIT(64'h556595A5596999A9)) 
    \stat[0]_i_22 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\rgf/sreg/sr [6]),
        .O(\stat[0]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_22__0 
       (.I0(\fch/ir0 [12]),
        .I1(\rgf/sreg/sr [4]),
        .O(\stat[0]_i_22__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000410151515151)) 
    \stat[0]_i_23 
       (.I0(\ctl0/stat [2]),
        .I1(\ctl0/stat [0]),
        .I2(brdy),
        .I3(\fch/ir0 [0]),
        .I4(\stat[0]_i_35_n_0 ),
        .I5(\stat[0]_i_36__0_n_0 ),
        .O(\stat[0]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_23__0 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [14]),
        .O(\stat[0]_i_23__0_n_0 ));
  LUT5 #(
    .INIT(32'h0A22A088)) 
    \stat[0]_i_24 
       (.I0(\fch/ir0 [13]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [11]),
        .O(\stat[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF8CBB)) 
    \stat[0]_i_24__0 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [2]),
        .I2(\rgf/sreg/sr [10]),
        .I3(\fch/ir1 [1]),
        .I4(\stat[0]_i_31__0_n_0 ),
        .I5(\stat[0]_i_32__0_n_0 ),
        .O(\stat[0]_i_24__0_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBB8BBBB)) 
    \stat[0]_i_25 
       (.I0(crdy),
        .I1(\ccmd[4]_INST_0_i_13_n_0 ),
        .I2(brdy),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [9]),
        .I5(\ccmd[4]_INST_0_i_16_n_0 ),
        .O(\stat[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000ABFEABFF)) 
    \stat[0]_i_25__0 
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [2]),
        .I3(\ctl1/stat [0]),
        .I4(\pc0[15]_i_3_n_0 ),
        .I5(\stat[0]_i_33__0_n_0 ),
        .O(\stat[0]_i_25__0_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \stat[0]_i_26 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(crdy),
        .I3(\fch/ir0 [8]),
        .O(\stat[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000D500D500D500)) 
    \stat[0]_i_26__0 
       (.I0(\fch/ir1 [12]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [11]),
        .I3(\stat[0]_i_34_n_0 ),
        .I4(\bdatw[15]_INST_0_i_42_n_0 ),
        .I5(\rgf/sreg/sr [10]),
        .O(\stat[0]_i_26__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \stat[0]_i_27 
       (.I0(\fch/ir1 [1]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [2]),
        .O(\stat[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0800080000000400)) 
    \stat[0]_i_27__0 
       (.I0(\fch/ir0 [5]),
        .I1(\badrx[15]_INST_0_i_4_n_0 ),
        .I2(brdy),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [6]),
        .O(\stat[0]_i_27__0_n_0 ));
  LUT5 #(
    .INIT(32'h7F3FFF3F)) 
    \stat[0]_i_28 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [10]),
        .O(\stat[0]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \stat[0]_i_28__0 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .I1(brdy),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [9]),
        .O(\stat[0]_i_28__0_n_0 ));
  LUT5 #(
    .INIT(32'hF2000000)) 
    \stat[0]_i_29 
       (.I0(brdy),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(\badr[15]_INST_0_i_215_n_0 ),
        .I3(\stat[0]_i_35__0_n_0 ),
        .I4(\fch/ir1 [11]),
        .O(\stat[0]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_29__0 
       (.I0(\ccmd[4]_INST_0_i_13_n_0 ),
        .I1(crdy),
        .O(\stat[0]_i_29__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55550030)) 
    \stat[0]_i_2__0 
       (.I0(\stat[0]_i_6_n_0 ),
        .I1(\stat[0]_i_7__0_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\stat[0]_i_8__0_n_0 ),
        .I4(\stat[0]_i_9__1_n_0 ),
        .I5(\stat[0]_i_10__1_n_0 ),
        .O(\stat[0]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_2__1 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\stat[1]_i_2__0_n_0 ),
        .O(\stat[0]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h1010101000000001)) 
    \stat[0]_i_2__2 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [11]),
        .O(\stat[0]_i_2__2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_3 
       (.I0(\stat[2]_i_9_n_0 ),
        .I1(\stat[2]_i_4_n_0 ),
        .O(\stat[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \stat[0]_i_30 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(brdy),
        .O(\stat[0]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \stat[0]_i_30__0 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [11]),
        .O(\stat[0]_i_30__0_n_0 ));
  LUT6 #(
    .INIT(64'h4F404F4F45404540)) 
    \stat[0]_i_31 
       (.I0(\rgf_selc0_wb[0]_i_14_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [11]),
        .I3(crdy),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\stat[0]_i_30_n_0 ),
        .O(\stat[0]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \stat[0]_i_31__0 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\stat[2]_i_5__0_n_0 ),
        .I5(\bdatw[11]_INST_0_i_27_n_0 ),
        .O(\stat[0]_i_31__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_32 
       (.I0(\fch/ir0 [9]),
        .I1(crdy),
        .O(\stat[0]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \stat[0]_i_32__0 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [10]),
        .O(\stat[0]_i_32__0_n_0 ));
  LUT6 #(
    .INIT(64'h8900010000000100)) 
    \stat[0]_i_33 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [4]),
        .I3(\stat[0]_i_37_n_0 ),
        .I4(\fch/ir0 [3]),
        .I5(brdy),
        .O(\stat[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4F4F4C4)) 
    \stat[0]_i_33__0 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\ctl1/stat [2]),
        .I3(\fch/ir1 [1]),
        .I4(\ctl1/stat [1]),
        .I5(\stat[0]_i_36_n_0 ),
        .O(\stat[0]_i_33__0_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_34 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .O(\stat[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000140000)) 
    \stat[0]_i_34__0 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\ctl0/stat [2]),
        .I4(\fch/ir0 [2]),
        .I5(\stat[0]_i_38_n_0 ),
        .O(\stat[0]_i_34__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF1)) 
    \stat[0]_i_35 
       (.I0(\ccmd[4]_INST_0_i_8_n_0 ),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [12]),
        .O(\stat[0]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h8000000080000088)) 
    \stat[0]_i_35__0 
       (.I0(\fch/ir1 [7]),
        .I1(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [4]),
        .O(\stat[0]_i_35__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[0]_i_36 
       (.I0(\badr[15]_INST_0_i_296_n_0 ),
        .I1(ctl_fetch1_fl_i_17_n_0),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [10]),
        .O(\stat[0]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFEF)) 
    \stat[0]_i_36__0 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [13]),
        .I2(\ctl0/stat [0]),
        .I3(\rgf/ivec/iv [0]),
        .O(\stat[0]_i_36__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_37 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [7]),
        .O(\stat[0]_i_37_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_38 
       (.I0(\ctl0/stat [1]),
        .I1(crdy),
        .O(\stat[0]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_3__0 
       (.I0(\fch/ir1 [14]),
        .I1(\ctl1/stat [2]),
        .O(\stat[0]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_3__1 
       (.I0(\fch/stat [1]),
        .I1(\fch/stat [2]),
        .O(\stat[0]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h77BF0000FFFFFFFF)) 
    \stat[0]_i_3__2 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\stat[0]_i_7__1_n_0 ),
        .I5(\stat[0]_i_8__1_n_0 ),
        .O(\stat[0]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'hEAAAEAAAEAAAEAFF)) 
    \stat[0]_i_4 
       (.I0(\stat[0]_i_12__1_n_0 ),
        .I1(\stat[0]_i_13_n_0 ),
        .I2(\stat[0]_i_14_n_0 ),
        .I3(\stat[0]_i_15__0_n_0 ),
        .I4(\stat[0]_i_16_n_0 ),
        .I5(\stat[0]_i_17_n_0 ),
        .O(\stat[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEFFFFFE)) 
    \stat[0]_i_4__0 
       (.I0(\stat[0]_i_9_n_0 ),
        .I1(\stat[0]_i_10__0_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [12]),
        .I5(\stat[0]_i_11__1_n_0 ),
        .O(\stat[0]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAA8288)) 
    \stat[0]_i_4__1 
       (.I0(\stat[0]_i_11__0_n_0 ),
        .I1(\ctl1/stat [0]),
        .I2(\bcmd[2]_INST_0_i_1_n_0 ),
        .I3(brdy),
        .I4(\ctl1/stat [2]),
        .I5(\stat[0]_i_12__0_n_0 ),
        .O(\stat[0]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000800000)) 
    \stat[0]_i_5 
       (.I0(\fch/ir0 [10]),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(\stat[0]_i_18__0_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\rgf/sreg/sr [11]),
        .I5(\fch/ir0 [11]),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFEEEEEFFEEEEEEEE)) 
    \stat[0]_i_5__0 
       (.I0(\stat[0]_i_12_n_0 ),
        .I1(\bcmd[1]_INST_0_i_11_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [10]),
        .I5(\stat[0]_i_13__1_n_0 ),
        .O(\stat[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000800080000)) 
    \stat[0]_i_5__1 
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(\stat[0]_i_13__0_n_0 ),
        .I2(\fch/ir1 [7]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [11]),
        .I5(\rgf/sreg/sr [11]),
        .O(\stat[0]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hA030AF3FAF3FA030)) 
    \stat[0]_i_6 
       (.I0(\stat[0]_i_14__0_n_0 ),
        .I1(\stat[0]_i_15_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [10]),
        .I4(\stat[0]_i_16__0_n_0 ),
        .I5(\rgf/sreg/sr [5]),
        .O(\stat[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hE0FFE0E0)) 
    \stat[0]_i_6__0 
       (.I0(\fch/fch_irq_req_fl ),
        .I1(\fch/ir0_id ),
        .I2(fch_memacc1),
        .I3(\mem/bctl/ctl/p_0_in [4]),
        .I4(\mem/bctl/ctl/p_0_in [5]),
        .O(\stat[0]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h7F0000007F7F7F7F)) 
    \stat[0]_i_6__1 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .I2(\rgf/sreg/sr [10]),
        .I3(\fch/ir0 [11]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\fch/ir0 [12]),
        .O(\stat[0]_i_6__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000005F1F1010)) 
    \stat[0]_i_7 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [1]),
        .I3(\rgf/sreg/sr [10]),
        .I4(crdy),
        .I5(\stat[0]_i_19_n_0 ),
        .O(\stat[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hA2220000A2228000)) 
    \stat[0]_i_7__0 
       (.I0(brdy),
        .I1(\mem/bctl/fch_term_fl ),
        .I2(\stat[0]_i_17__0_n_0 ),
        .I3(fch_memacc1),
        .I4(\mem/bctl/ctl/p_0_in [4]),
        .I5(\mem/bctl/ctl/p_0_in [5]),
        .O(\stat[0]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_7__1 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .O(\stat[0]_i_7__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBAB)) 
    \stat[0]_i_8 
       (.I0(\stat[0]_i_20_n_0 ),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [2]),
        .I3(\ctl0/stat [0]),
        .I4(\ctl0/stat [1]),
        .I5(\fch/ir0 [9]),
        .O(\stat[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h5550555555505515)) 
    \stat[0]_i_8__0 
       (.I0(\stat[0]_i_18_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [10]),
        .I3(\stat[0]_i_19__0_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .O(\stat[0]_i_8__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_8__1 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .O(\stat[0]_i_8__1_n_0 ));
  LUT6 #(
    .INIT(64'hAA5FFE5EFF5FFEFE)) 
    \stat[0]_i_9 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [12]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [11]),
        .O(\stat[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF54015400)) 
    \stat[0]_i_9__0 
       (.I0(\ctl0/stat [2]),
        .I1(\ctl0/stat [1]),
        .I2(\fch/ir0 [2]),
        .I3(\ctl0/stat [0]),
        .I4(\pc0[15]_i_3_n_0 ),
        .I5(\stat[0]_i_21_n_0 ),
        .O(\stat[0]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h80300030FFFFFFFF)) 
    \stat[0]_i_9__1 
       (.I0(ctl_fetch1_fl_i_11_n_0),
        .I1(\fch/ir1 [8]),
        .I2(\stat[0]_i_20__0_n_0 ),
        .I3(\stat[0]_i_7__0_n_0 ),
        .I4(\stat[0]_i_21__0_n_0 ),
        .I5(\ctl1/stat [0]),
        .O(\stat[0]_i_9__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000001111FF0F)) 
    \stat[1]_i_1 
       (.I0(\stat[1]_i_2_n_0 ),
        .I1(\ctl0/stat [2]),
        .I2(\stat[1]_i_3_n_0 ),
        .I3(\stat_reg[1]_i_4_n_0 ),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [15]),
        .O(\ctl0/stat_nx [1]));
  LUT6 #(
    .INIT(64'h00FF00FF822282A2)) 
    \stat[1]_i_10 
       (.I0(\stat[1]_i_18_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\stat[1]_i_19__0_n_0 ),
        .I3(\ctl0/stat [1]),
        .I4(\rgf/sreg/sr [10]),
        .I5(\fch/ir0 [11]),
        .O(\stat[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h1111111100101000)) 
    \stat[1]_i_10__0 
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [1]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [11]),
        .O(\stat[1]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFCFCFC0CC5757)) 
    \stat[1]_i_11 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [0]),
        .I3(\rgf/sreg/sr [10]),
        .I4(\fch/ir1 [2]),
        .I5(\ctl1/stat [2]),
        .O(\stat[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAAA2A)) 
    \stat[1]_i_11__0 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [11]),
        .I2(\rgf/sreg/sr [4]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [13]),
        .O(\stat[1]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \stat[1]_i_12 
       (.I0(\ctl0/stat [1]),
        .I1(\fch/ir0 [11]),
        .I2(\ctl0/stat [2]),
        .I3(\ctl0/stat [0]),
        .I4(\fch/ir0 [13]),
        .I5(\rgf/sreg/sr [6]),
        .O(\stat[1]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAAA2A)) 
    \stat[1]_i_12__0 
       (.I0(\fch/ir1 [12]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [11]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [13]),
        .O(\stat[1]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h4400000400440004)) 
    \stat[1]_i_13 
       (.I0(\ctl0/stat [2]),
        .I1(\ccmd[4]_INST_0_i_8_n_0 ),
        .I2(\rgf/sreg/sr [4]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [13]),
        .I5(\rgf/sreg/sr [7]),
        .O(\stat[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \stat[1]_i_13__0 
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [0]),
        .I2(\ctl1/stat [1]),
        .I3(\fch/ir1 [13]),
        .I4(\rgf/sreg/sr [6]),
        .I5(\fch/ir1 [11]),
        .O(\stat[1]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000084870000)) 
    \stat[1]_i_14 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [11]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\badr[15]_INST_0_i_144_n_0 ),
        .I5(\ctl1/stat [2]),
        .O(\stat[1]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_14__0 
       (.I0(\ctl0/stat [1]),
        .I1(\ctl0/stat [0]),
        .O(\stat[1]_i_14__0_n_0 ));
  LUT6 #(
    .INIT(64'h00C0500000000000)) 
    \stat[1]_i_15 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .I2(\stat[1]_i_20_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\ctl0/stat [0]),
        .I5(\stat[1]_i_21_n_0 ),
        .O(\stat[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[1]_i_15__0 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .O(\stat[1]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000C0500)) 
    \stat[1]_i_16 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [10]),
        .I2(\stat[1]_i_19_n_0 ),
        .I3(\fch/ir1 [9]),
        .I4(\ctl1/stat [0]),
        .I5(\stat[1]_i_20__0_n_0 ),
        .O(\stat[1]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00000024)) 
    \stat[1]_i_16__0 
       (.I0(\ctl0/stat [0]),
        .I1(\ctl0/stat [1]),
        .I2(brdy),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [9]),
        .O(\stat[1]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'h80808F8020202020)) 
    \stat[1]_i_17 
       (.I0(\stat[1]_i_22_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [9]),
        .I3(\stat[1]_i_23_n_0 ),
        .I4(\ctl0/stat [1]),
        .I5(\ctl0/stat [0]),
        .O(\stat[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000057555757)) 
    \stat[1]_i_17__0 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [1]),
        .I3(\ctl1/stat [1]),
        .I4(\rgf/sreg/sr [10]),
        .I5(\rgf_selc1_wb[1]_i_33_n_0 ),
        .O(\stat[1]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \stat[1]_i_18 
       (.I0(\stat[1]_i_24_n_0 ),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [8]),
        .O(\stat[1]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_18__0 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [1]),
        .O(\stat[1]_i_18__0_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[1]_i_19 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [7]),
        .O(\stat[1]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_19__0 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .O(\stat[1]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'hFF00040000000400)) 
    \stat[1]_i_1__0 
       (.I0(\fch/stat [0]),
        .I1(\fch/stat [1]),
        .I2(\stat[1]_i_2__0_n_0 ),
        .I3(\fadr[15]_INST_0_i_5_n_0 ),
        .I4(\stat[1]_i_3__1_n_0 ),
        .I5(\stat[1]_i_4_n_0 ),
        .O(\fch/fctl/stat_nx [1]));
  LUT6 #(
    .INIT(64'h000000001111FF0F)) 
    \stat[1]_i_1__1 
       (.I0(\stat[1]_i_2__1_n_0 ),
        .I1(\ctl1/stat [2]),
        .I2(\stat[1]_i_3__0_n_0 ),
        .I3(\stat_reg[1]_i_4__0_n_0 ),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [15]),
        .O(\ctl1/stat_nx [1]));
  LUT6 #(
    .INIT(64'hF2F2F222AAAAAAAA)) 
    \stat[1]_i_1__2 
       (.I0(\mem/bctl/ctl/p_0_in [5]),
        .I1(\mem/bctl/ctl/p_0_in [4]),
        .I2(fch_memacc1),
        .I3(\fch/ir0_id ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(\mem/bctl/fch_term_fl ),
        .O(\mem/bctl/ctl/stat_nx [1]));
  LUT6 #(
    .INIT(64'h00FE00FE000000FE)) 
    \stat[1]_i_2 
       (.I0(\fch/ir0 [11]),
        .I1(\bcmd[2]_INST_0_i_7_n_0 ),
        .I2(\stat[1]_i_5_n_0 ),
        .I3(\stat[0]_i_3_n_0 ),
        .I4(\stat_reg[1]_i_6_n_0 ),
        .I5(\stat[1]_i_7_n_0 ),
        .O(\stat[1]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_20 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .O(\stat[1]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \stat[1]_i_20__0 
       (.I0(\fch/ir1 [8]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [13]),
        .O(\stat[1]_i_20__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_21 
       (.I0(crdy),
        .I1(\ctl0/stat [1]),
        .O(\stat[1]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[1]_i_22 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .O(\stat[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[1]_i_23 
       (.I0(crdy),
        .I1(\rgf/sreg/sr [10]),
        .O(\stat[1]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[1]_i_24 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .O(\stat[1]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[1]_i_2__0 
       (.I0(fch_term),
        .I1(\fadr[15]_INST_0_i_8_n_0 ),
        .O(\stat[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EAEAFFEA)) 
    \stat[1]_i_2__1 
       (.I0(\stat[1]_i_5__0_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\ctl1/stat [1]),
        .I3(\stat[1]_i_6_n_0 ),
        .I4(\stat[1]_i_7__0_n_0 ),
        .I5(\stat[1]_i_8_n_0 ),
        .O(\stat[1]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF2AAAFFFFFFFF)) 
    \stat[1]_i_3 
       (.I0(\stat[1]_i_8__0_n_0 ),
        .I1(\ctl0/stat [0]),
        .I2(\ccmd[0]_INST_0_i_15_n_0 ),
        .I3(\stat[1]_i_9__0_n_0 ),
        .I4(\stat[2]_i_8__0_n_0 ),
        .I5(\stat[1]_i_10_n_0 ),
        .O(\stat[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBABB)) 
    \stat[1]_i_3__0 
       (.I0(\stat[1]_i_9_n_0 ),
        .I1(\stat[1]_i_10__0_n_0 ),
        .I2(\ctl1/stat [1]),
        .I3(\ctl1/stat [0]),
        .I4(\fch/ir1 [11]),
        .I5(\stat[1]_i_11_n_0 ),
        .O(\stat[1]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'hFF00FF47)) 
    \stat[1]_i_3__1 
       (.I0(\fch/fch_issu1 ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_issu1_fl ),
        .I3(\fch/stat [2]),
        .I4(\fch/stat [0]),
        .O(\stat[1]_i_3__1_n_0 ));
  LUT5 #(
    .INIT(32'h74300047)) 
    \stat[1]_i_4 
       (.I0(\fadr[15]_INST_0_i_8_n_0 ),
        .I1(fch_term),
        .I2(\fadr[15]_INST_0_i_4_n_0 ),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .O(\stat[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFF0DDDDFFFF)) 
    \stat[1]_i_5 
       (.I0(\stat[1]_i_14__0_n_0 ),
        .I1(crdy),
        .I2(\rgf/sreg/sr [10]),
        .I3(\fch/ir0 [9]),
        .I4(\ccmd[4]_INST_0_i_13_n_0 ),
        .I5(\stat[1]_i_15_n_0 ),
        .O(\stat[1]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \stat[1]_i_5__0 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [10]),
        .O(\stat[1]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDFFFBFFFDFFFD)) 
    \stat[1]_i_6 
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [0]),
        .I2(\stat[1]_i_15__0_n_0 ),
        .I3(\fch/ir1 [9]),
        .I4(\bcmd[2]_INST_0_i_1_n_0 ),
        .I5(brdy),
        .O(\stat[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF7F7F7F)) 
    \stat[1]_i_7 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [7]),
        .I3(\ctl0/stat [1]),
        .I4(\fch/ir0 [9]),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\stat[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \stat[1]_i_7__0 
       (.I0(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I1(\rgf/sreg/sr [10]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(\stat[2]_i_12__0_n_0 ),
        .O(\stat[1]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF444F44444444)) 
    \stat[1]_i_8 
       (.I0(\stat[2]_i_3__0_n_0 ),
        .I1(\stat[2]_i_10__0_n_0 ),
        .I2(\rgf/sreg/sr [10]),
        .I3(\fch/ir1 [9]),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\stat[1]_i_16_n_0 ),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEFFEFEFFF)) 
    \stat[1]_i_8__0 
       (.I0(\ctl0/stat [0]),
        .I1(\ctl0/stat [2]),
        .I2(\ctl0/stat [1]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [0]),
        .I5(\fch/ir0 [11]),
        .O(\stat[1]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0F055D5)) 
    \stat[1]_i_9 
       (.I0(\stat[1]_i_17__0_n_0 ),
        .I1(\stat[1]_i_18__0_n_0 ),
        .I2(\ctl1/stat [1]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [11]),
        .I5(\stat[2]_i_7__0_n_0 ),
        .O(\stat[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h023E0E0C023E020C)) 
    \stat[1]_i_9__0 
       (.I0(brdy),
        .I1(\fch/ir0 [2]),
        .I2(\ctl0/stat [2]),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [0]),
        .I5(\rgf/sreg/sr [10]),
        .O(\stat[1]_i_9__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1 
       (.I0(rst_n),
        .O(\rgf/treg/p_0_in ));
  LUT4 #(
    .INIT(16'h8000)) 
    \stat[2]_i_10 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .O(\stat[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0103030003000103)) 
    \stat[2]_i_10__0 
       (.I0(\fch/ir1 [12]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [13]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir1 [11]),
        .I5(\rgf/sreg/sr [5]),
        .O(\stat[2]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'h00000040)) 
    \stat[2]_i_11 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [6]),
        .O(\stat[2]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \stat[2]_i_11__0 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [6]),
        .O(\stat[2]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h004000F0000CF000)) 
    \stat[2]_i_12 
       (.I0(\ctl0/stat [0]),
        .I1(brdy),
        .I2(\fch/ir0 [0]),
        .I3(\ctl0/stat [2]),
        .I4(\fch/ir0 [1]),
        .I5(\ctl0/stat [1]),
        .O(\stat[2]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h9000)) 
    \stat[2]_i_12__0 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .O(\stat[2]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \stat[2]_i_13 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [10]),
        .O(\stat[2]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \stat[2]_i_13__0 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [3]),
        .O(\stat[2]_i_13__0_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[2]_i_14 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .O(\stat[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[2]_i_1__0 
       (.I0(\stat[2]_i_2__1_n_0 ),
        .I1(\stat[2]_i_3__0_n_0 ),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [14]),
        .I4(\ctl1/stat [2]),
        .I5(\stat[2]_i_4__0_n_0 ),
        .O(\ctl1/stat_nx [2]));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1__1 
       (.I0(\fch/rst_n_fl ),
        .O(\stat[2]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[2]_i_2 
       (.I0(\stat[2]_i_3_n_0 ),
        .I1(\stat[2]_i_4_n_0 ),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [14]),
        .I4(\ctl0/stat [2]),
        .I5(\stat[2]_i_5_n_0 ),
        .O(\ctl0/stat_nx [2]));
  LUT6 #(
    .INIT(64'h00000000FF005557)) 
    \stat[2]_i_2__0 
       (.I0(\fch/stat [0]),
        .I1(\fch/fch_issu1_ir ),
        .I2(\fch/stat [1]),
        .I3(\fch/stat [2]),
        .I4(\fadr[15]_INST_0_i_4_n_0 ),
        .I5(\stat[2]_i_3__1_n_0 ),
        .O(\fch/fctl/stat_nx [2]));
  LUT6 #(
    .INIT(64'h5551550055515551)) 
    \stat[2]_i_2__1 
       (.I0(\stat_reg[1]_i_4__0_n_0 ),
        .I1(\stat[2]_i_5__0_n_0 ),
        .I2(\stat[2]_i_6__0_n_0 ),
        .I3(\stat[2]_i_7__0_n_0 ),
        .I4(\stat[2]_i_8_n_0 ),
        .I5(\stat[2]_i_9__0_n_0 ),
        .O(\stat[2]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF00DF)) 
    \stat[2]_i_3 
       (.I0(\stat[2]_i_6_n_0 ),
        .I1(\ctl0/stat [0]),
        .I2(\fch/ir0 [11]),
        .I3(\stat[2]_i_7_n_0 ),
        .I4(\stat[2]_i_8__0_n_0 ),
        .I5(\stat_reg[1]_i_4_n_0 ),
        .O(\stat[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAFAEAFAFAFAFAFAE)) 
    \stat[2]_i_3__0 
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [0]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [11]),
        .I5(\rgf/sreg/sr [5]),
        .O(\stat[2]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[2]_i_3__1 
       (.I0(fch_term),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\stat[2]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAFFFFAAAAFFBE)) 
    \stat[2]_i_4 
       (.I0(\ctl0/stat [1]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [12]),
        .I5(\ctl0/stat [0]),
        .O(\stat[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEAAAAAAAAAAA)) 
    \stat[2]_i_4__0 
       (.I0(\stat[2]_i_10__0_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [10]),
        .I4(\stat[2]_i_11__0_n_0 ),
        .I5(\stat[2]_i_12__0_n_0 ),
        .O(\stat[2]_i_4__0_n_0 ));
  LUT5 #(
    .INIT(32'hEBAAAAAA)) 
    \stat[2]_i_5 
       (.I0(\stat[2]_i_9_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\ctl0/stat [0]),
        .I3(\stat[2]_i_10_n_0 ),
        .I4(\stat[2]_i_11_n_0 ),
        .O(\stat[2]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_5__0 
       (.I0(\ctl1/stat [2]),
        .I1(\ctl1/stat [1]),
        .O(\stat[2]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_6 
       (.I0(\ctl0/stat [1]),
        .I1(\ctl0/stat [2]),
        .O(\stat[2]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[2]_i_6__0 
       (.I0(\ctl1/stat [0]),
        .I1(\fch/ir1 [11]),
        .O(\stat[2]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h0202020000000000)) 
    \stat[2]_i_7 
       (.I0(\stat[2]_i_12_n_0 ),
        .I1(\ccmd[2]_INST_0_i_5_n_0 ),
        .I2(\stat[2]_i_13__0_n_0 ),
        .I3(\fch/ir0 [0]),
        .I4(\ctl0/stat [0]),
        .I5(\stat[2]_i_14_n_0 ),
        .O(\stat[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFCFFFCCCC44CC)) 
    \stat[2]_i_7__0 
       (.I0(\rgf/sreg/sr [4]),
        .I1(\fch/ir1 [12]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir1 [11]),
        .I4(\ctl1/stat [0]),
        .I5(\fch/ir1 [13]),
        .O(\stat[2]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFFFFFFFFFF)) 
    \stat[2]_i_8 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [0]),
        .I4(\ctl1/stat [0]),
        .I5(\fadr[15]_INST_0_i_20_n_0 ),
        .O(\stat[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFCFFFCCCC44CC)) 
    \stat[2]_i_8__0 
       (.I0(\rgf/sreg/sr [4]),
        .I1(\fch/ir0 [12]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir0 [11]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [13]),
        .O(\stat[2]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000007CD3)) 
    \stat[2]_i_9 
       (.I0(\fch/ir0 [12]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir0 [11]),
        .I4(\ctl0/stat [0]),
        .I5(\fch/ir0 [13]),
        .O(\stat[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h004F00000F0000C0)) 
    \stat[2]_i_9__0 
       (.I0(\ctl1/stat [0]),
        .I1(\stat[0]_i_7__0_n_0 ),
        .I2(\fch/ir1 [1]),
        .I3(\ctl1/stat [2]),
        .I4(\fch/ir1 [0]),
        .I5(\ctl1/stat [1]),
        .O(\stat[2]_i_9__0_n_0 ));
  MUXF7 \stat_reg[1]_i_4 
       (.I0(\stat[1]_i_12_n_0 ),
        .I1(\stat[1]_i_13_n_0 ),
        .O(\stat_reg[1]_i_4_n_0 ),
        .S(\stat[1]_i_11__0_n_0 ));
  MUXF7 \stat_reg[1]_i_4__0 
       (.I0(\stat[1]_i_13__0_n_0 ),
        .I1(\stat[1]_i_14_n_0 ),
        .O(\stat_reg[1]_i_4__0_n_0 ),
        .S(\stat[1]_i_12__0_n_0 ));
  MUXF7 \stat_reg[1]_i_6 
       (.I0(\stat[1]_i_16__0_n_0 ),
        .I1(\stat[1]_i_17_n_0 ),
        .O(\stat_reg[1]_i_6_n_0 ),
        .S(\fch/ir0 [8]));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .O(tout__1_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[14]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[6]),
        .O(tout__1_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .O(tout__1_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[13]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[5]),
        .O(tout__1_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_3
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(tout__1_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_3__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[4]),
        .O(tout__1_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__0_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(tout__1_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__0_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[3]),
        .O(tout__1_carry__0_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_5
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[7]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .I3(tout__1_carry__0_i_1_n_0),
        .O(tout__1_carry__0_i_5_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_5__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[15]_INST_0_i_18_n_0 ),
        .I2(a1bus_0[7]),
        .I3(tout__1_carry__0_i_1__0_n_0),
        .O(tout__1_carry__0_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .I3(tout__1_carry__0_i_2_n_0),
        .O(tout__1_carry__0_i_6_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[14]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[6]),
        .I3(tout__1_carry__0_i_2__0_n_0),
        .O(tout__1_carry__0_i_6__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_7
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .I3(tout__1_carry__0_i_3_n_0),
        .O(tout__1_carry__0_i_7_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_7__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[13]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[5]),
        .I3(tout__1_carry__0_i_3__0_n_0),
        .O(tout__1_carry__0_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__0_i_8
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .I3(tout__1_carry__0_i_4_n_0),
        .O(tout__1_carry__0_i_8_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__0_i_8__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[12]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[4]),
        .I3(tout__1_carry__0_i_4__0_n_0),
        .O(tout__1_carry__0_i_8__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[10]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(tout__1_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[10]),
        .O(tout__1_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[9]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(tout__1_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[9]),
        .O(tout__1_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_3
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[8]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(tout__1_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__1_i_3__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[8]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[8]),
        .O(tout__1_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[7]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .O(tout__1_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__1_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[15]_INST_0_i_18_n_0 ),
        .I2(a1bus_0[7]),
        .O(tout__1_carry__1_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_5
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[11]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .I3(tout__1_carry__1_i_1_n_0),
        .O(tout__1_carry__1_i_5_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_5__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[11]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[11]),
        .I3(tout__1_carry__1_i_1__0_n_0),
        .O(tout__1_carry__1_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[10]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .I3(tout__1_carry__1_i_2_n_0),
        .O(tout__1_carry__1_i_6_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[10]),
        .I3(tout__1_carry__1_i_2__0_n_0),
        .O(tout__1_carry__1_i_6__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_7
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[9]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .I3(tout__1_carry__1_i_3_n_0),
        .O(tout__1_carry__1_i_7_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_7__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[9]),
        .I3(tout__1_carry__1_i_3__0_n_0),
        .O(tout__1_carry__1_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__1_i_8
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[8]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .I3(tout__1_carry__1_i_4_n_0),
        .O(tout__1_carry__1_i_8_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__1_i_8__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[8]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[8]),
        .I3(tout__1_carry__1_i_4__0_n_0),
        .O(tout__1_carry__1_i_8__0_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    tout__1_carry__2_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(tout__1_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    tout__1_carry__2_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[15]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[15]),
        .O(tout__1_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[13]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .O(tout__1_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[13]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[13]),
        .O(tout__1_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_3
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[12]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .O(tout__1_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_3__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[12]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[12]),
        .O(tout__1_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry__2_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[11]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .O(tout__1_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry__2_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[11]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[11]),
        .O(tout__1_carry__2_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hC33C5AA5)) 
    tout__1_carry__2_i_5
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[14]_INST_0_i_2_n_0 ),
        .I2(\bdatw[15]_INST_0_i_2_n_0 ),
        .I3(a1bus_0[15]),
        .I4(a1bus_0[14]),
        .O(tout__1_carry__2_i_5_n_0));
  LUT5 #(
    .INIT(32'hC33C9696)) 
    tout__1_carry__2_i_5__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\bdatw[14]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[14]),
        .O(tout__1_carry__2_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[14]_INST_0_i_1_n_0 ),
        .I2(tout__1_carry__2_i_2_n_0),
        .I3(a0bus_0[14]),
        .O(tout__1_carry__2_i_6_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[14]_INST_0_i_2_n_0 ),
        .I2(tout__1_carry__2_i_2__0_n_0),
        .I3(a1bus_0[14]),
        .O(tout__1_carry__2_i_6__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_7
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[13]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .I3(tout__1_carry__2_i_3_n_0),
        .O(tout__1_carry__2_i_7_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_7__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[13]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[13]),
        .I3(tout__1_carry__2_i_3__0_n_0),
        .O(tout__1_carry__2_i_7__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry__2_i_8
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[12]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .I3(tout__1_carry__2_i_4_n_0),
        .O(tout__1_carry__2_i_8_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry__2_i_8__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[12]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[12]),
        .I3(tout__1_carry__2_i_4__0_n_0),
        .O(tout__1_carry__2_i_8__0_n_0));
  LUT3 #(
    .INIT(8'h6F)) 
    tout__1_carry__3_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(tout__1_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h9F)) 
    tout__1_carry__3_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[15]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[15]),
        .O(tout__1_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h96)) 
    tout__1_carry__3_i_2
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[15]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[15]),
        .O(tout__1_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    tout__1_carry__3_i_2__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(tout__1_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'hF9)) 
    tout__1_carry__3_i_3
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[15]_INST_0_i_2_n_0 ),
        .I2(a1bus_0[15]),
        .O(tout__1_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'hF6)) 
    tout__1_carry__3_i_3__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bdatw[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(tout__1_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_1
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(tout__1_carry_i_1_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    tout__1_carry_i_10
       (.I0(\ccmd[2]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .O(tout__1_carry_i_10_n_0));
  LUT4 #(
    .INIT(16'h0010)) 
    tout__1_carry_i_10__0
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .O(tout__1_carry_i_10__0_n_0));
  LUT6 #(
    .INIT(64'h4000400040004055)) 
    tout__1_carry_i_11
       (.I0(\ctl0/stat [2]),
        .I1(\ccmd[0]_INST_0_i_7_n_0 ),
        .I2(\ccmd[0]_INST_0_i_6_n_0 ),
        .I3(\ccmd[0]_INST_0_i_5_n_0 ),
        .I4(\ccmd[0]_INST_0_i_4_n_0 ),
        .I5(tout__1_carry_i_13_n_0),
        .O(tout__1_carry_i_11_n_0));
  LUT4 #(
    .INIT(16'hFFEF)) 
    tout__1_carry_i_11__0
       (.I0(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(tout__1_carry_i_11__0_n_0));
  LUT6 #(
    .INIT(64'h000000000000DD0D)) 
    tout__1_carry_i_12
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(tout__1_carry_i_13__0_n_0),
        .I2(\rgf_selc1_wb[0]_i_7_n_0 ),
        .I3(tout__1_carry_i_14_n_0),
        .I4(tout__1_carry_i_15_n_0),
        .I5(tout__1_carry_i_16_n_0),
        .O(tout__1_carry_i_12_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    tout__1_carry_i_12__0
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .O(tout__1_carry_i_12__0_n_0));
  LUT6 #(
    .INIT(64'hA200A2000000A200)) 
    tout__1_carry_i_13
       (.I0(\ccmd[0]_INST_0_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_36_n_0 ),
        .I2(\ccmd[0]_INST_0_i_9_n_0 ),
        .I3(\bdatw[8]_INST_0_i_17_n_0 ),
        .I4(\fch/ir0 [13]),
        .I5(\bcmd[1]_INST_0_i_1_n_0 ),
        .O(tout__1_carry_i_13_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00F8F8)) 
    tout__1_carry_i_13__0
       (.I0(\ctl1/stat [1]),
        .I1(\ctl1/stat [0]),
        .I2(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I3(tout__1_carry_i_17_n_0),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [15]),
        .O(tout__1_carry_i_13__0_n_0));
  LUT6 #(
    .INIT(64'hFFFBFFFBF00BFFFF)) 
    tout__1_carry_i_14
       (.I0(\ctl1/stat [0]),
        .I1(\ctl1/stat [1]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [0]),
        .O(tout__1_carry_i_14_n_0));
  LUT6 #(
    .INIT(64'h50007000A0000000)) 
    tout__1_carry_i_15
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [11]),
        .I2(\badr[15]_INST_0_i_144_n_0 ),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [14]),
        .O(tout__1_carry_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000000000002400)) 
    tout__1_carry_i_16
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I4(\ctl1/stat [0]),
        .I5(\ctl1/stat [1]),
        .O(tout__1_carry_i_16_n_0));
  LUT6 #(
    .INIT(64'h00F700FF000000FF)) 
    tout__1_carry_i_17
       (.I0(\fch/ir1 [7]),
        .I1(\badr[15]_INST_0_i_213_n_0 ),
        .I2(tout__1_carry_i_18_n_0),
        .I3(tout__1_carry_i_19_n_0),
        .I4(\fch/ir1 [8]),
        .I5(\rgf_selc1_wb[0]_i_11_n_0 ),
        .O(tout__1_carry_i_17_n_0));
  LUT6 #(
    .INIT(64'hAAAAAA8AAAAA02A8)) 
    tout__1_carry_i_18
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [5]),
        .I5(\ctl1/stat [0]),
        .O(tout__1_carry_i_18_n_0));
  LUT6 #(
    .INIT(64'h0000030003001111)) 
    tout__1_carry_i_19
       (.I0(tout__1_carry_i_20_n_0),
        .I1(\ctl1/stat [1]),
        .I2(\ctl1/stat [0]),
        .I3(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(tout__1_carry_i_19_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry_i_1__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .O(tout__1_carry_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h90)) 
    tout__1_carry_i_2
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(tout__1_carry_i_2_n_0));
  LUT4 #(
    .INIT(16'hFFF7)) 
    tout__1_carry_i_20
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [9]),
        .I3(\ctl1/stat [0]),
        .O(tout__1_carry_i_20_n_0));
  LUT3 #(
    .INIT(8'h60)) 
    tout__1_carry_i_2__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(a1bus_0[1]),
        .O(tout__1_carry_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hF9F999FF90900099)) 
    tout__1_carry_i_3
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(tout__1_carry_i_8_n_0),
        .I2(tout__1_carry_i_9__0_n_0),
        .I3(tout__1_carry_i_10__0_n_0),
        .I4(\rgf/sreg/sr [6]),
        .I5(a1bus_0[0]),
        .O(tout__1_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h6F06)) 
    tout__1_carry_i_3__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(tout__1_carry_i_9_n_0),
        .I3(a0bus_0[0]),
        .O(tout__1_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_4
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .I3(tout__1_carry_i_1_n_0),
        .O(tout__1_carry_i_4_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_4__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[11]_INST_0_i_16_n_0 ),
        .I2(a1bus_0[3]),
        .I3(tout__1_carry_i_1__0_n_0),
        .O(tout__1_carry_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_5
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .I3(tout__1_carry_i_2_n_0),
        .O(tout__1_carry_i_5_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_5__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[10]_INST_0_i_14_n_0 ),
        .I2(a1bus_0[2]),
        .I3(tout__1_carry_i_2__0_n_0),
        .O(tout__1_carry_i_5__0_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_6
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .I3(tout__1_carry_i_3__0_n_0),
        .O(tout__1_carry_i_6_n_0));
  LUT4 #(
    .INIT(16'h6996)) 
    tout__1_carry_i_6__0
       (.I0(tout__1_carry_i_8_n_0),
        .I1(\bdatw[9]_INST_0_i_13_n_0 ),
        .I2(a1bus_0[1]),
        .I3(tout__1_carry_i_3_n_0),
        .O(tout__1_carry_i_6__0_n_0));
  LUT6 #(
    .INIT(64'h9696669969699966)) 
    tout__1_carry_i_7
       (.I0(\bdatw[8]_INST_0_i_14_n_0 ),
        .I1(tout__1_carry_i_8_n_0),
        .I2(tout__1_carry_i_9__0_n_0),
        .I3(tout__1_carry_i_10__0_n_0),
        .I4(\rgf/sreg/sr [6]),
        .I5(a1bus_0[0]),
        .O(tout__1_carry_i_7_n_0));
  LUT4 #(
    .INIT(16'h9669)) 
    tout__1_carry_i_7__0
       (.I0(tout__1_carry_i_8__0_n_0),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(tout__1_carry_i_9_n_0),
        .I3(a0bus_0[0]),
        .O(tout__1_carry_i_7__0_n_0));
  LUT3 #(
    .INIT(8'h45)) 
    tout__1_carry_i_8
       (.I0(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I1(tout__1_carry_i_9__0_n_0),
        .I2(tout__1_carry_i_11__0_n_0),
        .O(tout__1_carry_i_8_n_0));
  LUT6 #(
    .INIT(64'hEEEEFFEEFFFEFFFE)) 
    tout__1_carry_i_8__0
       (.I0(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .I2(tout__1_carry_i_10_n_0),
        .I3(tout__1_carry_i_11_n_0),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .O(tout__1_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'h0002FF02)) 
    tout__1_carry_i_9
       (.I0(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I3(\rgf/sreg/sr [6]),
        .I4(tout__1_carry_i_12__0_n_0),
        .O(tout__1_carry_i_9_n_0));
  LUT4 #(
    .INIT(16'h0E00)) 
    tout__1_carry_i_9__0
       (.I0(\ctl1/stat [2]),
        .I1(tout__1_carry_i_12_n_0),
        .I2(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .O(tout__1_carry_i_9__0_n_0));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [0]),
        .O(\rgf/treg/p_1_in [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [10]),
        .O(\rgf/treg/p_1_in [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [11]),
        .O(\rgf/treg/p_1_in [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [12]),
        .O(\rgf/treg/p_1_in [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [13]),
        .O(\rgf/treg/p_1_in [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [14]),
        .O(\rgf/treg/p_1_in [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [15]),
        .O(\rgf/treg/p_1_in [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\sr[11]_i_9_n_0 ),
        .O(\rgf/c1bus_sel_cr [4]));
  LUT4 #(
    .INIT(16'h0010)) 
    \tr[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\pc[15]_i_7_n_0 ),
        .O(\rgf/c0bus_sel_cr [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [1]),
        .O(\rgf/treg/p_1_in [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [2]),
        .O(\rgf/treg/p_1_in [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [3]),
        .O(\rgf/treg/p_1_in [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [4]),
        .O(\rgf/treg/p_1_in [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [5]),
        .O(\rgf/treg/p_1_in [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [6]),
        .O(\rgf/treg/p_1_in [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [7]),
        .O(\rgf/treg/p_1_in [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [8]),
        .O(\rgf/treg/p_1_in [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [9]),
        .O(\rgf/treg/p_1_in [9]));
endmodule
