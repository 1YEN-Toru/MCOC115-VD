
(* STRUCTURAL_NETLIST = "yes" *)
module nihoniumss
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdat,
    bdatr,
    .fadr({\^fadr [15],\^fadr [14],\^fadr [13],\^fadr [12],\^fadr [11],\^fadr [10],\^fadr [9],\^fadr [8],\^fadr [7],\^fadr [6],\^fadr [5],\^fadr [4],\^fadr [3],\^fadr [2],\^fadr [1],\rgf/pcnt/pc [0]}),
    bcmd,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o,
    niss_dsp_c0,
    niss_dsp_c1,
    niss_dsp_a0,
    niss_dsp_a1,
    niss_dsp_b0,
    niss_dsp_b1);
//
//	Nihonium-SS 16/32 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2023/10/28	ver.1.16
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.14
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.12
//		instruction: divur, divsr, mulur, mulsr
//
//	2023/03/18	ver.1.10
//		instruction: jall, rtnl, pushcl, popcl
//
//	2023/03/11	ver.1.08
//		corresponding to 32 bit memory bus
//
//	2023/02/11	ver.1.06
//		instruction: fdown
//
//	2022/10/22	ver.1.04
//		corresponding to interrupt vector / level
//
//	2022/06/04	ver.1.02
//		instruction: csft, csfti
//
//	2022/05/21	ver.1.00
//		Nihonium-SS: Super Scalar Edition
//
// ================================
//
//	2022/04/09	ver.1.00
//		external 16 bit / internal 32 bit CPU
//		32 bit divider from divc32 ver.1.00
//		extended instructions:
//			link, unlk, brn, ldli, cendl, pushl, popl,
//			exsgl, exzrl, ldl, stl, ldlsp, stlsp
//
// ================================
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [31:0]fdat;
  input [31:0]bdatr;
  output [3:0]bcmd;
  output [31:0]badr;
  output [31:0]bdatw;
  input crdy;
  input [31:0]cbus_i;
  output [4:0]ccmd;
  output [31:0]abus_o;
  output [31:0]bbus_o;
  input [65:0]niss_dsp_c0;
  input [65:0]niss_dsp_c1;
  output [32:0]niss_dsp_a0;
  output [32:0]niss_dsp_a1;
  output [32:0]niss_dsp_b0;
  output [32:0]niss_dsp_b1;
     output [15:1]\^fadr ;
     output [15:0]\rgf/pcnt/pc ;

  wire \<const0> ;
  wire \<const1> ;
  wire [31:0]a0bus_0;
  wire [31:0]a1bus_0;
  wire [31:0]abus_o;
  wire [4:0]acmd1;
  wire add_out0_carry__0_i_13__0_n_0;
  wire add_out0_carry__0_i_13_n_0;
  wire add_out0_carry__0_i_14__0_n_0;
  wire add_out0_carry__0_i_14_n_0;
  wire add_out0_carry__0_i_15__0_n_0;
  wire add_out0_carry__0_i_15_n_0;
  wire add_out0_carry__0_i_16__0_n_0;
  wire add_out0_carry__0_i_16_n_0;
  wire add_out0_carry__0_i_1__0_n_0;
  wire add_out0_carry__0_i_1_n_0;
  wire add_out0_carry__0_i_2__0_n_0;
  wire add_out0_carry__0_i_2_n_0;
  wire add_out0_carry__0_i_3__0_n_0;
  wire add_out0_carry__0_i_3_n_0;
  wire add_out0_carry__0_i_4__0_n_0;
  wire add_out0_carry__0_i_4_n_0;
  wire add_out0_carry__0_i_5__0_n_0;
  wire add_out0_carry__0_i_5_n_0;
  wire add_out0_carry__0_i_6__0_n_0;
  wire add_out0_carry__0_i_6_n_0;
  wire add_out0_carry__0_i_7__0_n_0;
  wire add_out0_carry__0_i_7_n_0;
  wire add_out0_carry__0_i_8__0_n_0;
  wire add_out0_carry__0_i_8_n_0;
  wire add_out0_carry__1_i_13__0_n_0;
  wire add_out0_carry__1_i_13_n_0;
  wire add_out0_carry__1_i_14__0_n_0;
  wire add_out0_carry__1_i_14_n_0;
  wire add_out0_carry__1_i_15__0_n_0;
  wire add_out0_carry__1_i_15_n_0;
  wire add_out0_carry__1_i_16__0_n_0;
  wire add_out0_carry__1_i_16_n_0;
  wire add_out0_carry__1_i_1__0_n_0;
  wire add_out0_carry__1_i_1_n_0;
  wire add_out0_carry__1_i_2__0_n_0;
  wire add_out0_carry__1_i_2_n_0;
  wire add_out0_carry__1_i_3__0_n_0;
  wire add_out0_carry__1_i_3_n_0;
  wire add_out0_carry__1_i_4__0_n_0;
  wire add_out0_carry__1_i_4_n_0;
  wire add_out0_carry__1_i_5__0_n_0;
  wire add_out0_carry__1_i_5_n_0;
  wire add_out0_carry__1_i_6__0_n_0;
  wire add_out0_carry__1_i_6_n_0;
  wire add_out0_carry__1_i_7__0_n_0;
  wire add_out0_carry__1_i_7_n_0;
  wire add_out0_carry__1_i_8__0_n_0;
  wire add_out0_carry__1_i_8_n_0;
  wire add_out0_carry__2_i_13__0_n_0;
  wire add_out0_carry__2_i_13_n_0;
  wire add_out0_carry__2_i_14__0_n_0;
  wire add_out0_carry__2_i_14_n_0;
  wire add_out0_carry__2_i_15__0_n_0;
  wire add_out0_carry__2_i_15_n_0;
  wire add_out0_carry__2_i_16__0_n_0;
  wire add_out0_carry__2_i_16_n_0;
  wire add_out0_carry__2_i_1__0_n_0;
  wire add_out0_carry__2_i_1_n_0;
  wire add_out0_carry__2_i_2__0_n_0;
  wire add_out0_carry__2_i_2_n_0;
  wire add_out0_carry__2_i_3__0_n_0;
  wire add_out0_carry__2_i_3_n_0;
  wire add_out0_carry__2_i_4__0_n_0;
  wire add_out0_carry__2_i_4_n_0;
  wire add_out0_carry__2_i_5__0_n_0;
  wire add_out0_carry__2_i_5_n_0;
  wire add_out0_carry__2_i_6__0_n_0;
  wire add_out0_carry__2_i_6_n_0;
  wire add_out0_carry__2_i_7__0_n_0;
  wire add_out0_carry__2_i_7_n_0;
  wire add_out0_carry__2_i_8__0_n_0;
  wire add_out0_carry__2_i_8_n_0;
  wire add_out0_carry__3_i_13__0_n_0;
  wire add_out0_carry__3_i_13_n_0;
  wire add_out0_carry__3_i_14__0_n_0;
  wire add_out0_carry__3_i_14_n_0;
  wire add_out0_carry__3_i_15__0_n_0;
  wire add_out0_carry__3_i_15_n_0;
  wire add_out0_carry__3_i_16__0_n_0;
  wire add_out0_carry__3_i_16_n_0;
  wire add_out0_carry__3_i_1__0_n_0;
  wire add_out0_carry__3_i_1_n_0;
  wire add_out0_carry__3_i_2__0_n_0;
  wire add_out0_carry__3_i_2_n_0;
  wire add_out0_carry__3_i_3__0_n_0;
  wire add_out0_carry__3_i_3_n_0;
  wire add_out0_carry__3_i_4__0_n_0;
  wire add_out0_carry__3_i_4_n_0;
  wire add_out0_carry__3_i_5__0_n_0;
  wire add_out0_carry__3_i_5_n_0;
  wire add_out0_carry__3_i_6__0_n_0;
  wire add_out0_carry__3_i_6_n_0;
  wire add_out0_carry__3_i_7__0_n_0;
  wire add_out0_carry__3_i_7_n_0;
  wire add_out0_carry__3_i_8__0_n_0;
  wire add_out0_carry__3_i_8_n_0;
  wire add_out0_carry__4_i_13__0_n_0;
  wire add_out0_carry__4_i_13_n_0;
  wire add_out0_carry__4_i_14__0_n_0;
  wire add_out0_carry__4_i_14_n_0;
  wire add_out0_carry__4_i_15__0_n_0;
  wire add_out0_carry__4_i_15_n_0;
  wire add_out0_carry__4_i_16__0_n_0;
  wire add_out0_carry__4_i_16_n_0;
  wire add_out0_carry__4_i_1__0_n_0;
  wire add_out0_carry__4_i_1_n_0;
  wire add_out0_carry__4_i_2__0_n_0;
  wire add_out0_carry__4_i_2_n_0;
  wire add_out0_carry__4_i_3__0_n_0;
  wire add_out0_carry__4_i_3_n_0;
  wire add_out0_carry__4_i_4__0_n_0;
  wire add_out0_carry__4_i_4_n_0;
  wire add_out0_carry__4_i_5__0_n_0;
  wire add_out0_carry__4_i_5_n_0;
  wire add_out0_carry__4_i_6__0_n_0;
  wire add_out0_carry__4_i_6_n_0;
  wire add_out0_carry__4_i_7__0_n_0;
  wire add_out0_carry__4_i_7_n_0;
  wire add_out0_carry__4_i_8__0_n_0;
  wire add_out0_carry__4_i_8_n_0;
  wire add_out0_carry__5_i_13__0_n_0;
  wire add_out0_carry__5_i_13_n_0;
  wire add_out0_carry__5_i_14__0_n_0;
  wire add_out0_carry__5_i_14_n_0;
  wire add_out0_carry__5_i_15__0_n_0;
  wire add_out0_carry__5_i_15_n_0;
  wire add_out0_carry__5_i_16__0_n_0;
  wire add_out0_carry__5_i_16_n_0;
  wire add_out0_carry__5_i_1__0_n_0;
  wire add_out0_carry__5_i_1_n_0;
  wire add_out0_carry__5_i_2__0_n_0;
  wire add_out0_carry__5_i_2_n_0;
  wire add_out0_carry__5_i_3__0_n_0;
  wire add_out0_carry__5_i_3_n_0;
  wire add_out0_carry__5_i_4__0_n_0;
  wire add_out0_carry__5_i_4_n_0;
  wire add_out0_carry__5_i_5__0_n_0;
  wire add_out0_carry__5_i_5_n_0;
  wire add_out0_carry__5_i_6__0_n_0;
  wire add_out0_carry__5_i_6_n_0;
  wire add_out0_carry__5_i_7__0_n_0;
  wire add_out0_carry__5_i_7_n_0;
  wire add_out0_carry__5_i_8__0_n_0;
  wire add_out0_carry__5_i_8_n_0;
  wire add_out0_carry__6_i_11__0_n_0;
  wire add_out0_carry__6_i_11_n_0;
  wire add_out0_carry__6_i_12__0_n_0;
  wire add_out0_carry__6_i_12_n_0;
  wire add_out0_carry__6_i_13__0_n_0;
  wire add_out0_carry__6_i_13_n_0;
  wire add_out0_carry__6_i_1__0_n_0;
  wire add_out0_carry__6_i_1_n_0;
  wire add_out0_carry__6_i_2__0_n_0;
  wire add_out0_carry__6_i_2_n_0;
  wire add_out0_carry__6_i_3__0_n_0;
  wire add_out0_carry__6_i_3_n_0;
  wire add_out0_carry__6_i_4__0_n_0;
  wire add_out0_carry__6_i_4_n_0;
  wire add_out0_carry__6_i_5__0_n_0;
  wire add_out0_carry__6_i_5_n_0;
  wire add_out0_carry__6_i_6__0_n_0;
  wire add_out0_carry__6_i_6_n_0;
  wire add_out0_carry__6_i_7__0_n_0;
  wire add_out0_carry__6_i_7_n_0;
  wire add_out0_carry_i_13__0_n_0;
  wire add_out0_carry_i_13_n_0;
  wire add_out0_carry_i_14__0_n_0;
  wire add_out0_carry_i_14_n_0;
  wire add_out0_carry_i_15__0_n_0;
  wire add_out0_carry_i_15_n_0;
  wire add_out0_carry_i_16__0_n_0;
  wire add_out0_carry_i_16_n_0;
  wire add_out0_carry_i_1__0_n_0;
  wire add_out0_carry_i_1_n_0;
  wire add_out0_carry_i_2__0_n_0;
  wire add_out0_carry_i_2_n_0;
  wire add_out0_carry_i_3__0_n_0;
  wire add_out0_carry_i_3_n_0;
  wire add_out0_carry_i_4__0_n_0;
  wire add_out0_carry_i_4_n_0;
  wire add_out0_carry_i_5__0_n_0;
  wire add_out0_carry_i_5_n_0;
  wire add_out0_carry_i_6__0_n_0;
  wire add_out0_carry_i_6_n_0;
  wire add_out0_carry_i_7__0_n_0;
  wire add_out0_carry_i_7_n_0;
  wire add_out0_carry_i_8__0_n_0;
  wire add_out0_carry_i_8_n_0;
  wire \alu0/art/add/p_0_in ;
  wire [34:18]\alu0/art/add/tout ;
  wire [32:32]\alu0/art/p_0_in__0 ;
  wire [16:16]\alu0/asr0 ;
  wire [31:0]\alu0/div/add_out ;
  wire \alu0/div/chg_quo_sgn ;
  wire \alu0/div/chg_rem_sgn ;
  wire \alu0/div/dadd/add_out0_carry__0_n_0 ;
  wire \alu0/div/dadd/add_out0_carry__0_n_1 ;
  wire \alu0/div/dadd/add_out0_carry__0_n_2 ;
  wire \alu0/div/dadd/add_out0_carry__0_n_3 ;
  wire \alu0/div/dadd/add_out0_carry__1_n_0 ;
  wire \alu0/div/dadd/add_out0_carry__1_n_1 ;
  wire \alu0/div/dadd/add_out0_carry__1_n_2 ;
  wire \alu0/div/dadd/add_out0_carry__1_n_3 ;
  wire \alu0/div/dadd/add_out0_carry__2_n_0 ;
  wire \alu0/div/dadd/add_out0_carry__2_n_1 ;
  wire \alu0/div/dadd/add_out0_carry__2_n_2 ;
  wire \alu0/div/dadd/add_out0_carry__2_n_3 ;
  wire \alu0/div/dadd/add_out0_carry__3_n_0 ;
  wire \alu0/div/dadd/add_out0_carry__3_n_1 ;
  wire \alu0/div/dadd/add_out0_carry__3_n_2 ;
  wire \alu0/div/dadd/add_out0_carry__3_n_3 ;
  wire \alu0/div/dadd/add_out0_carry__4_n_0 ;
  wire \alu0/div/dadd/add_out0_carry__4_n_1 ;
  wire \alu0/div/dadd/add_out0_carry__4_n_2 ;
  wire \alu0/div/dadd/add_out0_carry__4_n_3 ;
  wire \alu0/div/dadd/add_out0_carry__5_n_0 ;
  wire \alu0/div/dadd/add_out0_carry__5_n_1 ;
  wire \alu0/div/dadd/add_out0_carry__5_n_2 ;
  wire \alu0/div/dadd/add_out0_carry__5_n_3 ;
  wire \alu0/div/dadd/add_out0_carry__6_n_1 ;
  wire \alu0/div/dadd/add_out0_carry__6_n_2 ;
  wire \alu0/div/dadd/add_out0_carry__6_n_3 ;
  wire \alu0/div/dadd/add_out0_carry_n_0 ;
  wire \alu0/div/dadd/add_out0_carry_n_1 ;
  wire \alu0/div/dadd/add_out0_carry_n_2 ;
  wire \alu0/div/dadd/add_out0_carry_n_3 ;
  wire \alu0/div/dctl/dctl_long_f ;
  wire \alu0/div/dctl/dctl_sign ;
  wire \alu0/div/dctl/dctl_sign_f ;
  wire \alu0/div/dctl/fsm/chg_rem_sgn0 ;
  wire [3:0]\alu0/div/dctl/fsm/dctl_next ;
  wire \alu0/div/dctl/fsm/set_sgn ;
  wire \alu0/div/dctl_long ;
  wire [3:0]\alu0/div/dctl_stat ;
  wire [64:0]\alu0/div/den ;
  wire [3:3]\alu0/div/den2 ;
  wire [31:0]\alu0/div/dso_0 ;
  wire [0:0]\alu0/div/fdiv/p_1_in3_in ;
  wire [0:0]\alu0/div/fdiv/p_1_in5_in ;
  wire \alu0/div/fdiv/rem0_carry__0_n_0 ;
  wire \alu0/div/fdiv/rem0_carry__0_n_1 ;
  wire \alu0/div/fdiv/rem0_carry__0_n_2 ;
  wire \alu0/div/fdiv/rem0_carry__0_n_3 ;
  wire \alu0/div/fdiv/rem0_carry__1_n_0 ;
  wire \alu0/div/fdiv/rem0_carry__1_n_1 ;
  wire \alu0/div/fdiv/rem0_carry__1_n_2 ;
  wire \alu0/div/fdiv/rem0_carry__1_n_3 ;
  wire \alu0/div/fdiv/rem0_carry__2_n_0 ;
  wire \alu0/div/fdiv/rem0_carry__2_n_1 ;
  wire \alu0/div/fdiv/rem0_carry__2_n_2 ;
  wire \alu0/div/fdiv/rem0_carry__2_n_3 ;
  wire \alu0/div/fdiv/rem0_carry__3_n_0 ;
  wire \alu0/div/fdiv/rem0_carry__3_n_1 ;
  wire \alu0/div/fdiv/rem0_carry__3_n_2 ;
  wire \alu0/div/fdiv/rem0_carry__3_n_3 ;
  wire \alu0/div/fdiv/rem0_carry__4_n_0 ;
  wire \alu0/div/fdiv/rem0_carry__4_n_1 ;
  wire \alu0/div/fdiv/rem0_carry__4_n_2 ;
  wire \alu0/div/fdiv/rem0_carry__4_n_3 ;
  wire \alu0/div/fdiv/rem0_carry__5_n_0 ;
  wire \alu0/div/fdiv/rem0_carry__5_n_1 ;
  wire \alu0/div/fdiv/rem0_carry__5_n_2 ;
  wire \alu0/div/fdiv/rem0_carry__5_n_3 ;
  wire \alu0/div/fdiv/rem0_carry__6_n_0 ;
  wire \alu0/div/fdiv/rem0_carry__6_n_1 ;
  wire \alu0/div/fdiv/rem0_carry__6_n_2 ;
  wire \alu0/div/fdiv/rem0_carry__6_n_3 ;
  wire \alu0/div/fdiv/rem0_carry_n_0 ;
  wire \alu0/div/fdiv/rem0_carry_n_1 ;
  wire \alu0/div/fdiv/rem0_carry_n_2 ;
  wire \alu0/div/fdiv/rem0_carry_n_3 ;
  wire \alu0/div/fdiv/rem1_carry__0_n_0 ;
  wire \alu0/div/fdiv/rem1_carry__0_n_1 ;
  wire \alu0/div/fdiv/rem1_carry__0_n_2 ;
  wire \alu0/div/fdiv/rem1_carry__0_n_3 ;
  wire \alu0/div/fdiv/rem1_carry__1_n_0 ;
  wire \alu0/div/fdiv/rem1_carry__1_n_1 ;
  wire \alu0/div/fdiv/rem1_carry__1_n_2 ;
  wire \alu0/div/fdiv/rem1_carry__1_n_3 ;
  wire \alu0/div/fdiv/rem1_carry__2_n_0 ;
  wire \alu0/div/fdiv/rem1_carry__2_n_1 ;
  wire \alu0/div/fdiv/rem1_carry__2_n_2 ;
  wire \alu0/div/fdiv/rem1_carry__2_n_3 ;
  wire \alu0/div/fdiv/rem1_carry__3_n_0 ;
  wire \alu0/div/fdiv/rem1_carry__3_n_1 ;
  wire \alu0/div/fdiv/rem1_carry__3_n_2 ;
  wire \alu0/div/fdiv/rem1_carry__3_n_3 ;
  wire \alu0/div/fdiv/rem1_carry__4_n_0 ;
  wire \alu0/div/fdiv/rem1_carry__4_n_1 ;
  wire \alu0/div/fdiv/rem1_carry__4_n_2 ;
  wire \alu0/div/fdiv/rem1_carry__4_n_3 ;
  wire \alu0/div/fdiv/rem1_carry__5_n_0 ;
  wire \alu0/div/fdiv/rem1_carry__5_n_1 ;
  wire \alu0/div/fdiv/rem1_carry__5_n_2 ;
  wire \alu0/div/fdiv/rem1_carry__5_n_3 ;
  wire \alu0/div/fdiv/rem1_carry__6_n_0 ;
  wire \alu0/div/fdiv/rem1_carry__6_n_1 ;
  wire \alu0/div/fdiv/rem1_carry__6_n_2 ;
  wire \alu0/div/fdiv/rem1_carry__6_n_3 ;
  wire \alu0/div/fdiv/rem1_carry_n_0 ;
  wire \alu0/div/fdiv/rem1_carry_n_1 ;
  wire \alu0/div/fdiv/rem1_carry_n_2 ;
  wire \alu0/div/fdiv/rem1_carry_n_3 ;
  wire \alu0/div/fdiv/rem2_carry__0_n_0 ;
  wire \alu0/div/fdiv/rem2_carry__0_n_1 ;
  wire \alu0/div/fdiv/rem2_carry__0_n_2 ;
  wire \alu0/div/fdiv/rem2_carry__0_n_3 ;
  wire \alu0/div/fdiv/rem2_carry__1_n_0 ;
  wire \alu0/div/fdiv/rem2_carry__1_n_1 ;
  wire \alu0/div/fdiv/rem2_carry__1_n_2 ;
  wire \alu0/div/fdiv/rem2_carry__1_n_3 ;
  wire \alu0/div/fdiv/rem2_carry__2_n_0 ;
  wire \alu0/div/fdiv/rem2_carry__2_n_1 ;
  wire \alu0/div/fdiv/rem2_carry__2_n_2 ;
  wire \alu0/div/fdiv/rem2_carry__2_n_3 ;
  wire \alu0/div/fdiv/rem2_carry__3_n_0 ;
  wire \alu0/div/fdiv/rem2_carry__3_n_1 ;
  wire \alu0/div/fdiv/rem2_carry__3_n_2 ;
  wire \alu0/div/fdiv/rem2_carry__3_n_3 ;
  wire \alu0/div/fdiv/rem2_carry__4_n_0 ;
  wire \alu0/div/fdiv/rem2_carry__4_n_1 ;
  wire \alu0/div/fdiv/rem2_carry__4_n_2 ;
  wire \alu0/div/fdiv/rem2_carry__4_n_3 ;
  wire \alu0/div/fdiv/rem2_carry__5_n_0 ;
  wire \alu0/div/fdiv/rem2_carry__5_n_1 ;
  wire \alu0/div/fdiv/rem2_carry__5_n_2 ;
  wire \alu0/div/fdiv/rem2_carry__5_n_3 ;
  wire \alu0/div/fdiv/rem2_carry__6_n_0 ;
  wire \alu0/div/fdiv/rem2_carry__6_n_1 ;
  wire \alu0/div/fdiv/rem2_carry__6_n_2 ;
  wire \alu0/div/fdiv/rem2_carry__6_n_3 ;
  wire \alu0/div/fdiv/rem2_carry_n_0 ;
  wire \alu0/div/fdiv/rem2_carry_n_1 ;
  wire \alu0/div/fdiv/rem2_carry_n_2 ;
  wire \alu0/div/fdiv/rem2_carry_n_3 ;
  wire \alu0/div/fdiv/rem3_carry__0_n_0 ;
  wire \alu0/div/fdiv/rem3_carry__0_n_1 ;
  wire \alu0/div/fdiv/rem3_carry__0_n_2 ;
  wire \alu0/div/fdiv/rem3_carry__0_n_3 ;
  wire \alu0/div/fdiv/rem3_carry__1_n_0 ;
  wire \alu0/div/fdiv/rem3_carry__1_n_1 ;
  wire \alu0/div/fdiv/rem3_carry__1_n_2 ;
  wire \alu0/div/fdiv/rem3_carry__1_n_3 ;
  wire \alu0/div/fdiv/rem3_carry__2_n_0 ;
  wire \alu0/div/fdiv/rem3_carry__2_n_1 ;
  wire \alu0/div/fdiv/rem3_carry__2_n_2 ;
  wire \alu0/div/fdiv/rem3_carry__2_n_3 ;
  wire \alu0/div/fdiv/rem3_carry__3_n_0 ;
  wire \alu0/div/fdiv/rem3_carry__3_n_1 ;
  wire \alu0/div/fdiv/rem3_carry__3_n_2 ;
  wire \alu0/div/fdiv/rem3_carry__3_n_3 ;
  wire \alu0/div/fdiv/rem3_carry__4_n_0 ;
  wire \alu0/div/fdiv/rem3_carry__4_n_1 ;
  wire \alu0/div/fdiv/rem3_carry__4_n_2 ;
  wire \alu0/div/fdiv/rem3_carry__4_n_3 ;
  wire \alu0/div/fdiv/rem3_carry__5_n_0 ;
  wire \alu0/div/fdiv/rem3_carry__5_n_1 ;
  wire \alu0/div/fdiv/rem3_carry__5_n_2 ;
  wire \alu0/div/fdiv/rem3_carry__5_n_3 ;
  wire \alu0/div/fdiv/rem3_carry__6_n_0 ;
  wire \alu0/div/fdiv/rem3_carry__6_n_1 ;
  wire \alu0/div/fdiv/rem3_carry__6_n_2 ;
  wire \alu0/div/fdiv/rem3_carry__6_n_3 ;
  wire \alu0/div/fdiv/rem3_carry_n_0 ;
  wire \alu0/div/fdiv/rem3_carry_n_1 ;
  wire \alu0/div/fdiv/rem3_carry_n_2 ;
  wire \alu0/div/fdiv/rem3_carry_n_3 ;
  wire [31:0]\alu0/div/fdiv_rem ;
  wire \alu0/div/fdiv_rem_msb_f ;
  wire \alu0/div/p_0_in0 ;
  wire [31:0]\alu0/div/p_0_out ;
  wire [31:0]\alu0/div/p_2_in ;
  wire [27:0]\alu0/div/quo ;
  wire [31:28]\alu0/div/quo__0 ;
  wire [31:0]\alu0/div/rem ;
  wire [33:33]\alu0/div/rem1 ;
  wire [32:1]\alu0/div/rem1__0 ;
  wire [33:33]\alu0/div/rem2 ;
  wire [32:1]\alu0/div/rem2__0 ;
  wire [33:33]\alu0/div/rem3 ;
  wire [32:1]\alu0/div/rem3__0 ;
  wire [32:0]\alu0/mul/mul_a ;
  wire \alu0/mul/mul_b ;
  wire \alu0/mul/mul_b_reg_n_0_[0] ;
  wire \alu0/mul/mul_b_reg_n_0_[10] ;
  wire \alu0/mul/mul_b_reg_n_0_[11] ;
  wire \alu0/mul/mul_b_reg_n_0_[12] ;
  wire \alu0/mul/mul_b_reg_n_0_[13] ;
  wire \alu0/mul/mul_b_reg_n_0_[14] ;
  wire \alu0/mul/mul_b_reg_n_0_[15] ;
  wire \alu0/mul/mul_b_reg_n_0_[16] ;
  wire \alu0/mul/mul_b_reg_n_0_[17] ;
  wire \alu0/mul/mul_b_reg_n_0_[18] ;
  wire \alu0/mul/mul_b_reg_n_0_[19] ;
  wire \alu0/mul/mul_b_reg_n_0_[1] ;
  wire \alu0/mul/mul_b_reg_n_0_[20] ;
  wire \alu0/mul/mul_b_reg_n_0_[21] ;
  wire \alu0/mul/mul_b_reg_n_0_[22] ;
  wire \alu0/mul/mul_b_reg_n_0_[23] ;
  wire \alu0/mul/mul_b_reg_n_0_[24] ;
  wire \alu0/mul/mul_b_reg_n_0_[25] ;
  wire \alu0/mul/mul_b_reg_n_0_[26] ;
  wire \alu0/mul/mul_b_reg_n_0_[27] ;
  wire \alu0/mul/mul_b_reg_n_0_[28] ;
  wire \alu0/mul/mul_b_reg_n_0_[29] ;
  wire \alu0/mul/mul_b_reg_n_0_[2] ;
  wire \alu0/mul/mul_b_reg_n_0_[30] ;
  wire \alu0/mul/mul_b_reg_n_0_[31] ;
  wire \alu0/mul/mul_b_reg_n_0_[32] ;
  wire \alu0/mul/mul_b_reg_n_0_[3] ;
  wire \alu0/mul/mul_b_reg_n_0_[4] ;
  wire \alu0/mul/mul_b_reg_n_0_[5] ;
  wire \alu0/mul/mul_b_reg_n_0_[6] ;
  wire \alu0/mul/mul_b_reg_n_0_[7] ;
  wire \alu0/mul/mul_b_reg_n_0_[8] ;
  wire \alu0/mul/mul_b_reg_n_0_[9] ;
  wire \alu0/mul/mul_rslt ;
  wire \alu0/mul/mul_rslt0 ;
  wire [15:0]\alu0/mul/mulh ;
  wire [30:17]\alu0/mul_a_i ;
  wire \alu1/art/add/p_0_in ;
  wire [34:18]\alu1/art/add/tout ;
  wire [32:32]\alu1/art/p_0_in__0 ;
  wire [16:16]\alu1/asr0 ;
  wire [31:0]\alu1/div/add_out ;
  wire \alu1/div/chg_quo_sgn ;
  wire \alu1/div/chg_rem_sgn ;
  wire \alu1/div/dadd/add_out0_carry__0_n_0 ;
  wire \alu1/div/dadd/add_out0_carry__0_n_1 ;
  wire \alu1/div/dadd/add_out0_carry__0_n_2 ;
  wire \alu1/div/dadd/add_out0_carry__0_n_3 ;
  wire \alu1/div/dadd/add_out0_carry__1_n_0 ;
  wire \alu1/div/dadd/add_out0_carry__1_n_1 ;
  wire \alu1/div/dadd/add_out0_carry__1_n_2 ;
  wire \alu1/div/dadd/add_out0_carry__1_n_3 ;
  wire \alu1/div/dadd/add_out0_carry__2_n_0 ;
  wire \alu1/div/dadd/add_out0_carry__2_n_1 ;
  wire \alu1/div/dadd/add_out0_carry__2_n_2 ;
  wire \alu1/div/dadd/add_out0_carry__2_n_3 ;
  wire \alu1/div/dadd/add_out0_carry__3_n_0 ;
  wire \alu1/div/dadd/add_out0_carry__3_n_1 ;
  wire \alu1/div/dadd/add_out0_carry__3_n_2 ;
  wire \alu1/div/dadd/add_out0_carry__3_n_3 ;
  wire \alu1/div/dadd/add_out0_carry__4_n_0 ;
  wire \alu1/div/dadd/add_out0_carry__4_n_1 ;
  wire \alu1/div/dadd/add_out0_carry__4_n_2 ;
  wire \alu1/div/dadd/add_out0_carry__4_n_3 ;
  wire \alu1/div/dadd/add_out0_carry__5_n_0 ;
  wire \alu1/div/dadd/add_out0_carry__5_n_1 ;
  wire \alu1/div/dadd/add_out0_carry__5_n_2 ;
  wire \alu1/div/dadd/add_out0_carry__5_n_3 ;
  wire \alu1/div/dadd/add_out0_carry__6_n_1 ;
  wire \alu1/div/dadd/add_out0_carry__6_n_2 ;
  wire \alu1/div/dadd/add_out0_carry__6_n_3 ;
  wire \alu1/div/dadd/add_out0_carry_n_0 ;
  wire \alu1/div/dadd/add_out0_carry_n_1 ;
  wire \alu1/div/dadd/add_out0_carry_n_2 ;
  wire \alu1/div/dadd/add_out0_carry_n_3 ;
  wire \alu1/div/dctl/dctl_long_f ;
  wire \alu1/div/dctl/dctl_sign ;
  wire \alu1/div/dctl/dctl_sign_f ;
  wire \alu1/div/dctl/fsm/chg_rem_sgn0 ;
  wire [3:0]\alu1/div/dctl/fsm/dctl_next ;
  wire \alu1/div/dctl/fsm/set_sgn ;
  wire \alu1/div/dctl_long ;
  wire [3:0]\alu1/div/dctl_stat ;
  wire [64:0]\alu1/div/den ;
  wire [3:3]\alu1/div/den2 ;
  wire [31:0]\alu1/div/dso_0 ;
  wire [0:0]\alu1/div/fdiv/p_1_in3_in ;
  wire [0:0]\alu1/div/fdiv/p_1_in5_in ;
  wire \alu1/div/fdiv/rem0_carry__0_n_0 ;
  wire \alu1/div/fdiv/rem0_carry__0_n_1 ;
  wire \alu1/div/fdiv/rem0_carry__0_n_2 ;
  wire \alu1/div/fdiv/rem0_carry__0_n_3 ;
  wire \alu1/div/fdiv/rem0_carry__1_n_0 ;
  wire \alu1/div/fdiv/rem0_carry__1_n_1 ;
  wire \alu1/div/fdiv/rem0_carry__1_n_2 ;
  wire \alu1/div/fdiv/rem0_carry__1_n_3 ;
  wire \alu1/div/fdiv/rem0_carry__2_n_0 ;
  wire \alu1/div/fdiv/rem0_carry__2_n_1 ;
  wire \alu1/div/fdiv/rem0_carry__2_n_2 ;
  wire \alu1/div/fdiv/rem0_carry__2_n_3 ;
  wire \alu1/div/fdiv/rem0_carry__3_n_0 ;
  wire \alu1/div/fdiv/rem0_carry__3_n_1 ;
  wire \alu1/div/fdiv/rem0_carry__3_n_2 ;
  wire \alu1/div/fdiv/rem0_carry__3_n_3 ;
  wire \alu1/div/fdiv/rem0_carry__4_n_0 ;
  wire \alu1/div/fdiv/rem0_carry__4_n_1 ;
  wire \alu1/div/fdiv/rem0_carry__4_n_2 ;
  wire \alu1/div/fdiv/rem0_carry__4_n_3 ;
  wire \alu1/div/fdiv/rem0_carry__5_n_0 ;
  wire \alu1/div/fdiv/rem0_carry__5_n_1 ;
  wire \alu1/div/fdiv/rem0_carry__5_n_2 ;
  wire \alu1/div/fdiv/rem0_carry__5_n_3 ;
  wire \alu1/div/fdiv/rem0_carry__6_n_0 ;
  wire \alu1/div/fdiv/rem0_carry__6_n_1 ;
  wire \alu1/div/fdiv/rem0_carry__6_n_2 ;
  wire \alu1/div/fdiv/rem0_carry__6_n_3 ;
  wire \alu1/div/fdiv/rem0_carry_n_0 ;
  wire \alu1/div/fdiv/rem0_carry_n_1 ;
  wire \alu1/div/fdiv/rem0_carry_n_2 ;
  wire \alu1/div/fdiv/rem0_carry_n_3 ;
  wire \alu1/div/fdiv/rem1_carry__0_n_0 ;
  wire \alu1/div/fdiv/rem1_carry__0_n_1 ;
  wire \alu1/div/fdiv/rem1_carry__0_n_2 ;
  wire \alu1/div/fdiv/rem1_carry__0_n_3 ;
  wire \alu1/div/fdiv/rem1_carry__1_n_0 ;
  wire \alu1/div/fdiv/rem1_carry__1_n_1 ;
  wire \alu1/div/fdiv/rem1_carry__1_n_2 ;
  wire \alu1/div/fdiv/rem1_carry__1_n_3 ;
  wire \alu1/div/fdiv/rem1_carry__2_n_0 ;
  wire \alu1/div/fdiv/rem1_carry__2_n_1 ;
  wire \alu1/div/fdiv/rem1_carry__2_n_2 ;
  wire \alu1/div/fdiv/rem1_carry__2_n_3 ;
  wire \alu1/div/fdiv/rem1_carry__3_n_0 ;
  wire \alu1/div/fdiv/rem1_carry__3_n_1 ;
  wire \alu1/div/fdiv/rem1_carry__3_n_2 ;
  wire \alu1/div/fdiv/rem1_carry__3_n_3 ;
  wire \alu1/div/fdiv/rem1_carry__4_n_0 ;
  wire \alu1/div/fdiv/rem1_carry__4_n_1 ;
  wire \alu1/div/fdiv/rem1_carry__4_n_2 ;
  wire \alu1/div/fdiv/rem1_carry__4_n_3 ;
  wire \alu1/div/fdiv/rem1_carry__5_n_0 ;
  wire \alu1/div/fdiv/rem1_carry__5_n_1 ;
  wire \alu1/div/fdiv/rem1_carry__5_n_2 ;
  wire \alu1/div/fdiv/rem1_carry__5_n_3 ;
  wire \alu1/div/fdiv/rem1_carry__6_n_0 ;
  wire \alu1/div/fdiv/rem1_carry__6_n_1 ;
  wire \alu1/div/fdiv/rem1_carry__6_n_2 ;
  wire \alu1/div/fdiv/rem1_carry__6_n_3 ;
  wire \alu1/div/fdiv/rem1_carry_n_0 ;
  wire \alu1/div/fdiv/rem1_carry_n_1 ;
  wire \alu1/div/fdiv/rem1_carry_n_2 ;
  wire \alu1/div/fdiv/rem1_carry_n_3 ;
  wire \alu1/div/fdiv/rem2_carry__0_n_0 ;
  wire \alu1/div/fdiv/rem2_carry__0_n_1 ;
  wire \alu1/div/fdiv/rem2_carry__0_n_2 ;
  wire \alu1/div/fdiv/rem2_carry__0_n_3 ;
  wire \alu1/div/fdiv/rem2_carry__1_n_0 ;
  wire \alu1/div/fdiv/rem2_carry__1_n_1 ;
  wire \alu1/div/fdiv/rem2_carry__1_n_2 ;
  wire \alu1/div/fdiv/rem2_carry__1_n_3 ;
  wire \alu1/div/fdiv/rem2_carry__2_n_0 ;
  wire \alu1/div/fdiv/rem2_carry__2_n_1 ;
  wire \alu1/div/fdiv/rem2_carry__2_n_2 ;
  wire \alu1/div/fdiv/rem2_carry__2_n_3 ;
  wire \alu1/div/fdiv/rem2_carry__3_n_0 ;
  wire \alu1/div/fdiv/rem2_carry__3_n_1 ;
  wire \alu1/div/fdiv/rem2_carry__3_n_2 ;
  wire \alu1/div/fdiv/rem2_carry__3_n_3 ;
  wire \alu1/div/fdiv/rem2_carry__4_n_0 ;
  wire \alu1/div/fdiv/rem2_carry__4_n_1 ;
  wire \alu1/div/fdiv/rem2_carry__4_n_2 ;
  wire \alu1/div/fdiv/rem2_carry__4_n_3 ;
  wire \alu1/div/fdiv/rem2_carry__5_n_0 ;
  wire \alu1/div/fdiv/rem2_carry__5_n_1 ;
  wire \alu1/div/fdiv/rem2_carry__5_n_2 ;
  wire \alu1/div/fdiv/rem2_carry__5_n_3 ;
  wire \alu1/div/fdiv/rem2_carry__6_n_0 ;
  wire \alu1/div/fdiv/rem2_carry__6_n_1 ;
  wire \alu1/div/fdiv/rem2_carry__6_n_2 ;
  wire \alu1/div/fdiv/rem2_carry__6_n_3 ;
  wire \alu1/div/fdiv/rem2_carry_n_0 ;
  wire \alu1/div/fdiv/rem2_carry_n_1 ;
  wire \alu1/div/fdiv/rem2_carry_n_2 ;
  wire \alu1/div/fdiv/rem2_carry_n_3 ;
  wire \alu1/div/fdiv/rem3_carry__0_n_0 ;
  wire \alu1/div/fdiv/rem3_carry__0_n_1 ;
  wire \alu1/div/fdiv/rem3_carry__0_n_2 ;
  wire \alu1/div/fdiv/rem3_carry__0_n_3 ;
  wire \alu1/div/fdiv/rem3_carry__1_n_0 ;
  wire \alu1/div/fdiv/rem3_carry__1_n_1 ;
  wire \alu1/div/fdiv/rem3_carry__1_n_2 ;
  wire \alu1/div/fdiv/rem3_carry__1_n_3 ;
  wire \alu1/div/fdiv/rem3_carry__2_n_0 ;
  wire \alu1/div/fdiv/rem3_carry__2_n_1 ;
  wire \alu1/div/fdiv/rem3_carry__2_n_2 ;
  wire \alu1/div/fdiv/rem3_carry__2_n_3 ;
  wire \alu1/div/fdiv/rem3_carry__3_n_0 ;
  wire \alu1/div/fdiv/rem3_carry__3_n_1 ;
  wire \alu1/div/fdiv/rem3_carry__3_n_2 ;
  wire \alu1/div/fdiv/rem3_carry__3_n_3 ;
  wire \alu1/div/fdiv/rem3_carry__4_n_0 ;
  wire \alu1/div/fdiv/rem3_carry__4_n_1 ;
  wire \alu1/div/fdiv/rem3_carry__4_n_2 ;
  wire \alu1/div/fdiv/rem3_carry__4_n_3 ;
  wire \alu1/div/fdiv/rem3_carry__5_n_0 ;
  wire \alu1/div/fdiv/rem3_carry__5_n_1 ;
  wire \alu1/div/fdiv/rem3_carry__5_n_2 ;
  wire \alu1/div/fdiv/rem3_carry__5_n_3 ;
  wire \alu1/div/fdiv/rem3_carry__6_n_0 ;
  wire \alu1/div/fdiv/rem3_carry__6_n_1 ;
  wire \alu1/div/fdiv/rem3_carry__6_n_2 ;
  wire \alu1/div/fdiv/rem3_carry__6_n_3 ;
  wire \alu1/div/fdiv/rem3_carry_n_0 ;
  wire \alu1/div/fdiv/rem3_carry_n_1 ;
  wire \alu1/div/fdiv/rem3_carry_n_2 ;
  wire \alu1/div/fdiv/rem3_carry_n_3 ;
  wire [31:0]\alu1/div/fdiv_rem ;
  wire \alu1/div/fdiv_rem_msb_f ;
  wire \alu1/div/p_0_in0 ;
  wire \alu1/div/p_0_in__0 ;
  wire [31:0]\alu1/div/p_0_out ;
  wire [31:0]\alu1/div/p_2_in ;
  wire [27:0]\alu1/div/quo ;
  wire [31:28]\alu1/div/quo__0 ;
  wire [31:0]\alu1/div/rem ;
  wire [33:33]\alu1/div/rem1 ;
  wire [32:1]\alu1/div/rem1__0 ;
  wire [33:33]\alu1/div/rem2 ;
  wire [32:1]\alu1/div/rem2__0 ;
  wire [33:33]\alu1/div/rem3 ;
  wire [32:1]\alu1/div/rem3__0 ;
  wire [32:0]\alu1/mul/mul_a ;
  wire \alu1/mul/mul_b ;
  wire \alu1/mul/mul_b_reg_n_0_[0] ;
  wire \alu1/mul/mul_b_reg_n_0_[10] ;
  wire \alu1/mul/mul_b_reg_n_0_[11] ;
  wire \alu1/mul/mul_b_reg_n_0_[12] ;
  wire \alu1/mul/mul_b_reg_n_0_[13] ;
  wire \alu1/mul/mul_b_reg_n_0_[14] ;
  wire \alu1/mul/mul_b_reg_n_0_[15] ;
  wire \alu1/mul/mul_b_reg_n_0_[16] ;
  wire \alu1/mul/mul_b_reg_n_0_[17] ;
  wire \alu1/mul/mul_b_reg_n_0_[18] ;
  wire \alu1/mul/mul_b_reg_n_0_[19] ;
  wire \alu1/mul/mul_b_reg_n_0_[1] ;
  wire \alu1/mul/mul_b_reg_n_0_[20] ;
  wire \alu1/mul/mul_b_reg_n_0_[21] ;
  wire \alu1/mul/mul_b_reg_n_0_[22] ;
  wire \alu1/mul/mul_b_reg_n_0_[23] ;
  wire \alu1/mul/mul_b_reg_n_0_[24] ;
  wire \alu1/mul/mul_b_reg_n_0_[25] ;
  wire \alu1/mul/mul_b_reg_n_0_[26] ;
  wire \alu1/mul/mul_b_reg_n_0_[27] ;
  wire \alu1/mul/mul_b_reg_n_0_[28] ;
  wire \alu1/mul/mul_b_reg_n_0_[29] ;
  wire \alu1/mul/mul_b_reg_n_0_[2] ;
  wire \alu1/mul/mul_b_reg_n_0_[30] ;
  wire \alu1/mul/mul_b_reg_n_0_[31] ;
  wire \alu1/mul/mul_b_reg_n_0_[32] ;
  wire \alu1/mul/mul_b_reg_n_0_[3] ;
  wire \alu1/mul/mul_b_reg_n_0_[4] ;
  wire \alu1/mul/mul_b_reg_n_0_[5] ;
  wire \alu1/mul/mul_b_reg_n_0_[6] ;
  wire \alu1/mul/mul_b_reg_n_0_[7] ;
  wire \alu1/mul/mul_b_reg_n_0_[8] ;
  wire \alu1/mul/mul_b_reg_n_0_[9] ;
  wire \alu1/mul/mul_rslt ;
  wire \alu1/mul/mul_rslt0 ;
  wire [15:0]\alu1/mul/mulh ;
  wire [31:17]\alu1/mul_a_i ;
  wire [1:0]alu_sr_flag0;
  wire [3:0]alu_sr_flag1;
  wire \art/add/rgf_c0bus_wb[11]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[11]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[11]_i_31_n_0 ;
  wire \art/add/rgf_c0bus_wb[11]_i_32_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_31_n_0 ;
  wire \art/add/rgf_c0bus_wb[15]_i_32_n_0 ;
  wire \art/add/rgf_c0bus_wb[19]_i_28_n_0 ;
  wire \art/add/rgf_c0bus_wb[19]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[19]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[23]_i_38_n_0 ;
  wire \art/add/rgf_c0bus_wb[23]_i_39_n_0 ;
  wire \art/add/rgf_c0bus_wb[27]_i_40_n_0 ;
  wire \art/add/rgf_c0bus_wb[27]_i_41_n_0 ;
  wire \art/add/rgf_c0bus_wb[29]_i_29_n_0 ;
  wire \art/add/rgf_c0bus_wb[29]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_23_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_24_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_25_n_0 ;
  wire \art/add/rgf_c0bus_wb[3]_i_26_n_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_30_n_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_31_n_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_32_n_0 ;
  wire \art/add/rgf_c0bus_wb[7]_i_33_n_0 ;
  wire \art/add/rgf_c1bus_wb[11]_i_26_n_0 ;
  wire \art/add/rgf_c1bus_wb[11]_i_27_n_0 ;
  wire \art/add/rgf_c1bus_wb[11]_i_28_n_0 ;
  wire \art/add/rgf_c1bus_wb[11]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_23_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_24_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_25_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_26_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_35_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_36_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_37_n_0 ;
  wire \art/add/rgf_c1bus_wb[19]_i_38_n_0 ;
  wire \art/add/rgf_c1bus_wb[23]_i_27_n_0 ;
  wire \art/add/rgf_c1bus_wb[23]_i_28_n_0 ;
  wire \art/add/rgf_c1bus_wb[23]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_21_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_22_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_23_n_0 ;
  wire \art/add/rgf_c1bus_wb[27]_i_24_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_30_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_31_n_0 ;
  wire \art/add/rgf_c1bus_wb[31]_i_32_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_27_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_28_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_29_n_0 ;
  wire \art/add/rgf_c1bus_wb[3]_i_30_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_31_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_32_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_33_n_0 ;
  wire \art/add/rgf_c1bus_wb[7]_i_34_n_0 ;
  wire \art/add/sr[6]_i_29_n_0 ;
  wire [31:0]b0bus_0;
  wire [31:0]b1bus_0;
  wire [31:0]badr;
  wire \badr[0]_INST_0_i_25_n_0 ;
  wire \badr[0]_INST_0_i_3_n_0 ;
  wire \badr[0]_INST_0_i_44_n_0 ;
  wire \badr[0]_INST_0_i_45_n_0 ;
  wire \badr[0]_INST_0_i_46_n_0 ;
  wire \badr[0]_INST_0_i_47_n_0 ;
  wire \badr[0]_INST_0_i_7_n_0 ;
  wire \badr[10]_INST_0_i_17_n_0 ;
  wire \badr[10]_INST_0_i_21_n_0 ;
  wire \badr[10]_INST_0_i_3_n_0 ;
  wire \badr[10]_INST_0_i_45_n_0 ;
  wire \badr[10]_INST_0_i_46_n_0 ;
  wire \badr[10]_INST_0_i_47_n_0 ;
  wire \badr[10]_INST_0_i_48_n_0 ;
  wire \badr[10]_INST_0_i_9_n_0 ;
  wire \badr[11]_INST_0_i_17_n_0 ;
  wire \badr[11]_INST_0_i_21_n_0 ;
  wire \badr[11]_INST_0_i_3_n_0 ;
  wire \badr[11]_INST_0_i_45_n_0 ;
  wire \badr[11]_INST_0_i_46_n_0 ;
  wire \badr[11]_INST_0_i_47_n_0 ;
  wire \badr[11]_INST_0_i_48_n_0 ;
  wire \badr[11]_INST_0_i_9_n_0 ;
  wire \badr[12]_INST_0_i_17_n_0 ;
  wire \badr[12]_INST_0_i_21_n_0 ;
  wire \badr[12]_INST_0_i_29_n_0 ;
  wire \badr[12]_INST_0_i_29_n_1 ;
  wire \badr[12]_INST_0_i_29_n_2 ;
  wire \badr[12]_INST_0_i_29_n_3 ;
  wire \badr[12]_INST_0_i_3_n_0 ;
  wire \badr[12]_INST_0_i_46_n_0 ;
  wire \badr[12]_INST_0_i_47_n_0 ;
  wire \badr[12]_INST_0_i_48_n_0 ;
  wire \badr[12]_INST_0_i_49_n_0 ;
  wire \badr[12]_INST_0_i_50_n_0 ;
  wire \badr[12]_INST_0_i_51_n_0 ;
  wire \badr[12]_INST_0_i_52_n_0 ;
  wire \badr[12]_INST_0_i_53_n_0 ;
  wire \badr[12]_INST_0_i_9_n_0 ;
  wire \badr[13]_INST_0_i_15_n_0 ;
  wire \badr[13]_INST_0_i_19_n_0 ;
  wire \badr[13]_INST_0_i_24_n_0 ;
  wire \badr[13]_INST_0_i_3_n_0 ;
  wire \badr[13]_INST_0_i_46_n_0 ;
  wire \badr[13]_INST_0_i_49_n_0 ;
  wire \badr[13]_INST_0_i_50_n_0 ;
  wire \badr[13]_INST_0_i_51_n_0 ;
  wire \badr[13]_INST_0_i_52_n_0 ;
  wire \badr[13]_INST_0_i_9_n_0 ;
  wire \badr[14]_INST_0_i_43_n_0 ;
  wire \badr[14]_INST_0_i_44_n_0 ;
  wire \badr[14]_INST_0_i_45_n_0 ;
  wire \badr[14]_INST_0_i_46_n_0 ;
  wire \badr[14]_INST_0_i_7_n_0 ;
  wire \badr[15]_INST_0_i_100_n_0 ;
  wire \badr[15]_INST_0_i_103_n_0 ;
  wire \badr[15]_INST_0_i_104_n_0 ;
  wire \badr[15]_INST_0_i_113_n_0 ;
  wire \badr[15]_INST_0_i_114_n_0 ;
  wire \badr[15]_INST_0_i_115_n_0 ;
  wire \badr[15]_INST_0_i_116_n_0 ;
  wire \badr[15]_INST_0_i_117_n_0 ;
  wire \badr[15]_INST_0_i_118_n_0 ;
  wire \badr[15]_INST_0_i_119_n_0 ;
  wire \badr[15]_INST_0_i_120_n_0 ;
  wire \badr[15]_INST_0_i_121_n_0 ;
  wire \badr[15]_INST_0_i_122_n_0 ;
  wire \badr[15]_INST_0_i_123_n_0 ;
  wire \badr[15]_INST_0_i_124_n_0 ;
  wire \badr[15]_INST_0_i_125_n_0 ;
  wire \badr[15]_INST_0_i_126_n_0 ;
  wire \badr[15]_INST_0_i_127_n_0 ;
  wire \badr[15]_INST_0_i_128_n_0 ;
  wire \badr[15]_INST_0_i_129_n_0 ;
  wire \badr[15]_INST_0_i_131_n_0 ;
  wire \badr[15]_INST_0_i_132_n_0 ;
  wire \badr[15]_INST_0_i_133_n_0 ;
  wire \badr[15]_INST_0_i_134_n_0 ;
  wire \badr[15]_INST_0_i_135_n_0 ;
  wire \badr[15]_INST_0_i_136_n_0 ;
  wire \badr[15]_INST_0_i_137_n_0 ;
  wire \badr[15]_INST_0_i_138_n_0 ;
  wire \badr[15]_INST_0_i_139_n_0 ;
  wire \badr[15]_INST_0_i_140_n_0 ;
  wire \badr[15]_INST_0_i_141_n_0 ;
  wire \badr[15]_INST_0_i_142_n_0 ;
  wire \badr[15]_INST_0_i_143_n_0 ;
  wire \badr[15]_INST_0_i_144_n_0 ;
  wire \badr[15]_INST_0_i_145_n_0 ;
  wire \badr[15]_INST_0_i_146_n_0 ;
  wire \badr[15]_INST_0_i_147_n_0 ;
  wire \badr[15]_INST_0_i_148_n_0 ;
  wire \badr[15]_INST_0_i_149_n_0 ;
  wire \badr[15]_INST_0_i_14_n_0 ;
  wire \badr[15]_INST_0_i_150_n_0 ;
  wire \badr[15]_INST_0_i_151_n_0 ;
  wire \badr[15]_INST_0_i_15_n_0 ;
  wire \badr[15]_INST_0_i_29_n_0 ;
  wire \badr[15]_INST_0_i_47_n_0 ;
  wire \badr[15]_INST_0_i_48_n_0 ;
  wire \badr[15]_INST_0_i_49_n_0 ;
  wire \badr[15]_INST_0_i_50_n_0 ;
  wire \badr[15]_INST_0_i_51_n_0 ;
  wire \badr[15]_INST_0_i_52_n_0 ;
  wire \badr[15]_INST_0_i_8_n_0 ;
  wire \badr[15]_INST_0_i_99_n_0 ;
  wire \badr[16]_INST_0_i_15_n_0 ;
  wire \badr[16]_INST_0_i_16_n_0 ;
  wire \badr[16]_INST_0_i_18_n_0 ;
  wire \badr[16]_INST_0_i_19_n_0 ;
  wire \badr[16]_INST_0_i_21_n_0 ;
  wire \badr[16]_INST_0_i_21_n_1 ;
  wire \badr[16]_INST_0_i_21_n_2 ;
  wire \badr[16]_INST_0_i_21_n_3 ;
  wire \badr[16]_INST_0_i_22_n_0 ;
  wire \badr[16]_INST_0_i_23_n_0 ;
  wire \badr[16]_INST_0_i_24_n_0 ;
  wire \badr[16]_INST_0_i_25_n_0 ;
  wire \badr[16]_INST_0_i_26_n_0 ;
  wire \badr[16]_INST_0_i_27_n_0 ;
  wire \badr[16]_INST_0_i_28_n_0 ;
  wire \badr[16]_INST_0_i_29_n_0 ;
  wire \badr[16]_INST_0_i_30_n_0 ;
  wire \badr[16]_INST_0_i_31_n_0 ;
  wire \badr[16]_INST_0_i_32_n_0 ;
  wire \badr[16]_INST_0_i_33_n_0 ;
  wire \badr[16]_INST_0_i_3_n_0 ;
  wire \badr[16]_INST_0_i_9_n_0 ;
  wire \badr[17]_INST_0_i_15_n_0 ;
  wire \badr[17]_INST_0_i_16_n_0 ;
  wire \badr[17]_INST_0_i_18_n_0 ;
  wire \badr[17]_INST_0_i_19_n_0 ;
  wire \badr[17]_INST_0_i_21_n_0 ;
  wire \badr[17]_INST_0_i_22_n_0 ;
  wire \badr[17]_INST_0_i_23_n_0 ;
  wire \badr[17]_INST_0_i_24_n_0 ;
  wire \badr[17]_INST_0_i_25_n_0 ;
  wire \badr[17]_INST_0_i_26_n_0 ;
  wire \badr[17]_INST_0_i_27_n_0 ;
  wire \badr[17]_INST_0_i_28_n_0 ;
  wire \badr[17]_INST_0_i_3_n_0 ;
  wire \badr[17]_INST_0_i_9_n_0 ;
  wire \badr[18]_INST_0_i_15_n_0 ;
  wire \badr[18]_INST_0_i_16_n_0 ;
  wire \badr[18]_INST_0_i_18_n_0 ;
  wire \badr[18]_INST_0_i_19_n_0 ;
  wire \badr[18]_INST_0_i_21_n_0 ;
  wire \badr[18]_INST_0_i_22_n_0 ;
  wire \badr[18]_INST_0_i_23_n_0 ;
  wire \badr[18]_INST_0_i_24_n_0 ;
  wire \badr[18]_INST_0_i_25_n_0 ;
  wire \badr[18]_INST_0_i_26_n_0 ;
  wire \badr[18]_INST_0_i_27_n_0 ;
  wire \badr[18]_INST_0_i_28_n_0 ;
  wire \badr[18]_INST_0_i_3_n_0 ;
  wire \badr[18]_INST_0_i_9_n_0 ;
  wire \badr[19]_INST_0_i_15_n_0 ;
  wire \badr[19]_INST_0_i_16_n_0 ;
  wire \badr[19]_INST_0_i_18_n_0 ;
  wire \badr[19]_INST_0_i_19_n_0 ;
  wire \badr[19]_INST_0_i_21_n_0 ;
  wire \badr[19]_INST_0_i_22_n_0 ;
  wire \badr[19]_INST_0_i_23_n_0 ;
  wire \badr[19]_INST_0_i_24_n_0 ;
  wire \badr[19]_INST_0_i_25_n_0 ;
  wire \badr[19]_INST_0_i_26_n_0 ;
  wire \badr[19]_INST_0_i_27_n_0 ;
  wire \badr[19]_INST_0_i_28_n_0 ;
  wire \badr[19]_INST_0_i_3_n_0 ;
  wire \badr[19]_INST_0_i_9_n_0 ;
  wire \badr[1]_INST_0_i_43_n_0 ;
  wire \badr[1]_INST_0_i_44_n_0 ;
  wire \badr[1]_INST_0_i_45_n_0 ;
  wire \badr[1]_INST_0_i_46_n_0 ;
  wire \badr[1]_INST_0_i_7_n_0 ;
  wire \badr[20]_INST_0_i_15_n_0 ;
  wire \badr[20]_INST_0_i_16_n_0 ;
  wire \badr[20]_INST_0_i_18_n_0 ;
  wire \badr[20]_INST_0_i_19_n_0 ;
  wire \badr[20]_INST_0_i_21_n_0 ;
  wire \badr[20]_INST_0_i_21_n_1 ;
  wire \badr[20]_INST_0_i_21_n_2 ;
  wire \badr[20]_INST_0_i_21_n_3 ;
  wire \badr[20]_INST_0_i_22_n_0 ;
  wire \badr[20]_INST_0_i_23_n_0 ;
  wire \badr[20]_INST_0_i_24_n_0 ;
  wire \badr[20]_INST_0_i_25_n_0 ;
  wire \badr[20]_INST_0_i_26_n_0 ;
  wire \badr[20]_INST_0_i_27_n_0 ;
  wire \badr[20]_INST_0_i_28_n_0 ;
  wire \badr[20]_INST_0_i_29_n_0 ;
  wire \badr[20]_INST_0_i_30_n_0 ;
  wire \badr[20]_INST_0_i_31_n_0 ;
  wire \badr[20]_INST_0_i_32_n_0 ;
  wire \badr[20]_INST_0_i_33_n_0 ;
  wire \badr[20]_INST_0_i_3_n_0 ;
  wire \badr[20]_INST_0_i_9_n_0 ;
  wire \badr[21]_INST_0_i_15_n_0 ;
  wire \badr[21]_INST_0_i_16_n_0 ;
  wire \badr[21]_INST_0_i_18_n_0 ;
  wire \badr[21]_INST_0_i_19_n_0 ;
  wire \badr[21]_INST_0_i_21_n_0 ;
  wire \badr[21]_INST_0_i_22_n_0 ;
  wire \badr[21]_INST_0_i_23_n_0 ;
  wire \badr[21]_INST_0_i_24_n_0 ;
  wire \badr[21]_INST_0_i_25_n_0 ;
  wire \badr[21]_INST_0_i_26_n_0 ;
  wire \badr[21]_INST_0_i_27_n_0 ;
  wire \badr[21]_INST_0_i_28_n_0 ;
  wire \badr[21]_INST_0_i_3_n_0 ;
  wire \badr[21]_INST_0_i_9_n_0 ;
  wire \badr[22]_INST_0_i_15_n_0 ;
  wire \badr[22]_INST_0_i_16_n_0 ;
  wire \badr[22]_INST_0_i_18_n_0 ;
  wire \badr[22]_INST_0_i_19_n_0 ;
  wire \badr[22]_INST_0_i_21_n_0 ;
  wire \badr[22]_INST_0_i_22_n_0 ;
  wire \badr[22]_INST_0_i_23_n_0 ;
  wire \badr[22]_INST_0_i_24_n_0 ;
  wire \badr[22]_INST_0_i_25_n_0 ;
  wire \badr[22]_INST_0_i_26_n_0 ;
  wire \badr[22]_INST_0_i_27_n_0 ;
  wire \badr[22]_INST_0_i_28_n_0 ;
  wire \badr[22]_INST_0_i_3_n_0 ;
  wire \badr[22]_INST_0_i_9_n_0 ;
  wire \badr[23]_INST_0_i_15_n_0 ;
  wire \badr[23]_INST_0_i_16_n_0 ;
  wire \badr[23]_INST_0_i_18_n_0 ;
  wire \badr[23]_INST_0_i_19_n_0 ;
  wire \badr[23]_INST_0_i_21_n_0 ;
  wire \badr[23]_INST_0_i_22_n_0 ;
  wire \badr[23]_INST_0_i_23_n_0 ;
  wire \badr[23]_INST_0_i_24_n_0 ;
  wire \badr[23]_INST_0_i_25_n_0 ;
  wire \badr[23]_INST_0_i_26_n_0 ;
  wire \badr[23]_INST_0_i_27_n_0 ;
  wire \badr[23]_INST_0_i_28_n_0 ;
  wire \badr[23]_INST_0_i_3_n_0 ;
  wire \badr[23]_INST_0_i_9_n_0 ;
  wire \badr[24]_INST_0_i_15_n_0 ;
  wire \badr[24]_INST_0_i_16_n_0 ;
  wire \badr[24]_INST_0_i_18_n_0 ;
  wire \badr[24]_INST_0_i_19_n_0 ;
  wire \badr[24]_INST_0_i_21_n_0 ;
  wire \badr[24]_INST_0_i_21_n_1 ;
  wire \badr[24]_INST_0_i_21_n_2 ;
  wire \badr[24]_INST_0_i_21_n_3 ;
  wire \badr[24]_INST_0_i_22_n_0 ;
  wire \badr[24]_INST_0_i_23_n_0 ;
  wire \badr[24]_INST_0_i_24_n_0 ;
  wire \badr[24]_INST_0_i_25_n_0 ;
  wire \badr[24]_INST_0_i_26_n_0 ;
  wire \badr[24]_INST_0_i_27_n_0 ;
  wire \badr[24]_INST_0_i_28_n_0 ;
  wire \badr[24]_INST_0_i_29_n_0 ;
  wire \badr[24]_INST_0_i_30_n_0 ;
  wire \badr[24]_INST_0_i_31_n_0 ;
  wire \badr[24]_INST_0_i_32_n_0 ;
  wire \badr[24]_INST_0_i_33_n_0 ;
  wire \badr[24]_INST_0_i_3_n_0 ;
  wire \badr[24]_INST_0_i_9_n_0 ;
  wire \badr[25]_INST_0_i_15_n_0 ;
  wire \badr[25]_INST_0_i_16_n_0 ;
  wire \badr[25]_INST_0_i_18_n_0 ;
  wire \badr[25]_INST_0_i_19_n_0 ;
  wire \badr[25]_INST_0_i_21_n_0 ;
  wire \badr[25]_INST_0_i_22_n_0 ;
  wire \badr[25]_INST_0_i_23_n_0 ;
  wire \badr[25]_INST_0_i_24_n_0 ;
  wire \badr[25]_INST_0_i_25_n_0 ;
  wire \badr[25]_INST_0_i_26_n_0 ;
  wire \badr[25]_INST_0_i_27_n_0 ;
  wire \badr[25]_INST_0_i_28_n_0 ;
  wire \badr[25]_INST_0_i_3_n_0 ;
  wire \badr[25]_INST_0_i_9_n_0 ;
  wire \badr[26]_INST_0_i_15_n_0 ;
  wire \badr[26]_INST_0_i_16_n_0 ;
  wire \badr[26]_INST_0_i_18_n_0 ;
  wire \badr[26]_INST_0_i_19_n_0 ;
  wire \badr[26]_INST_0_i_21_n_0 ;
  wire \badr[26]_INST_0_i_22_n_0 ;
  wire \badr[26]_INST_0_i_23_n_0 ;
  wire \badr[26]_INST_0_i_24_n_0 ;
  wire \badr[26]_INST_0_i_25_n_0 ;
  wire \badr[26]_INST_0_i_26_n_0 ;
  wire \badr[26]_INST_0_i_27_n_0 ;
  wire \badr[26]_INST_0_i_28_n_0 ;
  wire \badr[26]_INST_0_i_3_n_0 ;
  wire \badr[26]_INST_0_i_9_n_0 ;
  wire \badr[27]_INST_0_i_15_n_0 ;
  wire \badr[27]_INST_0_i_16_n_0 ;
  wire \badr[27]_INST_0_i_18_n_0 ;
  wire \badr[27]_INST_0_i_19_n_0 ;
  wire \badr[27]_INST_0_i_21_n_0 ;
  wire \badr[27]_INST_0_i_22_n_0 ;
  wire \badr[27]_INST_0_i_23_n_0 ;
  wire \badr[27]_INST_0_i_24_n_0 ;
  wire \badr[27]_INST_0_i_25_n_0 ;
  wire \badr[27]_INST_0_i_26_n_0 ;
  wire \badr[27]_INST_0_i_27_n_0 ;
  wire \badr[27]_INST_0_i_28_n_0 ;
  wire \badr[27]_INST_0_i_3_n_0 ;
  wire \badr[27]_INST_0_i_9_n_0 ;
  wire \badr[28]_INST_0_i_15_n_0 ;
  wire \badr[28]_INST_0_i_16_n_0 ;
  wire \badr[28]_INST_0_i_18_n_0 ;
  wire \badr[28]_INST_0_i_19_n_0 ;
  wire \badr[28]_INST_0_i_21_n_0 ;
  wire \badr[28]_INST_0_i_21_n_1 ;
  wire \badr[28]_INST_0_i_21_n_2 ;
  wire \badr[28]_INST_0_i_21_n_3 ;
  wire \badr[28]_INST_0_i_22_n_0 ;
  wire \badr[28]_INST_0_i_23_n_0 ;
  wire \badr[28]_INST_0_i_24_n_0 ;
  wire \badr[28]_INST_0_i_25_n_0 ;
  wire \badr[28]_INST_0_i_26_n_0 ;
  wire \badr[28]_INST_0_i_27_n_0 ;
  wire \badr[28]_INST_0_i_28_n_0 ;
  wire \badr[28]_INST_0_i_29_n_0 ;
  wire \badr[28]_INST_0_i_30_n_0 ;
  wire \badr[28]_INST_0_i_31_n_0 ;
  wire \badr[28]_INST_0_i_32_n_0 ;
  wire \badr[28]_INST_0_i_33_n_0 ;
  wire \badr[28]_INST_0_i_3_n_0 ;
  wire \badr[28]_INST_0_i_9_n_0 ;
  wire \badr[29]_INST_0_i_15_n_0 ;
  wire \badr[29]_INST_0_i_16_n_0 ;
  wire \badr[29]_INST_0_i_18_n_0 ;
  wire \badr[29]_INST_0_i_19_n_0 ;
  wire \badr[29]_INST_0_i_21_n_0 ;
  wire \badr[29]_INST_0_i_22_n_0 ;
  wire \badr[29]_INST_0_i_23_n_0 ;
  wire \badr[29]_INST_0_i_24_n_0 ;
  wire \badr[29]_INST_0_i_25_n_0 ;
  wire \badr[29]_INST_0_i_26_n_0 ;
  wire \badr[29]_INST_0_i_27_n_0 ;
  wire \badr[29]_INST_0_i_28_n_0 ;
  wire \badr[29]_INST_0_i_3_n_0 ;
  wire \badr[29]_INST_0_i_9_n_0 ;
  wire \badr[2]_INST_0_i_43_n_0 ;
  wire \badr[2]_INST_0_i_44_n_0 ;
  wire \badr[2]_INST_0_i_45_n_0 ;
  wire \badr[2]_INST_0_i_46_n_0 ;
  wire \badr[2]_INST_0_i_7_n_0 ;
  wire \badr[30]_INST_0_i_15_n_0 ;
  wire \badr[30]_INST_0_i_16_n_0 ;
  wire \badr[30]_INST_0_i_18_n_0 ;
  wire \badr[30]_INST_0_i_19_n_0 ;
  wire \badr[30]_INST_0_i_21_n_0 ;
  wire \badr[30]_INST_0_i_22_n_0 ;
  wire \badr[30]_INST_0_i_23_n_0 ;
  wire \badr[30]_INST_0_i_24_n_0 ;
  wire \badr[30]_INST_0_i_25_n_0 ;
  wire \badr[30]_INST_0_i_26_n_0 ;
  wire \badr[30]_INST_0_i_27_n_0 ;
  wire \badr[30]_INST_0_i_28_n_0 ;
  wire \badr[30]_INST_0_i_3_n_0 ;
  wire \badr[30]_INST_0_i_9_n_0 ;
  wire \badr[31]_INST_0_i_100_n_0 ;
  wire \badr[31]_INST_0_i_101_n_0 ;
  wire \badr[31]_INST_0_i_102_n_0 ;
  wire \badr[31]_INST_0_i_103_n_0 ;
  wire \badr[31]_INST_0_i_104_n_0 ;
  wire \badr[31]_INST_0_i_105_n_0 ;
  wire \badr[31]_INST_0_i_106_n_0 ;
  wire \badr[31]_INST_0_i_107_n_0 ;
  wire \badr[31]_INST_0_i_108_n_0 ;
  wire \badr[31]_INST_0_i_109_n_0 ;
  wire \badr[31]_INST_0_i_110_n_0 ;
  wire \badr[31]_INST_0_i_111_n_0 ;
  wire \badr[31]_INST_0_i_112_n_0 ;
  wire \badr[31]_INST_0_i_113_n_0 ;
  wire \badr[31]_INST_0_i_114_n_0 ;
  wire \badr[31]_INST_0_i_115_n_0 ;
  wire \badr[31]_INST_0_i_116_n_0 ;
  wire \badr[31]_INST_0_i_117_n_0 ;
  wire \badr[31]_INST_0_i_118_n_0 ;
  wire \badr[31]_INST_0_i_119_n_0 ;
  wire \badr[31]_INST_0_i_11_n_0 ;
  wire \badr[31]_INST_0_i_120_n_0 ;
  wire \badr[31]_INST_0_i_121_n_0 ;
  wire \badr[31]_INST_0_i_122_n_0 ;
  wire \badr[31]_INST_0_i_123_n_0 ;
  wire \badr[31]_INST_0_i_124_n_0 ;
  wire \badr[31]_INST_0_i_125_n_0 ;
  wire \badr[31]_INST_0_i_126_n_0 ;
  wire \badr[31]_INST_0_i_127_n_0 ;
  wire \badr[31]_INST_0_i_128_n_0 ;
  wire \badr[31]_INST_0_i_129_n_0 ;
  wire \badr[31]_INST_0_i_130_n_0 ;
  wire \badr[31]_INST_0_i_131_n_0 ;
  wire \badr[31]_INST_0_i_132_n_0 ;
  wire \badr[31]_INST_0_i_133_n_0 ;
  wire \badr[31]_INST_0_i_134_n_0 ;
  wire \badr[31]_INST_0_i_135_n_0 ;
  wire \badr[31]_INST_0_i_136_n_0 ;
  wire \badr[31]_INST_0_i_137_n_0 ;
  wire \badr[31]_INST_0_i_138_n_0 ;
  wire \badr[31]_INST_0_i_139_n_0 ;
  wire \badr[31]_INST_0_i_140_n_0 ;
  wire \badr[31]_INST_0_i_141_n_0 ;
  wire \badr[31]_INST_0_i_142_n_0 ;
  wire \badr[31]_INST_0_i_143_n_0 ;
  wire \badr[31]_INST_0_i_144_n_0 ;
  wire \badr[31]_INST_0_i_145_n_0 ;
  wire \badr[31]_INST_0_i_146_n_0 ;
  wire \badr[31]_INST_0_i_147_n_0 ;
  wire \badr[31]_INST_0_i_148_n_0 ;
  wire \badr[31]_INST_0_i_149_n_0 ;
  wire \badr[31]_INST_0_i_150_n_0 ;
  wire \badr[31]_INST_0_i_151_n_0 ;
  wire \badr[31]_INST_0_i_152_n_0 ;
  wire \badr[31]_INST_0_i_153_n_0 ;
  wire \badr[31]_INST_0_i_154_n_0 ;
  wire \badr[31]_INST_0_i_155_n_0 ;
  wire \badr[31]_INST_0_i_156_n_0 ;
  wire \badr[31]_INST_0_i_157_n_0 ;
  wire \badr[31]_INST_0_i_158_n_0 ;
  wire \badr[31]_INST_0_i_159_n_0 ;
  wire \badr[31]_INST_0_i_160_n_0 ;
  wire \badr[31]_INST_0_i_161_n_0 ;
  wire \badr[31]_INST_0_i_162_n_0 ;
  wire \badr[31]_INST_0_i_163_n_0 ;
  wire \badr[31]_INST_0_i_164_n_0 ;
  wire \badr[31]_INST_0_i_165_n_0 ;
  wire \badr[31]_INST_0_i_166_n_0 ;
  wire \badr[31]_INST_0_i_167_n_0 ;
  wire \badr[31]_INST_0_i_168_n_0 ;
  wire \badr[31]_INST_0_i_169_n_0 ;
  wire \badr[31]_INST_0_i_170_n_0 ;
  wire \badr[31]_INST_0_i_171_n_0 ;
  wire \badr[31]_INST_0_i_172_n_0 ;
  wire \badr[31]_INST_0_i_173_n_0 ;
  wire \badr[31]_INST_0_i_174_n_0 ;
  wire \badr[31]_INST_0_i_175_n_0 ;
  wire \badr[31]_INST_0_i_176_n_0 ;
  wire \badr[31]_INST_0_i_177_n_0 ;
  wire \badr[31]_INST_0_i_178_n_0 ;
  wire \badr[31]_INST_0_i_179_n_0 ;
  wire \badr[31]_INST_0_i_17_n_0 ;
  wire \badr[31]_INST_0_i_180_n_0 ;
  wire \badr[31]_INST_0_i_181_n_0 ;
  wire \badr[31]_INST_0_i_182_n_0 ;
  wire \badr[31]_INST_0_i_183_n_0 ;
  wire \badr[31]_INST_0_i_184_n_0 ;
  wire \badr[31]_INST_0_i_185_n_0 ;
  wire \badr[31]_INST_0_i_186_n_0 ;
  wire \badr[31]_INST_0_i_187_n_0 ;
  wire \badr[31]_INST_0_i_188_n_0 ;
  wire \badr[31]_INST_0_i_189_n_0 ;
  wire \badr[31]_INST_0_i_18_n_0 ;
  wire \badr[31]_INST_0_i_190_n_0 ;
  wire \badr[31]_INST_0_i_191_n_0 ;
  wire \badr[31]_INST_0_i_192_n_0 ;
  wire \badr[31]_INST_0_i_193_n_0 ;
  wire \badr[31]_INST_0_i_194_n_0 ;
  wire \badr[31]_INST_0_i_195_n_0 ;
  wire \badr[31]_INST_0_i_196_n_0 ;
  wire \badr[31]_INST_0_i_197_n_0 ;
  wire \badr[31]_INST_0_i_198_n_0 ;
  wire \badr[31]_INST_0_i_199_n_0 ;
  wire \badr[31]_INST_0_i_19_n_0 ;
  wire \badr[31]_INST_0_i_1_n_0 ;
  wire \badr[31]_INST_0_i_200_n_0 ;
  wire \badr[31]_INST_0_i_201_n_0 ;
  wire \badr[31]_INST_0_i_202_n_0 ;
  wire \badr[31]_INST_0_i_203_n_0 ;
  wire \badr[31]_INST_0_i_204_n_0 ;
  wire \badr[31]_INST_0_i_205_n_0 ;
  wire \badr[31]_INST_0_i_206_n_0 ;
  wire \badr[31]_INST_0_i_207_n_0 ;
  wire \badr[31]_INST_0_i_208_n_0 ;
  wire \badr[31]_INST_0_i_209_n_0 ;
  wire \badr[31]_INST_0_i_20_n_0 ;
  wire \badr[31]_INST_0_i_210_n_0 ;
  wire \badr[31]_INST_0_i_211_n_0 ;
  wire \badr[31]_INST_0_i_212_n_0 ;
  wire \badr[31]_INST_0_i_213_n_0 ;
  wire \badr[31]_INST_0_i_214_n_0 ;
  wire \badr[31]_INST_0_i_215_n_0 ;
  wire \badr[31]_INST_0_i_216_n_0 ;
  wire \badr[31]_INST_0_i_217_n_0 ;
  wire \badr[31]_INST_0_i_218_n_0 ;
  wire \badr[31]_INST_0_i_219_n_0 ;
  wire \badr[31]_INST_0_i_220_n_0 ;
  wire \badr[31]_INST_0_i_23_n_0 ;
  wire \badr[31]_INST_0_i_24_n_0 ;
  wire \badr[31]_INST_0_i_30_n_0 ;
  wire \badr[31]_INST_0_i_31_n_0 ;
  wire \badr[31]_INST_0_i_36_n_2 ;
  wire \badr[31]_INST_0_i_36_n_3 ;
  wire \badr[31]_INST_0_i_38_n_0 ;
  wire \badr[31]_INST_0_i_39_n_0 ;
  wire \badr[31]_INST_0_i_40_n_0 ;
  wire \badr[31]_INST_0_i_43_n_0 ;
  wire \badr[31]_INST_0_i_44_n_0 ;
  wire \badr[31]_INST_0_i_47_n_0 ;
  wire \badr[31]_INST_0_i_48_n_0 ;
  wire \badr[31]_INST_0_i_4_n_0 ;
  wire \badr[31]_INST_0_i_51_n_0 ;
  wire \badr[31]_INST_0_i_52_n_0 ;
  wire \badr[31]_INST_0_i_55_n_0 ;
  wire \badr[31]_INST_0_i_56_n_0 ;
  wire \badr[31]_INST_0_i_57_n_0 ;
  wire \badr[31]_INST_0_i_58_n_0 ;
  wire \badr[31]_INST_0_i_59_n_0 ;
  wire \badr[31]_INST_0_i_5_n_0 ;
  wire \badr[31]_INST_0_i_60_n_0 ;
  wire \badr[31]_INST_0_i_62_n_0 ;
  wire \badr[31]_INST_0_i_63_n_0 ;
  wire \badr[31]_INST_0_i_64_n_0 ;
  wire \badr[31]_INST_0_i_65_n_0 ;
  wire \badr[31]_INST_0_i_67_n_0 ;
  wire \badr[31]_INST_0_i_68_n_0 ;
  wire \badr[31]_INST_0_i_70_n_0 ;
  wire \badr[31]_INST_0_i_71_n_0 ;
  wire \badr[31]_INST_0_i_72_n_0 ;
  wire \badr[31]_INST_0_i_73_n_0 ;
  wire \badr[31]_INST_0_i_74_n_0 ;
  wire \badr[31]_INST_0_i_75_n_0 ;
  wire \badr[31]_INST_0_i_77_n_0 ;
  wire \badr[31]_INST_0_i_78_n_0 ;
  wire \badr[31]_INST_0_i_79_n_0 ;
  wire \badr[31]_INST_0_i_80_n_0 ;
  wire \badr[31]_INST_0_i_81_n_0 ;
  wire \badr[31]_INST_0_i_82_n_0 ;
  wire \badr[31]_INST_0_i_83_n_0 ;
  wire \badr[31]_INST_0_i_84_n_0 ;
  wire \badr[31]_INST_0_i_85_n_0 ;
  wire \badr[31]_INST_0_i_86_n_0 ;
  wire \badr[31]_INST_0_i_87_n_0 ;
  wire \badr[31]_INST_0_i_88_n_0 ;
  wire \badr[31]_INST_0_i_89_n_0 ;
  wire \badr[31]_INST_0_i_90_n_0 ;
  wire \badr[31]_INST_0_i_91_n_0 ;
  wire \badr[31]_INST_0_i_92_n_0 ;
  wire \badr[31]_INST_0_i_93_n_0 ;
  wire \badr[31]_INST_0_i_94_n_0 ;
  wire \badr[31]_INST_0_i_95_n_0 ;
  wire \badr[31]_INST_0_i_96_n_0 ;
  wire \badr[31]_INST_0_i_97_n_0 ;
  wire \badr[31]_INST_0_i_98_n_0 ;
  wire \badr[31]_INST_0_i_99_n_0 ;
  wire \badr[3]_INST_0_i_43_n_0 ;
  wire \badr[3]_INST_0_i_44_n_0 ;
  wire \badr[3]_INST_0_i_45_n_0 ;
  wire \badr[3]_INST_0_i_46_n_0 ;
  wire \badr[3]_INST_0_i_7_n_0 ;
  wire \badr[4]_INST_0_i_25_n_0 ;
  wire \badr[4]_INST_0_i_25_n_1 ;
  wire \badr[4]_INST_0_i_25_n_2 ;
  wire \badr[4]_INST_0_i_25_n_3 ;
  wire \badr[4]_INST_0_i_44_n_0 ;
  wire \badr[4]_INST_0_i_45_n_0 ;
  wire \badr[4]_INST_0_i_46_n_0 ;
  wire \badr[4]_INST_0_i_47_n_0 ;
  wire \badr[4]_INST_0_i_48_n_0 ;
  wire \badr[4]_INST_0_i_49_n_0 ;
  wire \badr[4]_INST_0_i_50_n_0 ;
  wire \badr[4]_INST_0_i_51_n_0 ;
  wire \badr[4]_INST_0_i_52_n_0 ;
  wire \badr[4]_INST_0_i_53_n_0 ;
  wire \badr[4]_INST_0_i_56_n_0 ;
  wire \badr[4]_INST_0_i_57_n_0 ;
  wire \badr[4]_INST_0_i_58_n_0 ;
  wire \badr[4]_INST_0_i_59_n_0 ;
  wire \badr[4]_INST_0_i_60_n_0 ;
  wire \badr[4]_INST_0_i_61_n_0 ;
  wire \badr[4]_INST_0_i_62_n_0 ;
  wire \badr[4]_INST_0_i_63_n_0 ;
  wire \badr[4]_INST_0_i_64_n_0 ;
  wire \badr[4]_INST_0_i_65_n_0 ;
  wire \badr[4]_INST_0_i_7_n_0 ;
  wire \badr[5]_INST_0_i_17_n_0 ;
  wire \badr[5]_INST_0_i_21_n_0 ;
  wire \badr[5]_INST_0_i_3_n_0 ;
  wire \badr[5]_INST_0_i_45_n_0 ;
  wire \badr[5]_INST_0_i_46_n_0 ;
  wire \badr[5]_INST_0_i_47_n_0 ;
  wire \badr[5]_INST_0_i_48_n_0 ;
  wire \badr[5]_INST_0_i_9_n_0 ;
  wire \badr[6]_INST_0_i_17_n_0 ;
  wire \badr[6]_INST_0_i_21_n_0 ;
  wire \badr[6]_INST_0_i_3_n_0 ;
  wire \badr[6]_INST_0_i_45_n_0 ;
  wire \badr[6]_INST_0_i_46_n_0 ;
  wire \badr[6]_INST_0_i_47_n_0 ;
  wire \badr[6]_INST_0_i_48_n_0 ;
  wire \badr[6]_INST_0_i_9_n_0 ;
  wire \badr[7]_INST_0_i_17_n_0 ;
  wire \badr[7]_INST_0_i_21_n_0 ;
  wire \badr[7]_INST_0_i_3_n_0 ;
  wire \badr[7]_INST_0_i_45_n_0 ;
  wire \badr[7]_INST_0_i_46_n_0 ;
  wire \badr[7]_INST_0_i_47_n_0 ;
  wire \badr[7]_INST_0_i_48_n_0 ;
  wire \badr[7]_INST_0_i_9_n_0 ;
  wire \badr[8]_INST_0_i_17_n_0 ;
  wire \badr[8]_INST_0_i_21_n_0 ;
  wire \badr[8]_INST_0_i_29_n_0 ;
  wire \badr[8]_INST_0_i_29_n_1 ;
  wire \badr[8]_INST_0_i_29_n_2 ;
  wire \badr[8]_INST_0_i_29_n_3 ;
  wire \badr[8]_INST_0_i_3_n_0 ;
  wire \badr[8]_INST_0_i_46_n_0 ;
  wire \badr[8]_INST_0_i_47_n_0 ;
  wire \badr[8]_INST_0_i_48_n_0 ;
  wire \badr[8]_INST_0_i_49_n_0 ;
  wire \badr[8]_INST_0_i_50_n_0 ;
  wire \badr[8]_INST_0_i_51_n_0 ;
  wire \badr[8]_INST_0_i_52_n_0 ;
  wire \badr[8]_INST_0_i_53_n_0 ;
  wire \badr[8]_INST_0_i_9_n_0 ;
  wire \badr[9]_INST_0_i_17_n_0 ;
  wire \badr[9]_INST_0_i_21_n_0 ;
  wire \badr[9]_INST_0_i_3_n_0 ;
  wire \badr[9]_INST_0_i_45_n_0 ;
  wire \badr[9]_INST_0_i_46_n_0 ;
  wire \badr[9]_INST_0_i_47_n_0 ;
  wire \badr[9]_INST_0_i_48_n_0 ;
  wire \badr[9]_INST_0_i_9_n_0 ;
  wire \bank02/a0buso/gr0_bus1 ;
  wire \bank02/a0buso/gr1_bus1 ;
  wire \bank02/a0buso/gr2_bus1 ;
  wire \bank02/a0buso/gr3_bus1 ;
  wire \bank02/a0buso/gr4_bus1 ;
  wire \bank02/a0buso/gr5_bus1 ;
  wire \bank02/a0buso/gr6_bus1 ;
  wire \bank02/a0buso/gr7_bus1 ;
  wire \bank02/a0buso2h/gr0_bus1 ;
  wire \bank02/a0buso2h/gr3_bus1 ;
  wire \bank02/a0buso2h/gr4_bus1 ;
  wire \bank02/a0buso2h/gr7_bus1 ;
  wire \bank02/a0buso2l/gr0_bus1 ;
  wire \bank02/a0buso2l/gr1_bus1 ;
  wire \bank02/a0buso2l/gr2_bus1 ;
  wire \bank02/a0buso2l/gr3_bus1 ;
  wire \bank02/a0buso2l/gr4_bus1 ;
  wire \bank02/a0buso2l/gr5_bus1 ;
  wire \bank02/a0buso2l/gr6_bus1 ;
  wire \bank02/a0buso2l/gr7_bus1 ;
  wire \bank02/a1buso/gr0_bus1 ;
  wire \bank02/a1buso/gr2_bus1 ;
  wire \bank02/a1buso/gr3_bus1 ;
  wire \bank02/a1buso/gr4_bus1 ;
  wire \bank02/a1buso/gr5_bus1 ;
  wire \bank02/a1buso/gr6_bus1 ;
  wire \bank02/a1buso/gr7_bus1 ;
  wire \bank02/a1buso2h/gr0_bus1 ;
  wire \bank02/a1buso2h/gr3_bus1 ;
  wire \bank02/a1buso2h/gr4_bus1 ;
  wire \bank02/a1buso2h/gr7_bus1 ;
  wire \bank02/a1buso2l/gr0_bus1 ;
  wire \bank02/a1buso2l/gr2_bus1 ;
  wire \bank02/a1buso2l/gr3_bus1 ;
  wire \bank02/a1buso2l/gr4_bus1 ;
  wire \bank02/a1buso2l/gr5_bus1 ;
  wire \bank02/a1buso2l/gr6_bus1 ;
  wire \bank02/a1buso2l/gr7_bus1 ;
  wire \bank02/b0buso/gr0_bus1 ;
  wire \bank02/b0buso/gr1_bus1 ;
  wire \bank02/b0buso/gr2_bus1 ;
  wire \bank02/b0buso/gr3_bus1 ;
  wire \bank02/b0buso/gr4_bus1 ;
  wire \bank02/b0buso/gr5_bus1 ;
  wire \bank02/b0buso/gr6_bus1 ;
  wire \bank02/b0buso/gr7_bus1 ;
  wire \bank02/b0buso2l/gr0_bus1 ;
  wire \bank02/b0buso2l/gr1_bus1 ;
  wire \bank02/b0buso2l/gr2_bus1 ;
  wire \bank02/b0buso2l/gr3_bus1 ;
  wire \bank02/b0buso2l/gr4_bus1 ;
  wire \bank02/b0buso2l/gr5_bus1 ;
  wire \bank02/b0buso2l/gr6_bus1 ;
  wire \bank02/b0buso2l/gr7_bus1 ;
  wire \bank02/b1buso/gr0_bus1 ;
  wire \bank02/b1buso/gr1_bus1 ;
  wire \bank02/b1buso/gr2_bus1 ;
  wire \bank02/b1buso/gr3_bus1 ;
  wire \bank02/b1buso/gr4_bus1 ;
  wire \bank02/b1buso/gr5_bus1 ;
  wire \bank02/b1buso/gr6_bus1 ;
  wire \bank02/b1buso/gr7_bus1 ;
  wire \bank02/b1buso2l/gr0_bus1 ;
  wire \bank02/b1buso2l/gr2_bus1 ;
  wire \bank02/b1buso2l/gr3_bus1 ;
  wire \bank02/b1buso2l/gr4_bus1 ;
  wire \bank02/b1buso2l/gr5_bus1 ;
  wire \bank02/b1buso2l/gr6_bus1 ;
  wire \bank02/b1buso2l/gr7_bus1 ;
  wire \bank13/a0buso/gr0_bus1 ;
  wire \bank13/a0buso/gr3_bus1 ;
  wire \bank13/a0buso/gr4_bus1 ;
  wire \bank13/a0buso/gr7_bus1 ;
  wire \bank13/a0buso2h/gr0_bus1 ;
  wire \bank13/a0buso2h/gr3_bus1 ;
  wire \bank13/a0buso2h/gr4_bus1 ;
  wire \bank13/a0buso2h/gr7_bus1 ;
  wire \bank13/a0buso2l/gr0_bus1 ;
  wire \bank13/a0buso2l/gr1_bus1 ;
  wire \bank13/a0buso2l/gr2_bus1 ;
  wire \bank13/a0buso2l/gr3_bus1 ;
  wire \bank13/a0buso2l/gr4_bus1 ;
  wire \bank13/a0buso2l/gr5_bus1 ;
  wire \bank13/a0buso2l/gr6_bus1 ;
  wire \bank13/a0buso2l/gr7_bus1 ;
  wire \bank13/a1buso/gr0_bus1 ;
  wire \bank13/a1buso/gr3_bus1 ;
  wire \bank13/a1buso/gr4_bus1 ;
  wire \bank13/a1buso/gr5_bus1 ;
  wire \bank13/a1buso/gr6_bus1 ;
  wire \bank13/a1buso/gr7_bus1 ;
  wire \bank13/a1buso2h/gr0_bus1 ;
  wire \bank13/a1buso2h/gr3_bus1 ;
  wire \bank13/a1buso2h/gr4_bus1 ;
  wire \bank13/a1buso2h/gr7_bus1 ;
  wire \bank13/a1buso2l/gr0_bus1 ;
  wire \bank13/a1buso2l/gr3_bus1 ;
  wire \bank13/a1buso2l/gr4_bus1 ;
  wire \bank13/a1buso2l/gr5_bus1 ;
  wire \bank13/a1buso2l/gr6_bus1 ;
  wire \bank13/a1buso2l/gr7_bus1 ;
  wire \bank13/b0buso/gr0_bus1 ;
  wire \bank13/b0buso/gr1_bus1 ;
  wire \bank13/b0buso/gr2_bus1 ;
  wire \bank13/b0buso/gr3_bus1 ;
  wire \bank13/b0buso/gr4_bus1 ;
  wire \bank13/b0buso/gr5_bus1 ;
  wire \bank13/b0buso/gr6_bus1 ;
  wire \bank13/b0buso/gr7_bus1 ;
  wire \bank13/b0buso2h/gr0_bus1 ;
  wire \bank13/b0buso2h/gr3_bus1 ;
  wire \bank13/b0buso2h/gr4_bus1 ;
  wire \bank13/b0buso2h/gr7_bus1 ;
  wire \bank13/b0buso2l/gr0_bus1 ;
  wire \bank13/b0buso2l/gr1_bus1 ;
  wire \bank13/b0buso2l/gr2_bus1 ;
  wire \bank13/b0buso2l/gr3_bus1 ;
  wire \bank13/b0buso2l/gr4_bus1 ;
  wire \bank13/b0buso2l/gr5_bus1 ;
  wire \bank13/b0buso2l/gr6_bus1 ;
  wire \bank13/b0buso2l/gr7_bus1 ;
  wire \bank13/b1buso/gr0_bus1 ;
  wire \bank13/b1buso/gr2_bus1 ;
  wire \bank13/b1buso/gr3_bus1 ;
  wire \bank13/b1buso/gr4_bus1 ;
  wire \bank13/b1buso/gr5_bus1 ;
  wire \bank13/b1buso/gr6_bus1 ;
  wire \bank13/b1buso/gr7_bus1 ;
  wire \bank13/b1buso2h/gr0_bus1 ;
  wire \bank13/b1buso2h/gr3_bus1 ;
  wire \bank13/b1buso2h/gr4_bus1 ;
  wire \bank13/b1buso2h/gr7_bus1 ;
  wire \bank13/b1buso2l/gr0_bus1 ;
  wire \bank13/b1buso2l/gr2_bus1 ;
  wire \bank13/b1buso2l/gr3_bus1 ;
  wire \bank13/b1buso2l/gr4_bus1 ;
  wire \bank13/b1buso2l/gr5_bus1 ;
  wire \bank13/b1buso2l/gr6_bus1 ;
  wire \bank13/b1buso2l/gr7_bus1 ;
  wire [31:0]bbus_o;
  wire \bbus_o[0]_INST_0_i_1_n_0 ;
  wire \bbus_o[0]_INST_0_i_2_n_0 ;
  wire \bbus_o[0]_INST_0_i_8_n_0 ;
  wire \bbus_o[1]_INST_0_i_1_n_0 ;
  wire \bbus_o[1]_INST_0_i_2_n_0 ;
  wire \bbus_o[2]_INST_0_i_1_n_0 ;
  wire \bbus_o[2]_INST_0_i_2_n_0 ;
  wire \bbus_o[3]_INST_0_i_1_n_0 ;
  wire \bbus_o[3]_INST_0_i_2_n_0 ;
  wire \bbus_o[3]_INST_0_i_7_n_0 ;
  wire \bbus_o[4]_INST_0_i_1_n_0 ;
  wire \bbus_o[4]_INST_0_i_2_n_0 ;
  wire \bbus_o[5]_INST_0_i_10_n_0 ;
  wire \bbus_o[5]_INST_0_i_11_n_0 ;
  wire \bbus_o[5]_INST_0_i_12_n_0 ;
  wire \bbus_o[5]_INST_0_i_13_n_0 ;
  wire \bbus_o[5]_INST_0_i_1_n_0 ;
  wire \bbus_o[5]_INST_0_i_24_n_0 ;
  wire \bbus_o[5]_INST_0_i_25_n_0 ;
  wire \bbus_o[5]_INST_0_i_26_n_0 ;
  wire \bbus_o[5]_INST_0_i_2_n_0 ;
  wire \bbus_o[5]_INST_0_i_3_n_0 ;
  wire \bbus_o[5]_INST_0_i_8_n_0 ;
  wire \bbus_o[5]_INST_0_i_9_n_0 ;
  wire \bbus_o[6]_INST_0_i_1_n_0 ;
  wire \bbus_o[6]_INST_0_i_2_n_0 ;
  wire \bbus_o[6]_INST_0_i_5_n_0 ;
  wire \bbus_o[7]_INST_0_i_2_n_0 ;
  wire \bbus_o[7]_INST_0_i_5_n_0 ;
  wire [3:0]bcmd;
  wire \bcmd[0]_INST_0_i_10_n_0 ;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_13_n_0 ;
  wire \bcmd[0]_INST_0_i_14_n_0 ;
  wire \bcmd[0]_INST_0_i_15_n_0 ;
  wire \bcmd[0]_INST_0_i_16_n_0 ;
  wire \bcmd[0]_INST_0_i_17_n_0 ;
  wire \bcmd[0]_INST_0_i_18_n_0 ;
  wire \bcmd[0]_INST_0_i_19_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_20_n_0 ;
  wire \bcmd[0]_INST_0_i_21_n_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_3_n_0 ;
  wire \bcmd[0]_INST_0_i_4_n_0 ;
  wire \bcmd[0]_INST_0_i_5_n_0 ;
  wire \bcmd[0]_INST_0_i_6_n_0 ;
  wire \bcmd[0]_INST_0_i_7_n_0 ;
  wire \bcmd[0]_INST_0_i_8_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_11_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_14_n_0 ;
  wire \bcmd[1]_INST_0_i_15_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_17_n_0 ;
  wire \bcmd[1]_INST_0_i_18_n_0 ;
  wire \bcmd[1]_INST_0_i_19_n_0 ;
  wire \bcmd[1]_INST_0_i_1_n_0 ;
  wire \bcmd[1]_INST_0_i_20_n_0 ;
  wire \bcmd[1]_INST_0_i_21_n_0 ;
  wire \bcmd[1]_INST_0_i_22_n_0 ;
  wire \bcmd[1]_INST_0_i_23_n_0 ;
  wire \bcmd[1]_INST_0_i_24_n_0 ;
  wire \bcmd[1]_INST_0_i_25_n_0 ;
  wire \bcmd[1]_INST_0_i_26_n_0 ;
  wire \bcmd[1]_INST_0_i_27_n_0 ;
  wire \bcmd[1]_INST_0_i_28_n_0 ;
  wire \bcmd[1]_INST_0_i_29_n_0 ;
  wire \bcmd[1]_INST_0_i_2_n_0 ;
  wire \bcmd[1]_INST_0_i_3_n_0 ;
  wire \bcmd[1]_INST_0_i_4_n_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_6_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_8_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2]_INST_0_i_1_n_0 ;
  wire \bcmd[2]_INST_0_i_2_n_0 ;
  wire \bcmd[2]_INST_0_i_3_n_0 ;
  wire \bcmd[2]_INST_0_i_4_n_0 ;
  wire \bcmd[2]_INST_0_i_5_n_0 ;
  wire \bcmd[2]_INST_0_i_6_n_0 ;
  wire \bcmd[2]_INST_0_i_7_n_0 ;
  wire \bcmd[2]_INST_0_i_8_n_0 ;
  wire \bcmd[3]_INST_0_i_10_n_0 ;
  wire \bcmd[3]_INST_0_i_11_n_0 ;
  wire \bcmd[3]_INST_0_i_12_n_0 ;
  wire \bcmd[3]_INST_0_i_13_n_0 ;
  wire \bcmd[3]_INST_0_i_14_n_0 ;
  wire \bcmd[3]_INST_0_i_15_n_0 ;
  wire \bcmd[3]_INST_0_i_16_n_0 ;
  wire \bcmd[3]_INST_0_i_17_n_0 ;
  wire \bcmd[3]_INST_0_i_18_n_0 ;
  wire \bcmd[3]_INST_0_i_19_n_0 ;
  wire \bcmd[3]_INST_0_i_1_n_0 ;
  wire \bcmd[3]_INST_0_i_20_n_0 ;
  wire \bcmd[3]_INST_0_i_21_n_0 ;
  wire \bcmd[3]_INST_0_i_22_n_0 ;
  wire \bcmd[3]_INST_0_i_23_n_0 ;
  wire \bcmd[3]_INST_0_i_24_n_0 ;
  wire \bcmd[3]_INST_0_i_2_n_0 ;
  wire \bcmd[3]_INST_0_i_3_n_0 ;
  wire \bcmd[3]_INST_0_i_4_n_0 ;
  wire \bcmd[3]_INST_0_i_5_n_0 ;
  wire \bcmd[3]_INST_0_i_6_n_0 ;
  wire \bcmd[3]_INST_0_i_7_n_0 ;
  wire \bcmd[3]_INST_0_i_8_n_0 ;
  wire \bcmd[3]_INST_0_i_9_n_0 ;
  wire [31:0]bdatr;
  wire [31:0]bdatw;
  wire \bdatw[10]_INST_0_i_12_n_0 ;
  wire \bdatw[10]_INST_0_i_13_n_0 ;
  wire \bdatw[10]_INST_0_i_19_n_0 ;
  wire \bdatw[10]_INST_0_i_3_n_0 ;
  wire \bdatw[10]_INST_0_i_4_n_0 ;
  wire \bdatw[10]_INST_0_i_5_n_0 ;
  wire \bdatw[10]_INST_0_i_9_n_0 ;
  wire \bdatw[11]_INST_0_i_12_n_0 ;
  wire \bdatw[11]_INST_0_i_18_n_0 ;
  wire \bdatw[11]_INST_0_i_19_n_0 ;
  wire \bdatw[11]_INST_0_i_3_n_0 ;
  wire \bdatw[11]_INST_0_i_4_n_0 ;
  wire \bdatw[11]_INST_0_i_5_n_0 ;
  wire \bdatw[11]_INST_0_i_9_n_0 ;
  wire \bdatw[12]_INST_0_i_11_n_0 ;
  wire \bdatw[12]_INST_0_i_1_n_0 ;
  wire \bdatw[12]_INST_0_i_22_n_0 ;
  wire \bdatw[12]_INST_0_i_23_n_0 ;
  wire \bdatw[12]_INST_0_i_29_n_0 ;
  wire \bdatw[12]_INST_0_i_33_n_0 ;
  wire \bdatw[12]_INST_0_i_34_n_0 ;
  wire \bdatw[12]_INST_0_i_4_n_0 ;
  wire \bdatw[12]_INST_0_i_5_n_0 ;
  wire \bdatw[12]_INST_0_i_60_n_0 ;
  wire \bdatw[12]_INST_0_i_61_n_0 ;
  wire \bdatw[12]_INST_0_i_62_n_0 ;
  wire \bdatw[12]_INST_0_i_63_n_0 ;
  wire \bdatw[12]_INST_0_i_64_n_0 ;
  wire \bdatw[12]_INST_0_i_65_n_0 ;
  wire \bdatw[12]_INST_0_i_66_n_0 ;
  wire \bdatw[12]_INST_0_i_67_n_0 ;
  wire \bdatw[12]_INST_0_i_8_n_0 ;
  wire \bdatw[13]_INST_0_i_1_n_0 ;
  wire \bdatw[13]_INST_0_i_4_n_0 ;
  wire \bdatw[13]_INST_0_i_7_n_0 ;
  wire \bdatw[14]_INST_0_i_3_n_0 ;
  wire \bdatw[14]_INST_0_i_4_n_0 ;
  wire \bdatw[14]_INST_0_i_8_n_0 ;
  wire \bdatw[15]_INST_0_i_11_n_0 ;
  wire \bdatw[15]_INST_0_i_14_n_0 ;
  wire \bdatw[15]_INST_0_i_1_n_0 ;
  wire \bdatw[15]_INST_0_i_22_n_0 ;
  wire \bdatw[15]_INST_0_i_4_n_0 ;
  wire \bdatw[15]_INST_0_i_5_n_0 ;
  wire \bdatw[15]_INST_0_i_63_n_0 ;
  wire \bdatw[15]_INST_0_i_64_n_0 ;
  wire \bdatw[15]_INST_0_i_6_n_0 ;
  wire \bdatw[15]_INST_0_i_7_n_0 ;
  wire \bdatw[15]_INST_0_i_90_n_0 ;
  wire \bdatw[15]_INST_0_i_91_n_0 ;
  wire \bdatw[15]_INST_0_i_92_n_0 ;
  wire \bdatw[15]_INST_0_i_93_n_0 ;
  wire \bdatw[15]_INST_0_i_94_n_0 ;
  wire \bdatw[15]_INST_0_i_95_n_0 ;
  wire \bdatw[15]_INST_0_i_96_n_0 ;
  wire \bdatw[16]_INST_0_i_10_n_0 ;
  wire \bdatw[16]_INST_0_i_13_n_0 ;
  wire \bdatw[16]_INST_0_i_14_n_0 ;
  wire \bdatw[16]_INST_0_i_15_n_0 ;
  wire \bdatw[16]_INST_0_i_16_n_0 ;
  wire \bdatw[16]_INST_0_i_19_n_0 ;
  wire \bdatw[16]_INST_0_i_20_n_0 ;
  wire \bdatw[16]_INST_0_i_21_n_0 ;
  wire \bdatw[16]_INST_0_i_22_n_0 ;
  wire \bdatw[16]_INST_0_i_7_n_0 ;
  wire \bdatw[16]_INST_0_i_8_n_0 ;
  wire \bdatw[16]_INST_0_i_9_n_0 ;
  wire \bdatw[17]_INST_0_i_10_n_0 ;
  wire \bdatw[17]_INST_0_i_13_n_0 ;
  wire \bdatw[17]_INST_0_i_14_n_0 ;
  wire \bdatw[17]_INST_0_i_15_n_0 ;
  wire \bdatw[17]_INST_0_i_16_n_0 ;
  wire \bdatw[17]_INST_0_i_19_n_0 ;
  wire \bdatw[17]_INST_0_i_20_n_0 ;
  wire \bdatw[17]_INST_0_i_21_n_0 ;
  wire \bdatw[17]_INST_0_i_22_n_0 ;
  wire \bdatw[17]_INST_0_i_7_n_0 ;
  wire \bdatw[17]_INST_0_i_8_n_0 ;
  wire \bdatw[17]_INST_0_i_9_n_0 ;
  wire \bdatw[18]_INST_0_i_10_n_0 ;
  wire \bdatw[18]_INST_0_i_13_n_0 ;
  wire \bdatw[18]_INST_0_i_14_n_0 ;
  wire \bdatw[18]_INST_0_i_15_n_0 ;
  wire \bdatw[18]_INST_0_i_16_n_0 ;
  wire \bdatw[18]_INST_0_i_19_n_0 ;
  wire \bdatw[18]_INST_0_i_20_n_0 ;
  wire \bdatw[18]_INST_0_i_21_n_0 ;
  wire \bdatw[18]_INST_0_i_22_n_0 ;
  wire \bdatw[18]_INST_0_i_7_n_0 ;
  wire \bdatw[18]_INST_0_i_8_n_0 ;
  wire \bdatw[18]_INST_0_i_9_n_0 ;
  wire \bdatw[19]_INST_0_i_10_n_0 ;
  wire \bdatw[19]_INST_0_i_13_n_0 ;
  wire \bdatw[19]_INST_0_i_14_n_0 ;
  wire \bdatw[19]_INST_0_i_15_n_0 ;
  wire \bdatw[19]_INST_0_i_16_n_0 ;
  wire \bdatw[19]_INST_0_i_19_n_0 ;
  wire \bdatw[19]_INST_0_i_20_n_0 ;
  wire \bdatw[19]_INST_0_i_21_n_0 ;
  wire \bdatw[19]_INST_0_i_22_n_0 ;
  wire \bdatw[19]_INST_0_i_7_n_0 ;
  wire \bdatw[19]_INST_0_i_8_n_0 ;
  wire \bdatw[19]_INST_0_i_9_n_0 ;
  wire \bdatw[20]_INST_0_i_10_n_0 ;
  wire \bdatw[20]_INST_0_i_13_n_0 ;
  wire \bdatw[20]_INST_0_i_14_n_0 ;
  wire \bdatw[20]_INST_0_i_15_n_0 ;
  wire \bdatw[20]_INST_0_i_16_n_0 ;
  wire \bdatw[20]_INST_0_i_19_n_0 ;
  wire \bdatw[20]_INST_0_i_20_n_0 ;
  wire \bdatw[20]_INST_0_i_21_n_0 ;
  wire \bdatw[20]_INST_0_i_22_n_0 ;
  wire \bdatw[20]_INST_0_i_7_n_0 ;
  wire \bdatw[20]_INST_0_i_8_n_0 ;
  wire \bdatw[20]_INST_0_i_9_n_0 ;
  wire \bdatw[21]_INST_0_i_10_n_0 ;
  wire \bdatw[21]_INST_0_i_13_n_0 ;
  wire \bdatw[21]_INST_0_i_14_n_0 ;
  wire \bdatw[21]_INST_0_i_15_n_0 ;
  wire \bdatw[21]_INST_0_i_16_n_0 ;
  wire \bdatw[21]_INST_0_i_19_n_0 ;
  wire \bdatw[21]_INST_0_i_20_n_0 ;
  wire \bdatw[21]_INST_0_i_21_n_0 ;
  wire \bdatw[21]_INST_0_i_22_n_0 ;
  wire \bdatw[21]_INST_0_i_7_n_0 ;
  wire \bdatw[21]_INST_0_i_8_n_0 ;
  wire \bdatw[21]_INST_0_i_9_n_0 ;
  wire \bdatw[22]_INST_0_i_10_n_0 ;
  wire \bdatw[22]_INST_0_i_13_n_0 ;
  wire \bdatw[22]_INST_0_i_14_n_0 ;
  wire \bdatw[22]_INST_0_i_15_n_0 ;
  wire \bdatw[22]_INST_0_i_16_n_0 ;
  wire \bdatw[22]_INST_0_i_19_n_0 ;
  wire \bdatw[22]_INST_0_i_20_n_0 ;
  wire \bdatw[22]_INST_0_i_21_n_0 ;
  wire \bdatw[22]_INST_0_i_22_n_0 ;
  wire \bdatw[22]_INST_0_i_7_n_0 ;
  wire \bdatw[22]_INST_0_i_8_n_0 ;
  wire \bdatw[22]_INST_0_i_9_n_0 ;
  wire \bdatw[23]_INST_0_i_10_n_0 ;
  wire \bdatw[23]_INST_0_i_13_n_0 ;
  wire \bdatw[23]_INST_0_i_14_n_0 ;
  wire \bdatw[23]_INST_0_i_15_n_0 ;
  wire \bdatw[23]_INST_0_i_16_n_0 ;
  wire \bdatw[23]_INST_0_i_19_n_0 ;
  wire \bdatw[23]_INST_0_i_20_n_0 ;
  wire \bdatw[23]_INST_0_i_21_n_0 ;
  wire \bdatw[23]_INST_0_i_22_n_0 ;
  wire \bdatw[23]_INST_0_i_7_n_0 ;
  wire \bdatw[23]_INST_0_i_8_n_0 ;
  wire \bdatw[23]_INST_0_i_9_n_0 ;
  wire \bdatw[24]_INST_0_i_10_n_0 ;
  wire \bdatw[24]_INST_0_i_13_n_0 ;
  wire \bdatw[24]_INST_0_i_14_n_0 ;
  wire \bdatw[24]_INST_0_i_15_n_0 ;
  wire \bdatw[24]_INST_0_i_16_n_0 ;
  wire \bdatw[24]_INST_0_i_19_n_0 ;
  wire \bdatw[24]_INST_0_i_20_n_0 ;
  wire \bdatw[24]_INST_0_i_21_n_0 ;
  wire \bdatw[24]_INST_0_i_22_n_0 ;
  wire \bdatw[24]_INST_0_i_7_n_0 ;
  wire \bdatw[24]_INST_0_i_8_n_0 ;
  wire \bdatw[24]_INST_0_i_9_n_0 ;
  wire \bdatw[25]_INST_0_i_10_n_0 ;
  wire \bdatw[25]_INST_0_i_13_n_0 ;
  wire \bdatw[25]_INST_0_i_14_n_0 ;
  wire \bdatw[25]_INST_0_i_15_n_0 ;
  wire \bdatw[25]_INST_0_i_16_n_0 ;
  wire \bdatw[25]_INST_0_i_19_n_0 ;
  wire \bdatw[25]_INST_0_i_20_n_0 ;
  wire \bdatw[25]_INST_0_i_21_n_0 ;
  wire \bdatw[25]_INST_0_i_22_n_0 ;
  wire \bdatw[25]_INST_0_i_7_n_0 ;
  wire \bdatw[25]_INST_0_i_8_n_0 ;
  wire \bdatw[25]_INST_0_i_9_n_0 ;
  wire \bdatw[26]_INST_0_i_10_n_0 ;
  wire \bdatw[26]_INST_0_i_13_n_0 ;
  wire \bdatw[26]_INST_0_i_14_n_0 ;
  wire \bdatw[26]_INST_0_i_15_n_0 ;
  wire \bdatw[26]_INST_0_i_16_n_0 ;
  wire \bdatw[26]_INST_0_i_19_n_0 ;
  wire \bdatw[26]_INST_0_i_20_n_0 ;
  wire \bdatw[26]_INST_0_i_21_n_0 ;
  wire \bdatw[26]_INST_0_i_22_n_0 ;
  wire \bdatw[26]_INST_0_i_7_n_0 ;
  wire \bdatw[26]_INST_0_i_8_n_0 ;
  wire \bdatw[26]_INST_0_i_9_n_0 ;
  wire \bdatw[27]_INST_0_i_10_n_0 ;
  wire \bdatw[27]_INST_0_i_13_n_0 ;
  wire \bdatw[27]_INST_0_i_14_n_0 ;
  wire \bdatw[27]_INST_0_i_15_n_0 ;
  wire \bdatw[27]_INST_0_i_16_n_0 ;
  wire \bdatw[27]_INST_0_i_19_n_0 ;
  wire \bdatw[27]_INST_0_i_20_n_0 ;
  wire \bdatw[27]_INST_0_i_21_n_0 ;
  wire \bdatw[27]_INST_0_i_22_n_0 ;
  wire \bdatw[27]_INST_0_i_7_n_0 ;
  wire \bdatw[27]_INST_0_i_8_n_0 ;
  wire \bdatw[27]_INST_0_i_9_n_0 ;
  wire \bdatw[28]_INST_0_i_10_n_0 ;
  wire \bdatw[28]_INST_0_i_13_n_0 ;
  wire \bdatw[28]_INST_0_i_14_n_0 ;
  wire \bdatw[28]_INST_0_i_15_n_0 ;
  wire \bdatw[28]_INST_0_i_16_n_0 ;
  wire \bdatw[28]_INST_0_i_19_n_0 ;
  wire \bdatw[28]_INST_0_i_20_n_0 ;
  wire \bdatw[28]_INST_0_i_21_n_0 ;
  wire \bdatw[28]_INST_0_i_22_n_0 ;
  wire \bdatw[28]_INST_0_i_7_n_0 ;
  wire \bdatw[28]_INST_0_i_8_n_0 ;
  wire \bdatw[28]_INST_0_i_9_n_0 ;
  wire \bdatw[29]_INST_0_i_10_n_0 ;
  wire \bdatw[29]_INST_0_i_13_n_0 ;
  wire \bdatw[29]_INST_0_i_14_n_0 ;
  wire \bdatw[29]_INST_0_i_15_n_0 ;
  wire \bdatw[29]_INST_0_i_16_n_0 ;
  wire \bdatw[29]_INST_0_i_19_n_0 ;
  wire \bdatw[29]_INST_0_i_20_n_0 ;
  wire \bdatw[29]_INST_0_i_21_n_0 ;
  wire \bdatw[29]_INST_0_i_22_n_0 ;
  wire \bdatw[29]_INST_0_i_7_n_0 ;
  wire \bdatw[29]_INST_0_i_8_n_0 ;
  wire \bdatw[29]_INST_0_i_9_n_0 ;
  wire \bdatw[30]_INST_0_i_10_n_0 ;
  wire \bdatw[30]_INST_0_i_13_n_0 ;
  wire \bdatw[30]_INST_0_i_14_n_0 ;
  wire \bdatw[30]_INST_0_i_15_n_0 ;
  wire \bdatw[30]_INST_0_i_16_n_0 ;
  wire \bdatw[30]_INST_0_i_19_n_0 ;
  wire \bdatw[30]_INST_0_i_20_n_0 ;
  wire \bdatw[30]_INST_0_i_21_n_0 ;
  wire \bdatw[30]_INST_0_i_22_n_0 ;
  wire \bdatw[30]_INST_0_i_7_n_0 ;
  wire \bdatw[30]_INST_0_i_8_n_0 ;
  wire \bdatw[30]_INST_0_i_9_n_0 ;
  wire \bdatw[31]_INST_0_i_100_n_0 ;
  wire \bdatw[31]_INST_0_i_101_n_0 ;
  wire \bdatw[31]_INST_0_i_102_n_0 ;
  wire \bdatw[31]_INST_0_i_103_n_0 ;
  wire \bdatw[31]_INST_0_i_104_n_0 ;
  wire \bdatw[31]_INST_0_i_105_n_0 ;
  wire \bdatw[31]_INST_0_i_106_n_0 ;
  wire \bdatw[31]_INST_0_i_107_n_0 ;
  wire \bdatw[31]_INST_0_i_108_n_0 ;
  wire \bdatw[31]_INST_0_i_109_n_0 ;
  wire \bdatw[31]_INST_0_i_110_n_0 ;
  wire \bdatw[31]_INST_0_i_111_n_0 ;
  wire \bdatw[31]_INST_0_i_112_n_0 ;
  wire \bdatw[31]_INST_0_i_113_n_0 ;
  wire \bdatw[31]_INST_0_i_114_n_0 ;
  wire \bdatw[31]_INST_0_i_115_n_0 ;
  wire \bdatw[31]_INST_0_i_116_n_0 ;
  wire \bdatw[31]_INST_0_i_117_n_0 ;
  wire \bdatw[31]_INST_0_i_118_n_0 ;
  wire \bdatw[31]_INST_0_i_119_n_0 ;
  wire \bdatw[31]_INST_0_i_11_n_0 ;
  wire \bdatw[31]_INST_0_i_120_n_0 ;
  wire \bdatw[31]_INST_0_i_121_n_0 ;
  wire \bdatw[31]_INST_0_i_122_n_0 ;
  wire \bdatw[31]_INST_0_i_123_n_0 ;
  wire \bdatw[31]_INST_0_i_124_n_0 ;
  wire \bdatw[31]_INST_0_i_125_n_0 ;
  wire \bdatw[31]_INST_0_i_126_n_0 ;
  wire \bdatw[31]_INST_0_i_127_n_0 ;
  wire \bdatw[31]_INST_0_i_128_n_0 ;
  wire \bdatw[31]_INST_0_i_129_n_0 ;
  wire \bdatw[31]_INST_0_i_12_n_0 ;
  wire \bdatw[31]_INST_0_i_130_n_0 ;
  wire \bdatw[31]_INST_0_i_131_n_0 ;
  wire \bdatw[31]_INST_0_i_132_n_0 ;
  wire \bdatw[31]_INST_0_i_133_n_0 ;
  wire \bdatw[31]_INST_0_i_134_n_0 ;
  wire \bdatw[31]_INST_0_i_135_n_0 ;
  wire \bdatw[31]_INST_0_i_136_n_0 ;
  wire \bdatw[31]_INST_0_i_137_n_0 ;
  wire \bdatw[31]_INST_0_i_138_n_0 ;
  wire \bdatw[31]_INST_0_i_139_n_0 ;
  wire \bdatw[31]_INST_0_i_13_n_0 ;
  wire \bdatw[31]_INST_0_i_140_n_0 ;
  wire \bdatw[31]_INST_0_i_141_n_0 ;
  wire \bdatw[31]_INST_0_i_142_n_0 ;
  wire \bdatw[31]_INST_0_i_143_n_0 ;
  wire \bdatw[31]_INST_0_i_144_n_0 ;
  wire \bdatw[31]_INST_0_i_145_n_0 ;
  wire \bdatw[31]_INST_0_i_146_n_0 ;
  wire \bdatw[31]_INST_0_i_147_n_0 ;
  wire \bdatw[31]_INST_0_i_148_n_0 ;
  wire \bdatw[31]_INST_0_i_149_n_0 ;
  wire \bdatw[31]_INST_0_i_14_n_0 ;
  wire \bdatw[31]_INST_0_i_150_n_0 ;
  wire \bdatw[31]_INST_0_i_151_n_0 ;
  wire \bdatw[31]_INST_0_i_152_n_0 ;
  wire \bdatw[31]_INST_0_i_153_n_0 ;
  wire \bdatw[31]_INST_0_i_154_n_0 ;
  wire \bdatw[31]_INST_0_i_155_n_0 ;
  wire \bdatw[31]_INST_0_i_156_n_0 ;
  wire \bdatw[31]_INST_0_i_157_n_0 ;
  wire \bdatw[31]_INST_0_i_158_n_0 ;
  wire \bdatw[31]_INST_0_i_159_n_0 ;
  wire \bdatw[31]_INST_0_i_15_n_0 ;
  wire \bdatw[31]_INST_0_i_160_n_0 ;
  wire \bdatw[31]_INST_0_i_161_n_0 ;
  wire \bdatw[31]_INST_0_i_162_n_0 ;
  wire \bdatw[31]_INST_0_i_163_n_0 ;
  wire \bdatw[31]_INST_0_i_164_n_0 ;
  wire \bdatw[31]_INST_0_i_165_n_0 ;
  wire \bdatw[31]_INST_0_i_166_n_0 ;
  wire \bdatw[31]_INST_0_i_167_n_0 ;
  wire \bdatw[31]_INST_0_i_168_n_0 ;
  wire \bdatw[31]_INST_0_i_169_n_0 ;
  wire \bdatw[31]_INST_0_i_16_n_0 ;
  wire \bdatw[31]_INST_0_i_170_n_0 ;
  wire \bdatw[31]_INST_0_i_171_n_0 ;
  wire \bdatw[31]_INST_0_i_172_n_0 ;
  wire \bdatw[31]_INST_0_i_173_n_0 ;
  wire \bdatw[31]_INST_0_i_174_n_0 ;
  wire \bdatw[31]_INST_0_i_17_n_0 ;
  wire \bdatw[31]_INST_0_i_24_n_0 ;
  wire \bdatw[31]_INST_0_i_25_n_0 ;
  wire \bdatw[31]_INST_0_i_26_n_0 ;
  wire \bdatw[31]_INST_0_i_27_n_0 ;
  wire \bdatw[31]_INST_0_i_28_n_0 ;
  wire \bdatw[31]_INST_0_i_30_n_0 ;
  wire \bdatw[31]_INST_0_i_31_n_0 ;
  wire \bdatw[31]_INST_0_i_32_n_0 ;
  wire \bdatw[31]_INST_0_i_33_n_0 ;
  wire \bdatw[31]_INST_0_i_34_n_0 ;
  wire \bdatw[31]_INST_0_i_3_n_0 ;
  wire \bdatw[31]_INST_0_i_41_n_0 ;
  wire \bdatw[31]_INST_0_i_42_n_0 ;
  wire \bdatw[31]_INST_0_i_43_n_0 ;
  wire \bdatw[31]_INST_0_i_44_n_0 ;
  wire \bdatw[31]_INST_0_i_45_n_0 ;
  wire \bdatw[31]_INST_0_i_59_n_0 ;
  wire \bdatw[31]_INST_0_i_62_n_0 ;
  wire \bdatw[31]_INST_0_i_63_n_0 ;
  wire \bdatw[31]_INST_0_i_64_n_0 ;
  wire \bdatw[31]_INST_0_i_65_n_0 ;
  wire \bdatw[31]_INST_0_i_66_n_0 ;
  wire \bdatw[31]_INST_0_i_67_n_0 ;
  wire \bdatw[31]_INST_0_i_68_n_0 ;
  wire \bdatw[31]_INST_0_i_69_n_0 ;
  wire \bdatw[31]_INST_0_i_6_n_0 ;
  wire \bdatw[31]_INST_0_i_70_n_0 ;
  wire \bdatw[31]_INST_0_i_71_n_0 ;
  wire \bdatw[31]_INST_0_i_72_n_0 ;
  wire \bdatw[31]_INST_0_i_73_n_0 ;
  wire \bdatw[31]_INST_0_i_74_n_0 ;
  wire \bdatw[31]_INST_0_i_75_n_0 ;
  wire \bdatw[31]_INST_0_i_76_n_0 ;
  wire \bdatw[31]_INST_0_i_77_n_0 ;
  wire \bdatw[31]_INST_0_i_78_n_0 ;
  wire \bdatw[31]_INST_0_i_79_n_0 ;
  wire \bdatw[31]_INST_0_i_7_n_0 ;
  wire \bdatw[31]_INST_0_i_80_n_0 ;
  wire \bdatw[31]_INST_0_i_81_n_0 ;
  wire \bdatw[31]_INST_0_i_82_n_0 ;
  wire \bdatw[31]_INST_0_i_83_n_0 ;
  wire \bdatw[31]_INST_0_i_84_n_0 ;
  wire \bdatw[31]_INST_0_i_85_n_0 ;
  wire \bdatw[31]_INST_0_i_8_n_0 ;
  wire \bdatw[31]_INST_0_i_96_n_0 ;
  wire \bdatw[31]_INST_0_i_99_n_0 ;
  wire \bdatw[8]_INST_0_i_10_n_0 ;
  wire \bdatw[8]_INST_0_i_1_n_0 ;
  wire \bdatw[8]_INST_0_i_21_n_0 ;
  wire \bdatw[8]_INST_0_i_22_n_0 ;
  wire \bdatw[8]_INST_0_i_4_n_0 ;
  wire \bdatw[8]_INST_0_i_9_n_0 ;
  wire \bdatw[9]_INST_0_i_10_n_0 ;
  wire \bdatw[9]_INST_0_i_11_n_0 ;
  wire \bdatw[9]_INST_0_i_17_n_0 ;
  wire \bdatw[9]_INST_0_i_1_n_0 ;
  wire \bdatw[9]_INST_0_i_4_n_0 ;
  wire \bdatw[9]_INST_0_i_7_n_0 ;
  wire brdy;
  wire [31:0]c0bus;
  wire [31:0]c1bus;
  wire [31:0]cbus_i;
  wire [4:0]ccmd;
  wire \ccmd[0]_INST_0_i_10_n_0 ;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_13_n_0 ;
  wire \ccmd[0]_INST_0_i_14_n_0 ;
  wire \ccmd[0]_INST_0_i_15_n_0 ;
  wire \ccmd[0]_INST_0_i_16_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_19_n_0 ;
  wire \ccmd[0]_INST_0_i_1_n_0 ;
  wire \ccmd[0]_INST_0_i_20_n_0 ;
  wire \ccmd[0]_INST_0_i_21_n_0 ;
  wire \ccmd[0]_INST_0_i_22_n_0 ;
  wire \ccmd[0]_INST_0_i_23_n_0 ;
  wire \ccmd[0]_INST_0_i_24_n_0 ;
  wire \ccmd[0]_INST_0_i_25_n_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_6_n_0 ;
  wire \ccmd[0]_INST_0_i_7_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1]_INST_0_i_10_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_12_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_15_n_0 ;
  wire \ccmd[1]_INST_0_i_16_n_0 ;
  wire \ccmd[1]_INST_0_i_17_n_0 ;
  wire \ccmd[1]_INST_0_i_1_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_6_n_0 ;
  wire \ccmd[1]_INST_0_i_7_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_10_n_0 ;
  wire \ccmd[2]_INST_0_i_11_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_13_n_0 ;
  wire \ccmd[2]_INST_0_i_14_n_0 ;
  wire \ccmd[2]_INST_0_i_15_n_0 ;
  wire \ccmd[2]_INST_0_i_16_n_0 ;
  wire \ccmd[2]_INST_0_i_17_n_0 ;
  wire \ccmd[2]_INST_0_i_18_n_0 ;
  wire \ccmd[2]_INST_0_i_19_n_0 ;
  wire \ccmd[2]_INST_0_i_1_n_0 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_3_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[2]_INST_0_i_7_n_0 ;
  wire \ccmd[2]_INST_0_i_8_n_0 ;
  wire \ccmd[2]_INST_0_i_9_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_12_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_14_n_0 ;
  wire \ccmd[3]_INST_0_i_15_n_0 ;
  wire \ccmd[3]_INST_0_i_16_n_0 ;
  wire \ccmd[3]_INST_0_i_17_n_0 ;
  wire \ccmd[3]_INST_0_i_18_n_0 ;
  wire \ccmd[3]_INST_0_i_19_n_0 ;
  wire \ccmd[3]_INST_0_i_1_n_0 ;
  wire \ccmd[3]_INST_0_i_20_n_0 ;
  wire \ccmd[3]_INST_0_i_21_n_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_8_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire \ccmd[4]_INST_0_i_1_n_0 ;
  wire \ccmd[4]_INST_0_i_2_n_0 ;
  wire \ccmd[4]_INST_0_i_3_n_0 ;
  wire \ccmd[4]_INST_0_i_4_n_0 ;
  wire chg_quo_sgn_i_1__0_n_0;
  wire chg_quo_sgn_i_1_n_0;
  wire chg_quo_sgn_i_2__0_n_0;
  wire chg_quo_sgn_i_2_n_0;
  wire chg_rem_sgn_i_1__0_n_0;
  wire chg_rem_sgn_i_1_n_0;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire [1:0]\ctl0/stat_nx ;
  wire [2:0]\ctl1/stat_nx ;
  wire \ctl1/stat_reg_n_0_[0] ;
  wire \ctl1/stat_reg_n_0_[1] ;
  wire \ctl1/stat_reg_n_0_[2] ;
  wire ctl_bcc_take0_fl_i_1_n_0;
  wire ctl_bcc_take0_fl_i_2_n_0;
  wire ctl_bcc_take1_fl_i_1_n_0;
  wire ctl_fetch0;
  wire ctl_fetch0_fl_i_10_n_0;
  wire ctl_fetch0_fl_i_11_n_0;
  wire ctl_fetch0_fl_i_12_n_0;
  wire ctl_fetch0_fl_i_13_n_0;
  wire ctl_fetch0_fl_i_14_n_0;
  wire ctl_fetch0_fl_i_15_n_0;
  wire ctl_fetch0_fl_i_16_n_0;
  wire ctl_fetch0_fl_i_17_n_0;
  wire ctl_fetch0_fl_i_18_n_0;
  wire ctl_fetch0_fl_i_19_n_0;
  wire ctl_fetch0_fl_i_20_n_0;
  wire ctl_fetch0_fl_i_21_n_0;
  wire ctl_fetch0_fl_i_22_n_0;
  wire ctl_fetch0_fl_i_23_n_0;
  wire ctl_fetch0_fl_i_24_n_0;
  wire ctl_fetch0_fl_i_25_n_0;
  wire ctl_fetch0_fl_i_26_n_0;
  wire ctl_fetch0_fl_i_27_n_0;
  wire ctl_fetch0_fl_i_28_n_0;
  wire ctl_fetch0_fl_i_29_n_0;
  wire ctl_fetch0_fl_i_2_n_0;
  wire ctl_fetch0_fl_i_30_n_0;
  wire ctl_fetch0_fl_i_31_n_0;
  wire ctl_fetch0_fl_i_32_n_0;
  wire ctl_fetch0_fl_i_33_n_0;
  wire ctl_fetch0_fl_i_34_n_0;
  wire ctl_fetch0_fl_i_35_n_0;
  wire ctl_fetch0_fl_i_36_n_0;
  wire ctl_fetch0_fl_i_37_n_0;
  wire ctl_fetch0_fl_i_38_n_0;
  wire ctl_fetch0_fl_i_39_n_0;
  wire ctl_fetch0_fl_i_3_n_0;
  wire ctl_fetch0_fl_i_40_n_0;
  wire ctl_fetch0_fl_i_41_n_0;
  wire ctl_fetch0_fl_i_42_n_0;
  wire ctl_fetch0_fl_i_43_n_0;
  wire ctl_fetch0_fl_i_44_n_0;
  wire ctl_fetch0_fl_i_45_n_0;
  wire ctl_fetch0_fl_i_46_n_0;
  wire ctl_fetch0_fl_i_47_n_0;
  wire ctl_fetch0_fl_i_48_n_0;
  wire ctl_fetch0_fl_i_49_n_0;
  wire ctl_fetch0_fl_i_4_n_0;
  wire ctl_fetch0_fl_i_50_n_0;
  wire ctl_fetch0_fl_i_51_n_0;
  wire ctl_fetch0_fl_i_5_n_0;
  wire ctl_fetch0_fl_i_6_n_0;
  wire ctl_fetch0_fl_i_7_n_0;
  wire ctl_fetch0_fl_i_8_n_0;
  wire ctl_fetch0_fl_i_9_n_0;
  wire ctl_fetch1;
  wire ctl_fetch1_fl_i_10_n_0;
  wire ctl_fetch1_fl_i_11_n_0;
  wire ctl_fetch1_fl_i_12_n_0;
  wire ctl_fetch1_fl_i_13_n_0;
  wire ctl_fetch1_fl_i_14_n_0;
  wire ctl_fetch1_fl_i_15_n_0;
  wire ctl_fetch1_fl_i_16_n_0;
  wire ctl_fetch1_fl_i_17_n_0;
  wire ctl_fetch1_fl_i_18_n_0;
  wire ctl_fetch1_fl_i_19_n_0;
  wire ctl_fetch1_fl_i_20_n_0;
  wire ctl_fetch1_fl_i_21_n_0;
  wire ctl_fetch1_fl_i_22_n_0;
  wire ctl_fetch1_fl_i_23_n_0;
  wire ctl_fetch1_fl_i_24_n_0;
  wire ctl_fetch1_fl_i_25_n_0;
  wire ctl_fetch1_fl_i_26_n_0;
  wire ctl_fetch1_fl_i_27_n_0;
  wire ctl_fetch1_fl_i_28_n_0;
  wire ctl_fetch1_fl_i_29_n_0;
  wire ctl_fetch1_fl_i_30_n_0;
  wire ctl_fetch1_fl_i_31_n_0;
  wire ctl_fetch1_fl_i_32_n_0;
  wire ctl_fetch1_fl_i_33_n_0;
  wire ctl_fetch1_fl_i_34_n_0;
  wire ctl_fetch1_fl_i_35_n_0;
  wire ctl_fetch1_fl_i_36_n_0;
  wire ctl_fetch1_fl_i_37_n_0;
  wire ctl_fetch1_fl_i_38_n_0;
  wire ctl_fetch1_fl_i_39_n_0;
  wire ctl_fetch1_fl_i_3_n_0;
  wire ctl_fetch1_fl_i_40_n_0;
  wire ctl_fetch1_fl_i_41_n_0;
  wire ctl_fetch1_fl_i_42_n_0;
  wire ctl_fetch1_fl_i_43_n_0;
  wire ctl_fetch1_fl_i_44_n_0;
  wire ctl_fetch1_fl_i_45_n_0;
  wire ctl_fetch1_fl_i_46_n_0;
  wire ctl_fetch1_fl_i_47_n_0;
  wire ctl_fetch1_fl_i_48_n_0;
  wire ctl_fetch1_fl_i_4_n_0;
  wire ctl_fetch1_fl_i_5_n_0;
  wire ctl_fetch1_fl_i_6_n_0;
  wire ctl_fetch1_fl_i_7_n_0;
  wire ctl_fetch1_fl_i_8_n_0;
  wire ctl_fetch1_fl_i_9_n_0;
  wire ctl_fetch1_fl_reg_i_2_n_0;
  wire ctl_fetch_ext0;
  wire ctl_fetch_ext1;
  wire ctl_fetch_lng0;
  wire ctl_fetch_lng1;
  wire [0:0]ctl_sela0;
  wire [1:1]ctl_sela0_rn;
  wire [0:0]ctl_sela1;
  wire [1:1]ctl_selb0_0;
  wire [2:0]ctl_selb0_rn;
  wire [2:1]ctl_selb1_0;
  wire [2:0]ctl_selb1_rn;
  wire [1:0]ctl_selc0;
  wire [0:0]ctl_selc0_rn;
  wire [1:0]ctl_selc1;
  wire [0:0]ctl_selc1_rn;
  wire ctl_sp_dec1;
  wire ctl_sp_id40;
  wire ctl_sp_inc0;
  wire ctl_sr_ldie0;
  wire ctl_sr_ldie1;
  wire ctl_sr_upd0;
  wire ctl_sr_upd1;
  wire dctl_sign_f_i_10_n_0;
  wire dctl_sign_f_i_11_n_0;
  wire dctl_sign_f_i_12_n_0;
  wire dctl_sign_f_i_13_n_0;
  wire dctl_sign_f_i_14_n_0;
  wire dctl_sign_f_i_2_n_0;
  wire dctl_sign_f_i_3_n_0;
  wire dctl_sign_f_i_4_n_0;
  wire dctl_sign_f_i_5_n_0;
  wire dctl_sign_f_i_6_n_0;
  wire dctl_sign_f_i_7_n_0;
  wire dctl_sign_f_i_8_n_0;
  wire dctl_sign_f_i_9_n_0;
  wire \dctl_stat[0]_i_2__0_n_0 ;
  wire \dctl_stat[0]_i_2_n_0 ;
  wire \dctl_stat[0]_i_3__0_n_0 ;
  wire \dctl_stat[0]_i_3_n_0 ;
  wire \dctl_stat[1]_i_2__0_n_0 ;
  wire \dctl_stat[1]_i_2_n_0 ;
  wire \dctl_stat[1]_i_3__0_n_0 ;
  wire \dctl_stat[1]_i_3_n_0 ;
  wire \dctl_stat[2]_i_2__0_n_0 ;
  wire \dctl_stat[2]_i_2_n_0 ;
  wire \dctl_stat[3]_i_2__0_n_0 ;
  wire \dctl_stat[3]_i_2_n_0 ;
  wire \dctl_stat[3]_i_4__0_n_0 ;
  wire \dctl_stat[3]_i_4_n_0 ;
  wire \dctl_stat[3]_i_5__0_n_0 ;
  wire \dctl_stat[3]_i_5_n_0 ;
  wire div_crdy0;
  wire div_crdy1;
  wire div_crdy_i_1__0_n_0;
  wire div_crdy_i_1_n_0;
  wire div_crdy_i_2__0_n_0;
  wire div_crdy_i_2_n_0;
  wire div_crdy_i_3__0_n_0;
  wire div_crdy_i_3_n_0;
  wire div_crdy_i_4__0_n_0;
  wire div_crdy_i_4_n_0;
  wire \dso[11]_i_10__0_n_0 ;
  wire \dso[11]_i_10_n_0 ;
  wire \dso[11]_i_11__0_n_0 ;
  wire \dso[11]_i_11_n_0 ;
  wire \dso[11]_i_12__0_n_0 ;
  wire \dso[11]_i_12_n_0 ;
  wire \dso[11]_i_13__0_n_0 ;
  wire \dso[11]_i_13_n_0 ;
  wire \dso[11]_i_2__0_n_0 ;
  wire \dso[11]_i_2_n_0 ;
  wire \dso[11]_i_3__0_n_0 ;
  wire \dso[11]_i_3_n_0 ;
  wire \dso[11]_i_4__0_n_0 ;
  wire \dso[11]_i_4_n_0 ;
  wire \dso[11]_i_5__0_n_0 ;
  wire \dso[11]_i_5_n_0 ;
  wire \dso[11]_i_6__0_n_0 ;
  wire \dso[11]_i_6_n_0 ;
  wire \dso[11]_i_7__0_n_0 ;
  wire \dso[11]_i_7_n_0 ;
  wire \dso[11]_i_8__0_n_0 ;
  wire \dso[11]_i_8_n_0 ;
  wire \dso[11]_i_9__0_n_0 ;
  wire \dso[11]_i_9_n_0 ;
  wire \dso[15]_i_10__0_n_0 ;
  wire \dso[15]_i_10_n_0 ;
  wire \dso[15]_i_11__0_n_0 ;
  wire \dso[15]_i_11_n_0 ;
  wire \dso[15]_i_12__0_n_0 ;
  wire \dso[15]_i_12_n_0 ;
  wire \dso[15]_i_13__0_n_0 ;
  wire \dso[15]_i_13_n_0 ;
  wire \dso[15]_i_14__0_n_0 ;
  wire \dso[15]_i_14_n_0 ;
  wire \dso[15]_i_2__0_n_0 ;
  wire \dso[15]_i_2_n_0 ;
  wire \dso[15]_i_3__0_n_0 ;
  wire \dso[15]_i_3_n_0 ;
  wire \dso[15]_i_4__0_n_0 ;
  wire \dso[15]_i_4_n_0 ;
  wire \dso[15]_i_5__0_n_0 ;
  wire \dso[15]_i_5_n_0 ;
  wire \dso[15]_i_6__0_n_0 ;
  wire \dso[15]_i_6_n_0 ;
  wire \dso[15]_i_7__0_n_0 ;
  wire \dso[15]_i_7_n_0 ;
  wire \dso[15]_i_8__0_n_0 ;
  wire \dso[15]_i_8_n_0 ;
  wire \dso[15]_i_9__0_n_0 ;
  wire \dso[15]_i_9_n_0 ;
  wire \dso[19]_i_10__0_n_0 ;
  wire \dso[19]_i_10_n_0 ;
  wire \dso[19]_i_11__0_n_0 ;
  wire \dso[19]_i_11_n_0 ;
  wire \dso[19]_i_12__0_n_0 ;
  wire \dso[19]_i_12_n_0 ;
  wire \dso[19]_i_13__0_n_0 ;
  wire \dso[19]_i_13_n_0 ;
  wire \dso[19]_i_2__0_n_0 ;
  wire \dso[19]_i_2_n_0 ;
  wire \dso[19]_i_3__0_n_0 ;
  wire \dso[19]_i_3_n_0 ;
  wire \dso[19]_i_4__0_n_0 ;
  wire \dso[19]_i_4_n_0 ;
  wire \dso[19]_i_5__0_n_0 ;
  wire \dso[19]_i_5_n_0 ;
  wire \dso[19]_i_6__0_n_0 ;
  wire \dso[19]_i_6_n_0 ;
  wire \dso[19]_i_7__0_n_0 ;
  wire \dso[19]_i_7_n_0 ;
  wire \dso[19]_i_8__0_n_0 ;
  wire \dso[19]_i_8_n_0 ;
  wire \dso[19]_i_9__0_n_0 ;
  wire \dso[19]_i_9_n_0 ;
  wire \dso[23]_i_10__0_n_0 ;
  wire \dso[23]_i_10_n_0 ;
  wire \dso[23]_i_11__0_n_0 ;
  wire \dso[23]_i_11_n_0 ;
  wire \dso[23]_i_12__0_n_0 ;
  wire \dso[23]_i_12_n_0 ;
  wire \dso[23]_i_13__0_n_0 ;
  wire \dso[23]_i_13_n_0 ;
  wire \dso[23]_i_2__0_n_0 ;
  wire \dso[23]_i_2_n_0 ;
  wire \dso[23]_i_3__0_n_0 ;
  wire \dso[23]_i_3_n_0 ;
  wire \dso[23]_i_4__0_n_0 ;
  wire \dso[23]_i_4_n_0 ;
  wire \dso[23]_i_5__0_n_0 ;
  wire \dso[23]_i_5_n_0 ;
  wire \dso[23]_i_6__0_n_0 ;
  wire \dso[23]_i_6_n_0 ;
  wire \dso[23]_i_7__0_n_0 ;
  wire \dso[23]_i_7_n_0 ;
  wire \dso[23]_i_8__0_n_0 ;
  wire \dso[23]_i_8_n_0 ;
  wire \dso[23]_i_9__0_n_0 ;
  wire \dso[23]_i_9_n_0 ;
  wire \dso[27]_i_10__0_n_0 ;
  wire \dso[27]_i_10_n_0 ;
  wire \dso[27]_i_11__0_n_0 ;
  wire \dso[27]_i_11_n_0 ;
  wire \dso[27]_i_12__0_n_0 ;
  wire \dso[27]_i_12_n_0 ;
  wire \dso[27]_i_13__0_n_0 ;
  wire \dso[27]_i_13_n_0 ;
  wire \dso[27]_i_2__0_n_0 ;
  wire \dso[27]_i_2_n_0 ;
  wire \dso[27]_i_3__0_n_0 ;
  wire \dso[27]_i_3_n_0 ;
  wire \dso[27]_i_4__0_n_0 ;
  wire \dso[27]_i_4_n_0 ;
  wire \dso[27]_i_5__0_n_0 ;
  wire \dso[27]_i_5_n_0 ;
  wire \dso[27]_i_6__0_n_0 ;
  wire \dso[27]_i_6_n_0 ;
  wire \dso[27]_i_7__0_n_0 ;
  wire \dso[27]_i_7_n_0 ;
  wire \dso[27]_i_8__0_n_0 ;
  wire \dso[27]_i_8_n_0 ;
  wire \dso[27]_i_9__0_n_0 ;
  wire \dso[27]_i_9_n_0 ;
  wire \dso[31]_i_10__0_n_0 ;
  wire \dso[31]_i_10_n_0 ;
  wire \dso[31]_i_11__0_n_0 ;
  wire \dso[31]_i_11_n_0 ;
  wire \dso[31]_i_12__0_n_0 ;
  wire \dso[31]_i_12_n_0 ;
  wire \dso[31]_i_13__0_n_0 ;
  wire \dso[31]_i_13_n_0 ;
  wire \dso[31]_i_14__0_n_0 ;
  wire \dso[31]_i_14_n_0 ;
  wire \dso[31]_i_15__0_n_0 ;
  wire \dso[31]_i_15_n_0 ;
  wire \dso[31]_i_17__0_n_0 ;
  wire \dso[31]_i_17_n_0 ;
  wire \dso[31]_i_18__0_n_0 ;
  wire \dso[31]_i_18_n_0 ;
  wire \dso[31]_i_19__0_n_0 ;
  wire \dso[31]_i_19_n_0 ;
  wire \dso[31]_i_1__0_n_0 ;
  wire \dso[31]_i_1_n_0 ;
  wire \dso[31]_i_20__0_n_0 ;
  wire \dso[31]_i_20_n_0 ;
  wire \dso[31]_i_21__0_n_0 ;
  wire \dso[31]_i_21_n_0 ;
  wire \dso[31]_i_3__0_n_0 ;
  wire \dso[31]_i_3_n_0 ;
  wire \dso[31]_i_4__0_n_0 ;
  wire \dso[31]_i_4_n_0 ;
  wire \dso[31]_i_5__0_n_0 ;
  wire \dso[31]_i_5_n_0 ;
  wire \dso[31]_i_6__0_n_0 ;
  wire \dso[31]_i_6_n_0 ;
  wire \dso[31]_i_7__0_n_0 ;
  wire \dso[31]_i_7_n_0 ;
  wire \dso[31]_i_8__0_n_0 ;
  wire \dso[31]_i_8_n_0 ;
  wire \dso[31]_i_9__0_n_0 ;
  wire \dso[31]_i_9_n_0 ;
  wire \dso[3]_i_10__0_n_0 ;
  wire \dso[3]_i_10_n_0 ;
  wire \dso[3]_i_11__0_n_0 ;
  wire \dso[3]_i_11_n_0 ;
  wire \dso[3]_i_12__0_n_0 ;
  wire \dso[3]_i_12_n_0 ;
  wire \dso[3]_i_13__0_n_0 ;
  wire \dso[3]_i_13_n_0 ;
  wire \dso[3]_i_2__0_n_0 ;
  wire \dso[3]_i_2_n_0 ;
  wire \dso[3]_i_3__0_n_0 ;
  wire \dso[3]_i_3_n_0 ;
  wire \dso[3]_i_4__0_n_0 ;
  wire \dso[3]_i_4_n_0 ;
  wire \dso[3]_i_5__0_n_0 ;
  wire \dso[3]_i_5_n_0 ;
  wire \dso[3]_i_6__0_n_0 ;
  wire \dso[3]_i_6_n_0 ;
  wire \dso[3]_i_7__0_n_0 ;
  wire \dso[3]_i_7_n_0 ;
  wire \dso[3]_i_8__0_n_0 ;
  wire \dso[3]_i_8_n_0 ;
  wire \dso[3]_i_9__0_n_0 ;
  wire \dso[3]_i_9_n_0 ;
  wire \dso[7]_i_10__0_n_0 ;
  wire \dso[7]_i_10_n_0 ;
  wire \dso[7]_i_11__0_n_0 ;
  wire \dso[7]_i_11_n_0 ;
  wire \dso[7]_i_12__0_n_0 ;
  wire \dso[7]_i_12_n_0 ;
  wire \dso[7]_i_13__0_n_0 ;
  wire \dso[7]_i_13_n_0 ;
  wire \dso[7]_i_2__0_n_0 ;
  wire \dso[7]_i_2_n_0 ;
  wire \dso[7]_i_3__0_n_0 ;
  wire \dso[7]_i_3_n_0 ;
  wire \dso[7]_i_4__0_n_0 ;
  wire \dso[7]_i_4_n_0 ;
  wire \dso[7]_i_5__0_n_0 ;
  wire \dso[7]_i_5_n_0 ;
  wire \dso[7]_i_6__0_n_0 ;
  wire \dso[7]_i_6_n_0 ;
  wire \dso[7]_i_7__0_n_0 ;
  wire \dso[7]_i_7_n_0 ;
  wire \dso[7]_i_8__0_n_0 ;
  wire \dso[7]_i_8_n_0 ;
  wire \dso[7]_i_9__0_n_0 ;
  wire \dso[7]_i_9_n_0 ;
  wire \dso_reg[11]_i_1__0_n_0 ;
  wire \dso_reg[11]_i_1__0_n_1 ;
  wire \dso_reg[11]_i_1__0_n_2 ;
  wire \dso_reg[11]_i_1__0_n_3 ;
  wire \dso_reg[11]_i_1__0_n_4 ;
  wire \dso_reg[11]_i_1__0_n_5 ;
  wire \dso_reg[11]_i_1__0_n_6 ;
  wire \dso_reg[11]_i_1__0_n_7 ;
  wire \dso_reg[11]_i_1_n_0 ;
  wire \dso_reg[11]_i_1_n_1 ;
  wire \dso_reg[11]_i_1_n_2 ;
  wire \dso_reg[11]_i_1_n_3 ;
  wire \dso_reg[11]_i_1_n_4 ;
  wire \dso_reg[11]_i_1_n_5 ;
  wire \dso_reg[11]_i_1_n_6 ;
  wire \dso_reg[11]_i_1_n_7 ;
  wire \dso_reg[15]_i_1__0_n_0 ;
  wire \dso_reg[15]_i_1__0_n_1 ;
  wire \dso_reg[15]_i_1__0_n_2 ;
  wire \dso_reg[15]_i_1__0_n_3 ;
  wire \dso_reg[15]_i_1__0_n_4 ;
  wire \dso_reg[15]_i_1__0_n_5 ;
  wire \dso_reg[15]_i_1__0_n_6 ;
  wire \dso_reg[15]_i_1__0_n_7 ;
  wire \dso_reg[15]_i_1_n_0 ;
  wire \dso_reg[15]_i_1_n_1 ;
  wire \dso_reg[15]_i_1_n_2 ;
  wire \dso_reg[15]_i_1_n_3 ;
  wire \dso_reg[15]_i_1_n_4 ;
  wire \dso_reg[15]_i_1_n_5 ;
  wire \dso_reg[15]_i_1_n_6 ;
  wire \dso_reg[15]_i_1_n_7 ;
  wire \dso_reg[19]_i_1__0_n_0 ;
  wire \dso_reg[19]_i_1__0_n_1 ;
  wire \dso_reg[19]_i_1__0_n_2 ;
  wire \dso_reg[19]_i_1__0_n_3 ;
  wire \dso_reg[19]_i_1__0_n_4 ;
  wire \dso_reg[19]_i_1__0_n_5 ;
  wire \dso_reg[19]_i_1__0_n_6 ;
  wire \dso_reg[19]_i_1__0_n_7 ;
  wire \dso_reg[19]_i_1_n_0 ;
  wire \dso_reg[19]_i_1_n_1 ;
  wire \dso_reg[19]_i_1_n_2 ;
  wire \dso_reg[19]_i_1_n_3 ;
  wire \dso_reg[19]_i_1_n_4 ;
  wire \dso_reg[19]_i_1_n_5 ;
  wire \dso_reg[19]_i_1_n_6 ;
  wire \dso_reg[19]_i_1_n_7 ;
  wire \dso_reg[23]_i_1__0_n_0 ;
  wire \dso_reg[23]_i_1__0_n_1 ;
  wire \dso_reg[23]_i_1__0_n_2 ;
  wire \dso_reg[23]_i_1__0_n_3 ;
  wire \dso_reg[23]_i_1__0_n_4 ;
  wire \dso_reg[23]_i_1__0_n_5 ;
  wire \dso_reg[23]_i_1__0_n_6 ;
  wire \dso_reg[23]_i_1__0_n_7 ;
  wire \dso_reg[23]_i_1_n_0 ;
  wire \dso_reg[23]_i_1_n_1 ;
  wire \dso_reg[23]_i_1_n_2 ;
  wire \dso_reg[23]_i_1_n_3 ;
  wire \dso_reg[23]_i_1_n_4 ;
  wire \dso_reg[23]_i_1_n_5 ;
  wire \dso_reg[23]_i_1_n_6 ;
  wire \dso_reg[23]_i_1_n_7 ;
  wire \dso_reg[27]_i_1__0_n_0 ;
  wire \dso_reg[27]_i_1__0_n_1 ;
  wire \dso_reg[27]_i_1__0_n_2 ;
  wire \dso_reg[27]_i_1__0_n_3 ;
  wire \dso_reg[27]_i_1__0_n_4 ;
  wire \dso_reg[27]_i_1__0_n_5 ;
  wire \dso_reg[27]_i_1__0_n_6 ;
  wire \dso_reg[27]_i_1__0_n_7 ;
  wire \dso_reg[27]_i_1_n_0 ;
  wire \dso_reg[27]_i_1_n_1 ;
  wire \dso_reg[27]_i_1_n_2 ;
  wire \dso_reg[27]_i_1_n_3 ;
  wire \dso_reg[27]_i_1_n_4 ;
  wire \dso_reg[27]_i_1_n_5 ;
  wire \dso_reg[27]_i_1_n_6 ;
  wire \dso_reg[27]_i_1_n_7 ;
  wire \dso_reg[31]_i_2__0_n_1 ;
  wire \dso_reg[31]_i_2__0_n_2 ;
  wire \dso_reg[31]_i_2__0_n_3 ;
  wire \dso_reg[31]_i_2__0_n_4 ;
  wire \dso_reg[31]_i_2__0_n_5 ;
  wire \dso_reg[31]_i_2__0_n_6 ;
  wire \dso_reg[31]_i_2__0_n_7 ;
  wire \dso_reg[31]_i_2_n_1 ;
  wire \dso_reg[31]_i_2_n_2 ;
  wire \dso_reg[31]_i_2_n_3 ;
  wire \dso_reg[31]_i_2_n_4 ;
  wire \dso_reg[31]_i_2_n_5 ;
  wire \dso_reg[31]_i_2_n_6 ;
  wire \dso_reg[31]_i_2_n_7 ;
  wire \dso_reg[3]_i_1__0_n_0 ;
  wire \dso_reg[3]_i_1__0_n_1 ;
  wire \dso_reg[3]_i_1__0_n_2 ;
  wire \dso_reg[3]_i_1__0_n_3 ;
  wire \dso_reg[3]_i_1__0_n_4 ;
  wire \dso_reg[3]_i_1__0_n_5 ;
  wire \dso_reg[3]_i_1__0_n_6 ;
  wire \dso_reg[3]_i_1__0_n_7 ;
  wire \dso_reg[3]_i_1_n_0 ;
  wire \dso_reg[3]_i_1_n_1 ;
  wire \dso_reg[3]_i_1_n_2 ;
  wire \dso_reg[3]_i_1_n_3 ;
  wire \dso_reg[3]_i_1_n_4 ;
  wire \dso_reg[3]_i_1_n_5 ;
  wire \dso_reg[3]_i_1_n_6 ;
  wire \dso_reg[3]_i_1_n_7 ;
  wire \dso_reg[7]_i_1__0_n_0 ;
  wire \dso_reg[7]_i_1__0_n_1 ;
  wire \dso_reg[7]_i_1__0_n_2 ;
  wire \dso_reg[7]_i_1__0_n_3 ;
  wire \dso_reg[7]_i_1__0_n_4 ;
  wire \dso_reg[7]_i_1__0_n_5 ;
  wire \dso_reg[7]_i_1__0_n_6 ;
  wire \dso_reg[7]_i_1__0_n_7 ;
  wire \dso_reg[7]_i_1_n_0 ;
  wire \dso_reg[7]_i_1_n_1 ;
  wire \dso_reg[7]_i_1_n_2 ;
  wire \dso_reg[7]_i_1_n_3 ;
  wire \dso_reg[7]_i_1_n_4 ;
  wire \dso_reg[7]_i_1_n_5 ;
  wire \dso_reg[7]_i_1_n_6 ;
  wire \dso_reg[7]_i_1_n_7 ;
  wire \eir_fl[1]_i_1_n_0 ;
  wire \eir_fl[2]_i_1_n_0 ;
  wire \eir_fl[31]_i_1_n_0 ;
  wire \eir_fl[3]_i_1_n_0 ;
  wire \eir_fl[4]_i_1_n_0 ;
  wire \eir_fl[5]_i_1_n_0 ;
  wire \eir_fl[6]_i_1_n_0 ;
  wire eir_inferred_i_33_n_0;
  wire eir_inferred_i_34_n_0;
  wire eir_inferred_i_35_n_0;
  wire eir_inferred_i_36_n_0;
  wire eir_inferred_i_37_n_0;
  wire eir_inferred_i_38_n_0;
  wire eir_inferred_i_39_n_0;
  wire eir_inferred_i_40_n_0;
  wire eir_inferred_i_41_n_0;
  wire eir_inferred_i_42_n_0;
  wire eir_inferred_i_43_n_0;
  wire eir_inferred_i_44_n_0;
  wire eir_inferred_i_45_n_0;
  wire eir_inferred_i_46_n_0;
  wire eir_inferred_i_47_n_0;
  wire eir_inferred_i_48_n_0;
  wire eir_inferred_i_49_n_0;
  wire eir_inferred_i_50_n_0;
  wire eir_inferred_i_51_n_0;
  wire eir_inferred_i_52_n_0;
  wire eir_inferred_i_53_n_0;
  wire eir_inferred_i_54_n_0;
  wire eir_inferred_i_55_n_0;
  wire eir_inferred_i_56_n_0;
  wire eir_inferred_i_57_n_0;
  wire eir_inferred_i_58_n_0;
  wire eir_inferred_i_59_n_0;
  wire eir_inferred_i_60_n_0;
  wire eir_inferred_i_61_n_0;
  wire eir_inferred_i_62_n_0;
  wire eir_inferred_i_63_n_0;
  wire eir_inferred_i_64_n_0;
  wire eir_inferred_i_65_n_0;
  wire eir_inferred_i_66_n_0;
  wire eir_inferred_i_67_n_0;
  wire eir_inferred_i_68_n_0;
  wire eir_inferred_i_69_n_0;
  wire eir_inferred_i_70_n_0;
  wire eir_inferred_i_71_n_0;
  wire eir_inferred_i_72_n_0;
  wire eir_inferred_i_73_n_0;
  wire eir_inferred_i_74_n_0;
  wire eir_inferred_i_75_n_0;
  wire eir_inferred_i_76_n_0;
  wire eir_inferred_i_77_n_0;
  wire eir_inferred_i_78_n_0;
  wire eir_inferred_i_79_n_0;
  wire eir_inferred_i_80_n_0;
  wire eir_inferred_i_81_n_0;
  wire eir_inferred_i_82_n_0;
  wire eir_inferred_i_83_n_0;
  wire eir_inferred_i_84_n_0;
  wire eir_inferred_i_85_n_0;
  wire eir_inferred_i_86_n_0;
  wire eir_inferred_i_87_n_0;
  wire eir_inferred_i_88_n_0;
  wire eir_inferred_i_89_n_0;
  wire [15:1]\^fadr ;
  wire \fadr[11]_INST_0_i_1_n_0 ;
  wire \fadr[11]_INST_0_i_1_n_1 ;
  wire \fadr[11]_INST_0_i_1_n_2 ;
  wire \fadr[11]_INST_0_i_1_n_3 ;
  wire \fadr[12]_INST_0_i_1_n_0 ;
  wire \fadr[12]_INST_0_i_1_n_1 ;
  wire \fadr[12]_INST_0_i_1_n_2 ;
  wire \fadr[12]_INST_0_i_1_n_3 ;
  wire \fadr[12]_INST_0_i_1_n_4 ;
  wire \fadr[12]_INST_0_i_1_n_5 ;
  wire \fadr[12]_INST_0_i_1_n_6 ;
  wire \fadr[12]_INST_0_i_1_n_7 ;
  wire \fadr[15]_INST_0_i_10_n_0 ;
  wire \fadr[15]_INST_0_i_11_n_0 ;
  wire \fadr[15]_INST_0_i_12_n_0 ;
  wire \fadr[15]_INST_0_i_13_n_0 ;
  wire \fadr[15]_INST_0_i_14_n_0 ;
  wire \fadr[15]_INST_0_i_15_n_0 ;
  wire \fadr[15]_INST_0_i_16_n_0 ;
  wire \fadr[15]_INST_0_i_17_n_0 ;
  wire \fadr[15]_INST_0_i_1_n_1 ;
  wire \fadr[15]_INST_0_i_1_n_2 ;
  wire \fadr[15]_INST_0_i_1_n_3 ;
  wire \fadr[15]_INST_0_i_2_n_0 ;
  wire \fadr[15]_INST_0_i_3_n_0 ;
  wire \fadr[15]_INST_0_i_4_n_2 ;
  wire \fadr[15]_INST_0_i_4_n_3 ;
  wire \fadr[15]_INST_0_i_4_n_5 ;
  wire \fadr[15]_INST_0_i_4_n_6 ;
  wire \fadr[15]_INST_0_i_4_n_7 ;
  wire \fadr[15]_INST_0_i_5_n_0 ;
  wire \fadr[15]_INST_0_i_6_n_0 ;
  wire \fadr[15]_INST_0_i_7_n_0 ;
  wire \fadr[15]_INST_0_i_8_n_0 ;
  wire \fadr[15]_INST_0_i_9_n_0 ;
  wire \fadr[3]_INST_0_i_1_n_0 ;
  wire \fadr[3]_INST_0_i_1_n_1 ;
  wire \fadr[3]_INST_0_i_1_n_2 ;
  wire \fadr[3]_INST_0_i_1_n_3 ;
  wire \fadr[3]_INST_0_i_2_n_0 ;
  wire \fadr[4]_INST_0_i_1_n_0 ;
  wire \fadr[4]_INST_0_i_1_n_1 ;
  wire \fadr[4]_INST_0_i_1_n_2 ;
  wire \fadr[4]_INST_0_i_1_n_3 ;
  wire \fadr[4]_INST_0_i_1_n_4 ;
  wire \fadr[4]_INST_0_i_1_n_5 ;
  wire \fadr[4]_INST_0_i_1_n_6 ;
  wire \fadr[4]_INST_0_i_1_n_7 ;
  wire \fadr[4]_INST_0_i_2_n_0 ;
  wire \fadr[7]_INST_0_i_1_n_0 ;
  wire \fadr[7]_INST_0_i_1_n_1 ;
  wire \fadr[7]_INST_0_i_1_n_2 ;
  wire \fadr[7]_INST_0_i_1_n_3 ;
  wire \fadr[8]_INST_0_i_1_n_0 ;
  wire \fadr[8]_INST_0_i_1_n_1 ;
  wire \fadr[8]_INST_0_i_1_n_2 ;
  wire \fadr[8]_INST_0_i_1_n_3 ;
  wire \fadr[8]_INST_0_i_1_n_4 ;
  wire \fadr[8]_INST_0_i_1_n_5 ;
  wire \fadr[8]_INST_0_i_1_n_6 ;
  wire \fadr[8]_INST_0_i_1_n_7 ;
  wire \fch/ctl_bcc_take0_fl ;
  wire \fch/ctl_bcc_take1_fl ;
  wire \fch/ctl_fetch0_fl ;
  wire \fch/ctl_fetch1_fl ;
  wire \fch/ctl_fetch_ext ;
  wire \fch/ctl_fetch_ext_fl ;
  wire \fch/ctl_fetch_lng ;
  wire \fch/ctl_fetch_lng_fl ;
  wire [31:0]\fch/data0 ;
  (* DONT_TOUCH *) wire [31:0]\fch/eir ;
  wire \fch/eir_fl_reg_n_0_[16] ;
  wire \fch/eir_fl_reg_n_0_[17] ;
  wire \fch/eir_fl_reg_n_0_[18] ;
  wire \fch/eir_fl_reg_n_0_[19] ;
  wire \fch/eir_fl_reg_n_0_[20] ;
  wire \fch/eir_fl_reg_n_0_[21] ;
  wire \fch/eir_fl_reg_n_0_[22] ;
  wire \fch/eir_fl_reg_n_0_[23] ;
  wire \fch/eir_fl_reg_n_0_[24] ;
  wire \fch/eir_fl_reg_n_0_[25] ;
  wire \fch/eir_fl_reg_n_0_[26] ;
  wire \fch/eir_fl_reg_n_0_[27] ;
  wire \fch/eir_fl_reg_n_0_[28] ;
  wire \fch/eir_fl_reg_n_0_[29] ;
  wire \fch/eir_fl_reg_n_0_[30] ;
  wire \fch/eir_fl_reg_n_0_[31] ;
  wire \fch/fadr_1_fl ;
  wire \fch/fch_heir_hir ;
  wire \fch/fch_heir_nir ;
  wire \fch/fch_irq_req_fl ;
  (* DONT_TOUCH *) wire \fch/fch_issu1 ;
  wire \fch/fch_issu1_fl ;
  wire \fch/fch_issu1_ir ;
  wire \fch/fch_leir_hir ;
  wire \fch/fch_leir_lir ;
  wire \fch/fch_leir_nir ;
  wire \fch/fch_term_fl ;
  wire \fch/fctl/fch_heir_hir_t ;
  wire \fch/fctl/fch_heir_nir_t ;
  wire \fch/fctl/fch_leir_hir_t ;
  wire \fch/fctl/fch_leir_lir_t ;
  wire \fch/fctl/fch_leir_nir_t ;
  wire \fch/fctl/fch_nir_lir ;
  wire [2:0]\fch/fctl/stat_nx ;
  (* DONT_TOUCH *) wire [15:0]\fch/ir0 ;
  wire [15:0]\fch/ir0_fl ;
  wire [21:20]\fch/ir0_id_fl ;
  (* DONT_TOUCH *) wire [15:0]\fch/ir1 ;
  wire [15:0]\fch/ir1_fl ;
  wire [21:20]\fch/ir1_id_fl ;
  wire [24:12]\fch/lir_id_0 ;
  wire [24:12]\fch/nir_id ;
  wire [15:1]\fch/p_2_in ;
  wire [15:0]\fch/p_2_in0_in ;
  wire \fch/rst_n_fl ;
  wire [2:0]\fch/stat ;
  wire fch_heir_nir_i_2_n_0;
  wire fch_heir_nir_i_3_n_0;
  wire fch_heir_nir_i_6_n_0;
  wire fch_heir_nir_i_7_n_0;
  wire fch_heir_nir_i_8_n_0;
  wire [1:0]fch_irq_lev;
  wire \fch_irq_lev[0]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_2_n_0 ;
  wire \fch_irq_lev[1]_i_3_n_0 ;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev[1]_i_5_n_0 ;
  wire \fch_irq_lev[1]_i_6_n_0 ;
  wire \fch_irq_lev[1]_i_7_n_0 ;
  wire \fch_irq_lev[1]_i_8_n_0 ;
  wire \fch_irq_lev[1]_i_9_n_0 ;
  wire fch_irq_req;
  wire fch_issu1_inferred_i_100_n_0;
  wire fch_issu1_inferred_i_101_n_0;
  wire fch_issu1_inferred_i_102_n_0;
  wire fch_issu1_inferred_i_103_n_0;
  wire fch_issu1_inferred_i_104_n_0;
  wire fch_issu1_inferred_i_105_n_0;
  wire fch_issu1_inferred_i_106_n_0;
  wire fch_issu1_inferred_i_107_n_0;
  wire fch_issu1_inferred_i_108_n_0;
  wire fch_issu1_inferred_i_109_n_0;
  wire fch_issu1_inferred_i_10_n_0;
  wire fch_issu1_inferred_i_110_n_0;
  wire fch_issu1_inferred_i_111_n_0;
  wire fch_issu1_inferred_i_112_n_0;
  wire fch_issu1_inferred_i_113_n_0;
  wire fch_issu1_inferred_i_114_n_0;
  wire fch_issu1_inferred_i_115_n_0;
  wire fch_issu1_inferred_i_116_n_0;
  wire fch_issu1_inferred_i_117_n_0;
  wire fch_issu1_inferred_i_118_n_0;
  wire fch_issu1_inferred_i_119_n_0;
  wire fch_issu1_inferred_i_11_n_0;
  wire fch_issu1_inferred_i_120_n_0;
  wire fch_issu1_inferred_i_121_n_0;
  wire fch_issu1_inferred_i_122_n_0;
  wire fch_issu1_inferred_i_123_n_0;
  wire fch_issu1_inferred_i_124_n_0;
  wire fch_issu1_inferred_i_125_n_0;
  wire fch_issu1_inferred_i_126_n_0;
  wire fch_issu1_inferred_i_127_n_0;
  wire fch_issu1_inferred_i_128_n_0;
  wire fch_issu1_inferred_i_129_n_0;
  wire fch_issu1_inferred_i_12_n_0;
  wire fch_issu1_inferred_i_130_n_0;
  wire fch_issu1_inferred_i_131_n_0;
  wire fch_issu1_inferred_i_132_n_0;
  wire fch_issu1_inferred_i_133_n_0;
  wire fch_issu1_inferred_i_134_n_0;
  wire fch_issu1_inferred_i_135_n_0;
  wire fch_issu1_inferred_i_136_n_0;
  wire fch_issu1_inferred_i_137_n_0;
  wire fch_issu1_inferred_i_138_n_0;
  wire fch_issu1_inferred_i_139_n_0;
  wire fch_issu1_inferred_i_13_n_0;
  wire fch_issu1_inferred_i_140_n_0;
  wire fch_issu1_inferred_i_141_n_0;
  wire fch_issu1_inferred_i_142_n_0;
  wire fch_issu1_inferred_i_143_n_0;
  wire fch_issu1_inferred_i_144_n_0;
  wire fch_issu1_inferred_i_145_n_0;
  wire fch_issu1_inferred_i_146_n_0;
  wire fch_issu1_inferred_i_147_n_0;
  wire fch_issu1_inferred_i_148_n_0;
  wire fch_issu1_inferred_i_149_n_0;
  wire fch_issu1_inferred_i_14_n_0;
  wire fch_issu1_inferred_i_150_n_0;
  wire fch_issu1_inferred_i_151_n_0;
  wire fch_issu1_inferred_i_152_n_0;
  wire fch_issu1_inferred_i_153_n_0;
  wire fch_issu1_inferred_i_154_n_0;
  wire fch_issu1_inferred_i_155_n_0;
  wire fch_issu1_inferred_i_156_n_0;
  wire fch_issu1_inferred_i_157_n_0;
  wire fch_issu1_inferred_i_158_n_0;
  wire fch_issu1_inferred_i_159_n_0;
  wire fch_issu1_inferred_i_15_n_0;
  wire fch_issu1_inferred_i_160_n_0;
  wire fch_issu1_inferred_i_161_n_0;
  wire fch_issu1_inferred_i_162_n_0;
  wire fch_issu1_inferred_i_163_n_0;
  wire fch_issu1_inferred_i_164_n_0;
  wire fch_issu1_inferred_i_165_n_0;
  wire fch_issu1_inferred_i_166_n_0;
  wire fch_issu1_inferred_i_167_n_0;
  wire fch_issu1_inferred_i_168_n_0;
  wire fch_issu1_inferred_i_169_n_0;
  wire fch_issu1_inferred_i_16_n_0;
  wire fch_issu1_inferred_i_170_n_0;
  wire fch_issu1_inferred_i_171_n_0;
  wire fch_issu1_inferred_i_172_n_0;
  wire fch_issu1_inferred_i_173_n_0;
  wire fch_issu1_inferred_i_174_n_0;
  wire fch_issu1_inferred_i_175_n_0;
  wire fch_issu1_inferred_i_176_n_0;
  wire fch_issu1_inferred_i_177_n_0;
  wire fch_issu1_inferred_i_178_n_0;
  wire fch_issu1_inferred_i_179_n_0;
  wire fch_issu1_inferred_i_17_n_0;
  wire fch_issu1_inferred_i_180_n_0;
  wire fch_issu1_inferred_i_181_n_0;
  wire fch_issu1_inferred_i_182_n_0;
  wire fch_issu1_inferred_i_183_n_0;
  wire fch_issu1_inferred_i_184_n_0;
  wire fch_issu1_inferred_i_185_n_0;
  wire fch_issu1_inferred_i_186_n_0;
  wire fch_issu1_inferred_i_187_n_0;
  wire fch_issu1_inferred_i_188_n_0;
  wire fch_issu1_inferred_i_189_n_0;
  wire fch_issu1_inferred_i_18_n_0;
  wire fch_issu1_inferred_i_190_n_0;
  wire fch_issu1_inferred_i_191_n_0;
  wire fch_issu1_inferred_i_192_n_0;
  wire fch_issu1_inferred_i_193_n_0;
  wire fch_issu1_inferred_i_194_n_0;
  wire fch_issu1_inferred_i_195_n_0;
  wire fch_issu1_inferred_i_196_n_0;
  wire fch_issu1_inferred_i_197_n_0;
  wire fch_issu1_inferred_i_198_n_0;
  wire fch_issu1_inferred_i_199_n_0;
  wire fch_issu1_inferred_i_19_n_0;
  wire fch_issu1_inferred_i_200_n_0;
  wire fch_issu1_inferred_i_201_n_0;
  wire fch_issu1_inferred_i_202_n_0;
  wire fch_issu1_inferred_i_203_n_0;
  wire fch_issu1_inferred_i_204_n_0;
  wire fch_issu1_inferred_i_20_n_0;
  wire fch_issu1_inferred_i_21_n_0;
  wire fch_issu1_inferred_i_22_n_0;
  wire fch_issu1_inferred_i_23_n_0;
  wire fch_issu1_inferred_i_24_n_0;
  wire fch_issu1_inferred_i_25_n_0;
  wire fch_issu1_inferred_i_26_n_0;
  wire fch_issu1_inferred_i_27_n_0;
  wire fch_issu1_inferred_i_28_n_0;
  wire fch_issu1_inferred_i_29_n_0;
  wire fch_issu1_inferred_i_2_n_0;
  wire fch_issu1_inferred_i_30_n_0;
  wire fch_issu1_inferred_i_31_n_0;
  wire fch_issu1_inferred_i_32_n_0;
  wire fch_issu1_inferred_i_33_n_0;
  wire fch_issu1_inferred_i_34_n_0;
  wire fch_issu1_inferred_i_35_n_0;
  wire fch_issu1_inferred_i_36_n_0;
  wire fch_issu1_inferred_i_37_n_0;
  wire fch_issu1_inferred_i_38_n_0;
  wire fch_issu1_inferred_i_39_n_0;
  wire fch_issu1_inferred_i_3_n_0;
  wire fch_issu1_inferred_i_40_n_0;
  wire fch_issu1_inferred_i_41_n_0;
  wire fch_issu1_inferred_i_42_n_0;
  wire fch_issu1_inferred_i_43_n_0;
  wire fch_issu1_inferred_i_44_n_0;
  wire fch_issu1_inferred_i_45_n_0;
  wire fch_issu1_inferred_i_46_n_0;
  wire fch_issu1_inferred_i_47_n_0;
  wire fch_issu1_inferred_i_48_n_0;
  wire fch_issu1_inferred_i_49_n_0;
  wire fch_issu1_inferred_i_4_n_0;
  wire fch_issu1_inferred_i_50_n_0;
  wire fch_issu1_inferred_i_51_n_0;
  wire fch_issu1_inferred_i_52_n_0;
  wire fch_issu1_inferred_i_53_n_0;
  wire fch_issu1_inferred_i_54_n_0;
  wire fch_issu1_inferred_i_55_n_0;
  wire fch_issu1_inferred_i_56_n_0;
  wire fch_issu1_inferred_i_57_n_0;
  wire fch_issu1_inferred_i_58_n_0;
  wire fch_issu1_inferred_i_59_n_0;
  wire fch_issu1_inferred_i_5_n_0;
  wire fch_issu1_inferred_i_60_n_0;
  wire fch_issu1_inferred_i_61_n_0;
  wire fch_issu1_inferred_i_62_n_0;
  wire fch_issu1_inferred_i_63_n_0;
  wire fch_issu1_inferred_i_64_n_0;
  wire fch_issu1_inferred_i_65_n_0;
  wire fch_issu1_inferred_i_66_n_0;
  wire fch_issu1_inferred_i_67_n_0;
  wire fch_issu1_inferred_i_68_n_0;
  wire fch_issu1_inferred_i_69_n_0;
  wire fch_issu1_inferred_i_6_n_0;
  wire fch_issu1_inferred_i_70_n_0;
  wire fch_issu1_inferred_i_71_n_0;
  wire fch_issu1_inferred_i_72_n_0;
  wire fch_issu1_inferred_i_73_n_0;
  wire fch_issu1_inferred_i_74_n_0;
  wire fch_issu1_inferred_i_75_n_0;
  wire fch_issu1_inferred_i_76_n_0;
  wire fch_issu1_inferred_i_77_n_0;
  wire fch_issu1_inferred_i_78_n_0;
  wire fch_issu1_inferred_i_79_n_0;
  wire fch_issu1_inferred_i_7_n_0;
  wire fch_issu1_inferred_i_80_n_0;
  wire fch_issu1_inferred_i_81_n_0;
  wire fch_issu1_inferred_i_82_n_0;
  wire fch_issu1_inferred_i_83_n_0;
  wire fch_issu1_inferred_i_84_n_0;
  wire fch_issu1_inferred_i_85_n_0;
  wire fch_issu1_inferred_i_86_n_0;
  wire fch_issu1_inferred_i_87_n_0;
  wire fch_issu1_inferred_i_88_n_0;
  wire fch_issu1_inferred_i_89_n_0;
  wire fch_issu1_inferred_i_8_n_0;
  wire fch_issu1_inferred_i_90_n_0;
  wire fch_issu1_inferred_i_91_n_0;
  wire fch_issu1_inferred_i_92_n_0;
  wire fch_issu1_inferred_i_93_n_0;
  wire fch_issu1_inferred_i_94_n_0;
  wire fch_issu1_inferred_i_95_n_0;
  wire fch_issu1_inferred_i_96_n_0;
  wire fch_issu1_inferred_i_97_n_0;
  wire fch_issu1_inferred_i_98_n_0;
  wire fch_issu1_inferred_i_99_n_0;
  wire fch_issu1_inferred_i_9_n_0;
  wire fch_leir_hir_i_2_n_0;
  wire fch_leir_nir_i_2_n_0;
  wire fch_memacc1;
  wire [15:0]fch_pc;
  wire [15:0]fch_pc0;
  wire [15:0]fch_pc1;
  (* DONT_TOUCH *) wire fch_term;
  wire fch_wrbufn0;
  wire fch_wrbufn1;
  wire [31:0]fdat;
  wire \grn[0]_i_1__0_n_0 ;
  wire \grn[0]_i_1__10_n_0 ;
  wire \grn[0]_i_1__11_n_0 ;
  wire \grn[0]_i_1__12_n_0 ;
  wire \grn[0]_i_1__13_n_0 ;
  wire \grn[0]_i_1__14_n_0 ;
  wire \grn[0]_i_1__15_n_0 ;
  wire \grn[0]_i_1__16_n_0 ;
  wire \grn[0]_i_1__17_n_0 ;
  wire \grn[0]_i_1__18_n_0 ;
  wire \grn[0]_i_1__19_n_0 ;
  wire \grn[0]_i_1__1_n_0 ;
  wire \grn[0]_i_1__20_n_0 ;
  wire \grn[0]_i_1__21_n_0 ;
  wire \grn[0]_i_1__22_n_0 ;
  wire \grn[0]_i_1__23_n_0 ;
  wire \grn[0]_i_1__24_n_0 ;
  wire \grn[0]_i_1__25_n_0 ;
  wire \grn[0]_i_1__26_n_0 ;
  wire \grn[0]_i_1__27_n_0 ;
  wire \grn[0]_i_1__28_n_0 ;
  wire \grn[0]_i_1__29_n_0 ;
  wire \grn[0]_i_1__2_n_0 ;
  wire \grn[0]_i_1__30_n_0 ;
  wire \grn[0]_i_1__3_n_0 ;
  wire \grn[0]_i_1__4_n_0 ;
  wire \grn[0]_i_1__5_n_0 ;
  wire \grn[0]_i_1__6_n_0 ;
  wire \grn[0]_i_1__7_n_0 ;
  wire \grn[0]_i_1__8_n_0 ;
  wire \grn[0]_i_1__9_n_0 ;
  wire \grn[10]_i_1__0_n_0 ;
  wire \grn[10]_i_1__10_n_0 ;
  wire \grn[10]_i_1__11_n_0 ;
  wire \grn[10]_i_1__12_n_0 ;
  wire \grn[10]_i_1__13_n_0 ;
  wire \grn[10]_i_1__14_n_0 ;
  wire \grn[10]_i_1__15_n_0 ;
  wire \grn[10]_i_1__16_n_0 ;
  wire \grn[10]_i_1__17_n_0 ;
  wire \grn[10]_i_1__18_n_0 ;
  wire \grn[10]_i_1__19_n_0 ;
  wire \grn[10]_i_1__1_n_0 ;
  wire \grn[10]_i_1__20_n_0 ;
  wire \grn[10]_i_1__21_n_0 ;
  wire \grn[10]_i_1__22_n_0 ;
  wire \grn[10]_i_1__23_n_0 ;
  wire \grn[10]_i_1__24_n_0 ;
  wire \grn[10]_i_1__25_n_0 ;
  wire \grn[10]_i_1__26_n_0 ;
  wire \grn[10]_i_1__27_n_0 ;
  wire \grn[10]_i_1__28_n_0 ;
  wire \grn[10]_i_1__29_n_0 ;
  wire \grn[10]_i_1__2_n_0 ;
  wire \grn[10]_i_1__30_n_0 ;
  wire \grn[10]_i_1__3_n_0 ;
  wire \grn[10]_i_1__4_n_0 ;
  wire \grn[10]_i_1__5_n_0 ;
  wire \grn[10]_i_1__6_n_0 ;
  wire \grn[10]_i_1__7_n_0 ;
  wire \grn[10]_i_1__8_n_0 ;
  wire \grn[10]_i_1__9_n_0 ;
  wire \grn[11]_i_1__0_n_0 ;
  wire \grn[11]_i_1__10_n_0 ;
  wire \grn[11]_i_1__11_n_0 ;
  wire \grn[11]_i_1__12_n_0 ;
  wire \grn[11]_i_1__13_n_0 ;
  wire \grn[11]_i_1__14_n_0 ;
  wire \grn[11]_i_1__15_n_0 ;
  wire \grn[11]_i_1__16_n_0 ;
  wire \grn[11]_i_1__17_n_0 ;
  wire \grn[11]_i_1__18_n_0 ;
  wire \grn[11]_i_1__19_n_0 ;
  wire \grn[11]_i_1__1_n_0 ;
  wire \grn[11]_i_1__20_n_0 ;
  wire \grn[11]_i_1__21_n_0 ;
  wire \grn[11]_i_1__22_n_0 ;
  wire \grn[11]_i_1__23_n_0 ;
  wire \grn[11]_i_1__24_n_0 ;
  wire \grn[11]_i_1__25_n_0 ;
  wire \grn[11]_i_1__26_n_0 ;
  wire \grn[11]_i_1__27_n_0 ;
  wire \grn[11]_i_1__28_n_0 ;
  wire \grn[11]_i_1__29_n_0 ;
  wire \grn[11]_i_1__2_n_0 ;
  wire \grn[11]_i_1__30_n_0 ;
  wire \grn[11]_i_1__3_n_0 ;
  wire \grn[11]_i_1__4_n_0 ;
  wire \grn[11]_i_1__5_n_0 ;
  wire \grn[11]_i_1__6_n_0 ;
  wire \grn[11]_i_1__7_n_0 ;
  wire \grn[11]_i_1__8_n_0 ;
  wire \grn[11]_i_1__9_n_0 ;
  wire \grn[12]_i_1__0_n_0 ;
  wire \grn[12]_i_1__10_n_0 ;
  wire \grn[12]_i_1__11_n_0 ;
  wire \grn[12]_i_1__12_n_0 ;
  wire \grn[12]_i_1__13_n_0 ;
  wire \grn[12]_i_1__14_n_0 ;
  wire \grn[12]_i_1__15_n_0 ;
  wire \grn[12]_i_1__16_n_0 ;
  wire \grn[12]_i_1__17_n_0 ;
  wire \grn[12]_i_1__18_n_0 ;
  wire \grn[12]_i_1__19_n_0 ;
  wire \grn[12]_i_1__1_n_0 ;
  wire \grn[12]_i_1__20_n_0 ;
  wire \grn[12]_i_1__21_n_0 ;
  wire \grn[12]_i_1__22_n_0 ;
  wire \grn[12]_i_1__23_n_0 ;
  wire \grn[12]_i_1__24_n_0 ;
  wire \grn[12]_i_1__25_n_0 ;
  wire \grn[12]_i_1__26_n_0 ;
  wire \grn[12]_i_1__27_n_0 ;
  wire \grn[12]_i_1__28_n_0 ;
  wire \grn[12]_i_1__29_n_0 ;
  wire \grn[12]_i_1__2_n_0 ;
  wire \grn[12]_i_1__30_n_0 ;
  wire \grn[12]_i_1__3_n_0 ;
  wire \grn[12]_i_1__4_n_0 ;
  wire \grn[12]_i_1__5_n_0 ;
  wire \grn[12]_i_1__6_n_0 ;
  wire \grn[12]_i_1__7_n_0 ;
  wire \grn[12]_i_1__8_n_0 ;
  wire \grn[12]_i_1__9_n_0 ;
  wire \grn[13]_i_1__0_n_0 ;
  wire \grn[13]_i_1__10_n_0 ;
  wire \grn[13]_i_1__11_n_0 ;
  wire \grn[13]_i_1__12_n_0 ;
  wire \grn[13]_i_1__13_n_0 ;
  wire \grn[13]_i_1__14_n_0 ;
  wire \grn[13]_i_1__15_n_0 ;
  wire \grn[13]_i_1__16_n_0 ;
  wire \grn[13]_i_1__17_n_0 ;
  wire \grn[13]_i_1__18_n_0 ;
  wire \grn[13]_i_1__19_n_0 ;
  wire \grn[13]_i_1__1_n_0 ;
  wire \grn[13]_i_1__20_n_0 ;
  wire \grn[13]_i_1__21_n_0 ;
  wire \grn[13]_i_1__22_n_0 ;
  wire \grn[13]_i_1__23_n_0 ;
  wire \grn[13]_i_1__24_n_0 ;
  wire \grn[13]_i_1__25_n_0 ;
  wire \grn[13]_i_1__26_n_0 ;
  wire \grn[13]_i_1__27_n_0 ;
  wire \grn[13]_i_1__28_n_0 ;
  wire \grn[13]_i_1__29_n_0 ;
  wire \grn[13]_i_1__2_n_0 ;
  wire \grn[13]_i_1__30_n_0 ;
  wire \grn[13]_i_1__3_n_0 ;
  wire \grn[13]_i_1__4_n_0 ;
  wire \grn[13]_i_1__5_n_0 ;
  wire \grn[13]_i_1__6_n_0 ;
  wire \grn[13]_i_1__7_n_0 ;
  wire \grn[13]_i_1__8_n_0 ;
  wire \grn[13]_i_1__9_n_0 ;
  wire \grn[14]_i_1__0_n_0 ;
  wire \grn[14]_i_1__10_n_0 ;
  wire \grn[14]_i_1__11_n_0 ;
  wire \grn[14]_i_1__12_n_0 ;
  wire \grn[14]_i_1__13_n_0 ;
  wire \grn[14]_i_1__14_n_0 ;
  wire \grn[14]_i_1__15_n_0 ;
  wire \grn[14]_i_1__16_n_0 ;
  wire \grn[14]_i_1__17_n_0 ;
  wire \grn[14]_i_1__18_n_0 ;
  wire \grn[14]_i_1__19_n_0 ;
  wire \grn[14]_i_1__1_n_0 ;
  wire \grn[14]_i_1__20_n_0 ;
  wire \grn[14]_i_1__21_n_0 ;
  wire \grn[14]_i_1__22_n_0 ;
  wire \grn[14]_i_1__23_n_0 ;
  wire \grn[14]_i_1__24_n_0 ;
  wire \grn[14]_i_1__25_n_0 ;
  wire \grn[14]_i_1__26_n_0 ;
  wire \grn[14]_i_1__27_n_0 ;
  wire \grn[14]_i_1__28_n_0 ;
  wire \grn[14]_i_1__29_n_0 ;
  wire \grn[14]_i_1__2_n_0 ;
  wire \grn[14]_i_1__30_n_0 ;
  wire \grn[14]_i_1__3_n_0 ;
  wire \grn[14]_i_1__4_n_0 ;
  wire \grn[14]_i_1__5_n_0 ;
  wire \grn[14]_i_1__6_n_0 ;
  wire \grn[14]_i_1__7_n_0 ;
  wire \grn[14]_i_1__8_n_0 ;
  wire \grn[14]_i_1__9_n_0 ;
  wire \grn[15]_i_1__0_n_0 ;
  wire \grn[15]_i_1__10_n_0 ;
  wire \grn[15]_i_1__11_n_0 ;
  wire \grn[15]_i_1__12_n_0 ;
  wire \grn[15]_i_1__13_n_0 ;
  wire \grn[15]_i_1__14_n_0 ;
  wire \grn[15]_i_1__15_n_0 ;
  wire \grn[15]_i_1__16_n_0 ;
  wire \grn[15]_i_1__17_n_0 ;
  wire \grn[15]_i_1__18_n_0 ;
  wire \grn[15]_i_1__19_n_0 ;
  wire \grn[15]_i_1__1_n_0 ;
  wire \grn[15]_i_1__20_n_0 ;
  wire \grn[15]_i_1__21_n_0 ;
  wire \grn[15]_i_1__22_n_0 ;
  wire \grn[15]_i_1__23_n_0 ;
  wire \grn[15]_i_1__24_n_0 ;
  wire \grn[15]_i_1__25_n_0 ;
  wire \grn[15]_i_1__26_n_0 ;
  wire \grn[15]_i_1__27_n_0 ;
  wire \grn[15]_i_1__28_n_0 ;
  wire \grn[15]_i_1__29_n_0 ;
  wire \grn[15]_i_1__2_n_0 ;
  wire \grn[15]_i_1__30_n_0 ;
  wire \grn[15]_i_1__3_n_0 ;
  wire \grn[15]_i_1__4_n_0 ;
  wire \grn[15]_i_1__5_n_0 ;
  wire \grn[15]_i_1__6_n_0 ;
  wire \grn[15]_i_1__7_n_0 ;
  wire \grn[15]_i_1__8_n_0 ;
  wire \grn[15]_i_1__9_n_0 ;
  wire \grn[15]_i_1_n_0 ;
  wire \grn[15]_i_2__0_n_0 ;
  wire \grn[15]_i_2__10_n_0 ;
  wire \grn[15]_i_2__11_n_0 ;
  wire \grn[15]_i_2__12_n_0 ;
  wire \grn[15]_i_2__13_n_0 ;
  wire \grn[15]_i_2__14_n_0 ;
  wire \grn[15]_i_2__15_n_0 ;
  wire \grn[15]_i_2__16_n_0 ;
  wire \grn[15]_i_2__17_n_0 ;
  wire \grn[15]_i_2__18_n_0 ;
  wire \grn[15]_i_2__19_n_0 ;
  wire \grn[15]_i_2__1_n_0 ;
  wire \grn[15]_i_2__20_n_0 ;
  wire \grn[15]_i_2__21_n_0 ;
  wire \grn[15]_i_2__22_n_0 ;
  wire \grn[15]_i_2__23_n_0 ;
  wire \grn[15]_i_2__24_n_0 ;
  wire \grn[15]_i_2__25_n_0 ;
  wire \grn[15]_i_2__26_n_0 ;
  wire \grn[15]_i_2__27_n_0 ;
  wire \grn[15]_i_2__28_n_0 ;
  wire \grn[15]_i_2__29_n_0 ;
  wire \grn[15]_i_2__2_n_0 ;
  wire \grn[15]_i_2__30_n_0 ;
  wire \grn[15]_i_2__3_n_0 ;
  wire \grn[15]_i_2__4_n_0 ;
  wire \grn[15]_i_2__5_n_0 ;
  wire \grn[15]_i_2__6_n_0 ;
  wire \grn[15]_i_2__7_n_0 ;
  wire \grn[15]_i_2__8_n_0 ;
  wire \grn[15]_i_2__9_n_0 ;
  wire \grn[15]_i_3__30_n_0 ;
  wire \grn[15]_i_3_n_0 ;
  wire \grn[15]_i_4__2_n_0 ;
  wire \grn[15]_i_4__6_n_0 ;
  wire \grn[15]_i_4__7_n_0 ;
  wire \grn[15]_i_5_n_0 ;
  wire \grn[15]_i_6__0_n_0 ;
  wire \grn[15]_i_6_n_0 ;
  wire \grn[15]_i_7__0_n_0 ;
  wire \grn[15]_i_7_n_0 ;
  wire \grn[1]_i_1__0_n_0 ;
  wire \grn[1]_i_1__10_n_0 ;
  wire \grn[1]_i_1__11_n_0 ;
  wire \grn[1]_i_1__12_n_0 ;
  wire \grn[1]_i_1__13_n_0 ;
  wire \grn[1]_i_1__14_n_0 ;
  wire \grn[1]_i_1__15_n_0 ;
  wire \grn[1]_i_1__16_n_0 ;
  wire \grn[1]_i_1__17_n_0 ;
  wire \grn[1]_i_1__18_n_0 ;
  wire \grn[1]_i_1__19_n_0 ;
  wire \grn[1]_i_1__1_n_0 ;
  wire \grn[1]_i_1__20_n_0 ;
  wire \grn[1]_i_1__21_n_0 ;
  wire \grn[1]_i_1__22_n_0 ;
  wire \grn[1]_i_1__23_n_0 ;
  wire \grn[1]_i_1__24_n_0 ;
  wire \grn[1]_i_1__25_n_0 ;
  wire \grn[1]_i_1__26_n_0 ;
  wire \grn[1]_i_1__27_n_0 ;
  wire \grn[1]_i_1__28_n_0 ;
  wire \grn[1]_i_1__29_n_0 ;
  wire \grn[1]_i_1__2_n_0 ;
  wire \grn[1]_i_1__30_n_0 ;
  wire \grn[1]_i_1__3_n_0 ;
  wire \grn[1]_i_1__4_n_0 ;
  wire \grn[1]_i_1__5_n_0 ;
  wire \grn[1]_i_1__6_n_0 ;
  wire \grn[1]_i_1__7_n_0 ;
  wire \grn[1]_i_1__8_n_0 ;
  wire \grn[1]_i_1__9_n_0 ;
  wire \grn[2]_i_1__0_n_0 ;
  wire \grn[2]_i_1__10_n_0 ;
  wire \grn[2]_i_1__11_n_0 ;
  wire \grn[2]_i_1__12_n_0 ;
  wire \grn[2]_i_1__13_n_0 ;
  wire \grn[2]_i_1__14_n_0 ;
  wire \grn[2]_i_1__15_n_0 ;
  wire \grn[2]_i_1__16_n_0 ;
  wire \grn[2]_i_1__17_n_0 ;
  wire \grn[2]_i_1__18_n_0 ;
  wire \grn[2]_i_1__19_n_0 ;
  wire \grn[2]_i_1__1_n_0 ;
  wire \grn[2]_i_1__20_n_0 ;
  wire \grn[2]_i_1__21_n_0 ;
  wire \grn[2]_i_1__22_n_0 ;
  wire \grn[2]_i_1__23_n_0 ;
  wire \grn[2]_i_1__24_n_0 ;
  wire \grn[2]_i_1__25_n_0 ;
  wire \grn[2]_i_1__26_n_0 ;
  wire \grn[2]_i_1__27_n_0 ;
  wire \grn[2]_i_1__28_n_0 ;
  wire \grn[2]_i_1__29_n_0 ;
  wire \grn[2]_i_1__2_n_0 ;
  wire \grn[2]_i_1__30_n_0 ;
  wire \grn[2]_i_1__3_n_0 ;
  wire \grn[2]_i_1__4_n_0 ;
  wire \grn[2]_i_1__5_n_0 ;
  wire \grn[2]_i_1__6_n_0 ;
  wire \grn[2]_i_1__7_n_0 ;
  wire \grn[2]_i_1__8_n_0 ;
  wire \grn[2]_i_1__9_n_0 ;
  wire \grn[3]_i_1__0_n_0 ;
  wire \grn[3]_i_1__10_n_0 ;
  wire \grn[3]_i_1__11_n_0 ;
  wire \grn[3]_i_1__12_n_0 ;
  wire \grn[3]_i_1__13_n_0 ;
  wire \grn[3]_i_1__14_n_0 ;
  wire \grn[3]_i_1__15_n_0 ;
  wire \grn[3]_i_1__16_n_0 ;
  wire \grn[3]_i_1__17_n_0 ;
  wire \grn[3]_i_1__18_n_0 ;
  wire \grn[3]_i_1__19_n_0 ;
  wire \grn[3]_i_1__1_n_0 ;
  wire \grn[3]_i_1__20_n_0 ;
  wire \grn[3]_i_1__21_n_0 ;
  wire \grn[3]_i_1__22_n_0 ;
  wire \grn[3]_i_1__23_n_0 ;
  wire \grn[3]_i_1__24_n_0 ;
  wire \grn[3]_i_1__25_n_0 ;
  wire \grn[3]_i_1__26_n_0 ;
  wire \grn[3]_i_1__27_n_0 ;
  wire \grn[3]_i_1__28_n_0 ;
  wire \grn[3]_i_1__29_n_0 ;
  wire \grn[3]_i_1__2_n_0 ;
  wire \grn[3]_i_1__30_n_0 ;
  wire \grn[3]_i_1__3_n_0 ;
  wire \grn[3]_i_1__4_n_0 ;
  wire \grn[3]_i_1__5_n_0 ;
  wire \grn[3]_i_1__6_n_0 ;
  wire \grn[3]_i_1__7_n_0 ;
  wire \grn[3]_i_1__8_n_0 ;
  wire \grn[3]_i_1__9_n_0 ;
  wire \grn[4]_i_1__0_n_0 ;
  wire \grn[4]_i_1__10_n_0 ;
  wire \grn[4]_i_1__11_n_0 ;
  wire \grn[4]_i_1__12_n_0 ;
  wire \grn[4]_i_1__13_n_0 ;
  wire \grn[4]_i_1__14_n_0 ;
  wire \grn[4]_i_1__15_n_0 ;
  wire \grn[4]_i_1__16_n_0 ;
  wire \grn[4]_i_1__17_n_0 ;
  wire \grn[4]_i_1__18_n_0 ;
  wire \grn[4]_i_1__19_n_0 ;
  wire \grn[4]_i_1__1_n_0 ;
  wire \grn[4]_i_1__20_n_0 ;
  wire \grn[4]_i_1__21_n_0 ;
  wire \grn[4]_i_1__22_n_0 ;
  wire \grn[4]_i_1__23_n_0 ;
  wire \grn[4]_i_1__24_n_0 ;
  wire \grn[4]_i_1__25_n_0 ;
  wire \grn[4]_i_1__26_n_0 ;
  wire \grn[4]_i_1__27_n_0 ;
  wire \grn[4]_i_1__28_n_0 ;
  wire \grn[4]_i_1__29_n_0 ;
  wire \grn[4]_i_1__2_n_0 ;
  wire \grn[4]_i_1__30_n_0 ;
  wire \grn[4]_i_1__3_n_0 ;
  wire \grn[4]_i_1__4_n_0 ;
  wire \grn[4]_i_1__5_n_0 ;
  wire \grn[4]_i_1__6_n_0 ;
  wire \grn[4]_i_1__7_n_0 ;
  wire \grn[4]_i_1__8_n_0 ;
  wire \grn[4]_i_1__9_n_0 ;
  wire \grn[5]_i_1__0_n_0 ;
  wire \grn[5]_i_1__10_n_0 ;
  wire \grn[5]_i_1__11_n_0 ;
  wire \grn[5]_i_1__12_n_0 ;
  wire \grn[5]_i_1__13_n_0 ;
  wire \grn[5]_i_1__14_n_0 ;
  wire \grn[5]_i_1__15_n_0 ;
  wire \grn[5]_i_1__16_n_0 ;
  wire \grn[5]_i_1__17_n_0 ;
  wire \grn[5]_i_1__18_n_0 ;
  wire \grn[5]_i_1__19_n_0 ;
  wire \grn[5]_i_1__1_n_0 ;
  wire \grn[5]_i_1__20_n_0 ;
  wire \grn[5]_i_1__21_n_0 ;
  wire \grn[5]_i_1__22_n_0 ;
  wire \grn[5]_i_1__23_n_0 ;
  wire \grn[5]_i_1__24_n_0 ;
  wire \grn[5]_i_1__25_n_0 ;
  wire \grn[5]_i_1__26_n_0 ;
  wire \grn[5]_i_1__27_n_0 ;
  wire \grn[5]_i_1__28_n_0 ;
  wire \grn[5]_i_1__29_n_0 ;
  wire \grn[5]_i_1__2_n_0 ;
  wire \grn[5]_i_1__30_n_0 ;
  wire \grn[5]_i_1__3_n_0 ;
  wire \grn[5]_i_1__4_n_0 ;
  wire \grn[5]_i_1__5_n_0 ;
  wire \grn[5]_i_1__6_n_0 ;
  wire \grn[5]_i_1__7_n_0 ;
  wire \grn[5]_i_1__8_n_0 ;
  wire \grn[5]_i_1__9_n_0 ;
  wire \grn[6]_i_1__0_n_0 ;
  wire \grn[6]_i_1__10_n_0 ;
  wire \grn[6]_i_1__11_n_0 ;
  wire \grn[6]_i_1__12_n_0 ;
  wire \grn[6]_i_1__13_n_0 ;
  wire \grn[6]_i_1__14_n_0 ;
  wire \grn[6]_i_1__15_n_0 ;
  wire \grn[6]_i_1__16_n_0 ;
  wire \grn[6]_i_1__17_n_0 ;
  wire \grn[6]_i_1__18_n_0 ;
  wire \grn[6]_i_1__19_n_0 ;
  wire \grn[6]_i_1__1_n_0 ;
  wire \grn[6]_i_1__20_n_0 ;
  wire \grn[6]_i_1__21_n_0 ;
  wire \grn[6]_i_1__22_n_0 ;
  wire \grn[6]_i_1__23_n_0 ;
  wire \grn[6]_i_1__24_n_0 ;
  wire \grn[6]_i_1__25_n_0 ;
  wire \grn[6]_i_1__26_n_0 ;
  wire \grn[6]_i_1__27_n_0 ;
  wire \grn[6]_i_1__28_n_0 ;
  wire \grn[6]_i_1__29_n_0 ;
  wire \grn[6]_i_1__2_n_0 ;
  wire \grn[6]_i_1__30_n_0 ;
  wire \grn[6]_i_1__3_n_0 ;
  wire \grn[6]_i_1__4_n_0 ;
  wire \grn[6]_i_1__5_n_0 ;
  wire \grn[6]_i_1__6_n_0 ;
  wire \grn[6]_i_1__7_n_0 ;
  wire \grn[6]_i_1__8_n_0 ;
  wire \grn[6]_i_1__9_n_0 ;
  wire \grn[7]_i_1__0_n_0 ;
  wire \grn[7]_i_1__10_n_0 ;
  wire \grn[7]_i_1__11_n_0 ;
  wire \grn[7]_i_1__12_n_0 ;
  wire \grn[7]_i_1__13_n_0 ;
  wire \grn[7]_i_1__14_n_0 ;
  wire \grn[7]_i_1__15_n_0 ;
  wire \grn[7]_i_1__16_n_0 ;
  wire \grn[7]_i_1__17_n_0 ;
  wire \grn[7]_i_1__18_n_0 ;
  wire \grn[7]_i_1__19_n_0 ;
  wire \grn[7]_i_1__1_n_0 ;
  wire \grn[7]_i_1__20_n_0 ;
  wire \grn[7]_i_1__21_n_0 ;
  wire \grn[7]_i_1__22_n_0 ;
  wire \grn[7]_i_1__23_n_0 ;
  wire \grn[7]_i_1__24_n_0 ;
  wire \grn[7]_i_1__25_n_0 ;
  wire \grn[7]_i_1__26_n_0 ;
  wire \grn[7]_i_1__27_n_0 ;
  wire \grn[7]_i_1__28_n_0 ;
  wire \grn[7]_i_1__29_n_0 ;
  wire \grn[7]_i_1__2_n_0 ;
  wire \grn[7]_i_1__30_n_0 ;
  wire \grn[7]_i_1__3_n_0 ;
  wire \grn[7]_i_1__4_n_0 ;
  wire \grn[7]_i_1__5_n_0 ;
  wire \grn[7]_i_1__6_n_0 ;
  wire \grn[7]_i_1__7_n_0 ;
  wire \grn[7]_i_1__8_n_0 ;
  wire \grn[7]_i_1__9_n_0 ;
  wire \grn[8]_i_1__0_n_0 ;
  wire \grn[8]_i_1__10_n_0 ;
  wire \grn[8]_i_1__11_n_0 ;
  wire \grn[8]_i_1__12_n_0 ;
  wire \grn[8]_i_1__13_n_0 ;
  wire \grn[8]_i_1__14_n_0 ;
  wire \grn[8]_i_1__15_n_0 ;
  wire \grn[8]_i_1__16_n_0 ;
  wire \grn[8]_i_1__17_n_0 ;
  wire \grn[8]_i_1__18_n_0 ;
  wire \grn[8]_i_1__19_n_0 ;
  wire \grn[8]_i_1__1_n_0 ;
  wire \grn[8]_i_1__20_n_0 ;
  wire \grn[8]_i_1__21_n_0 ;
  wire \grn[8]_i_1__22_n_0 ;
  wire \grn[8]_i_1__23_n_0 ;
  wire \grn[8]_i_1__24_n_0 ;
  wire \grn[8]_i_1__25_n_0 ;
  wire \grn[8]_i_1__26_n_0 ;
  wire \grn[8]_i_1__27_n_0 ;
  wire \grn[8]_i_1__28_n_0 ;
  wire \grn[8]_i_1__29_n_0 ;
  wire \grn[8]_i_1__2_n_0 ;
  wire \grn[8]_i_1__30_n_0 ;
  wire \grn[8]_i_1__3_n_0 ;
  wire \grn[8]_i_1__4_n_0 ;
  wire \grn[8]_i_1__5_n_0 ;
  wire \grn[8]_i_1__6_n_0 ;
  wire \grn[8]_i_1__7_n_0 ;
  wire \grn[8]_i_1__8_n_0 ;
  wire \grn[8]_i_1__9_n_0 ;
  wire \grn[9]_i_1__0_n_0 ;
  wire \grn[9]_i_1__10_n_0 ;
  wire \grn[9]_i_1__11_n_0 ;
  wire \grn[9]_i_1__12_n_0 ;
  wire \grn[9]_i_1__13_n_0 ;
  wire \grn[9]_i_1__14_n_0 ;
  wire \grn[9]_i_1__15_n_0 ;
  wire \grn[9]_i_1__16_n_0 ;
  wire \grn[9]_i_1__17_n_0 ;
  wire \grn[9]_i_1__18_n_0 ;
  wire \grn[9]_i_1__19_n_0 ;
  wire \grn[9]_i_1__1_n_0 ;
  wire \grn[9]_i_1__20_n_0 ;
  wire \grn[9]_i_1__21_n_0 ;
  wire \grn[9]_i_1__22_n_0 ;
  wire \grn[9]_i_1__23_n_0 ;
  wire \grn[9]_i_1__24_n_0 ;
  wire \grn[9]_i_1__25_n_0 ;
  wire \grn[9]_i_1__26_n_0 ;
  wire \grn[9]_i_1__27_n_0 ;
  wire \grn[9]_i_1__28_n_0 ;
  wire \grn[9]_i_1__29_n_0 ;
  wire \grn[9]_i_1__2_n_0 ;
  wire \grn[9]_i_1__30_n_0 ;
  wire \grn[9]_i_1__3_n_0 ;
  wire \grn[9]_i_1__4_n_0 ;
  wire \grn[9]_i_1__5_n_0 ;
  wire \grn[9]_i_1__6_n_0 ;
  wire \grn[9]_i_1__7_n_0 ;
  wire \grn[9]_i_1__8_n_0 ;
  wire \grn[9]_i_1__9_n_0 ;
  wire \ir0_id_fl[20]_i_1_n_0 ;
  wire \ir0_id_fl[20]_i_2_n_0 ;
  wire \ir0_id_fl[20]_i_3_n_0 ;
  wire \ir0_id_fl[20]_i_4_n_0 ;
  wire \ir0_id_fl[20]_i_5_n_0 ;
  wire \ir0_id_fl[20]_i_6_n_0 ;
  wire \ir0_id_fl[20]_i_7_n_0 ;
  wire \ir0_id_fl[20]_i_8_n_0 ;
  wire \ir0_id_fl[21]_i_10_n_0 ;
  wire \ir0_id_fl[21]_i_11_n_0 ;
  wire \ir0_id_fl[21]_i_1_n_0 ;
  wire \ir0_id_fl[21]_i_2_n_0 ;
  wire \ir0_id_fl[21]_i_3_n_0 ;
  wire \ir0_id_fl[21]_i_4_n_0 ;
  wire \ir0_id_fl[21]_i_5_n_0 ;
  wire \ir0_id_fl[21]_i_6_n_0 ;
  wire \ir0_id_fl[21]_i_7_n_0 ;
  wire \ir0_id_fl[21]_i_8_n_0 ;
  wire \ir0_id_fl[21]_i_9_n_0 ;
  wire ir0_inferred_i_17_n_0;
  wire ir0_inferred_i_18_n_0;
  wire ir0_inferred_i_19_n_0;
  wire ir0_inferred_i_20_n_0;
  wire ir0_inferred_i_21_n_0;
  wire ir0_inferred_i_22_n_0;
  wire ir0_inferred_i_23_n_0;
  wire ir0_inferred_i_24_n_0;
  wire ir0_inferred_i_25_n_0;
  wire ir0_inferred_i_26_n_0;
  wire ir0_inferred_i_27_n_0;
  wire ir0_inferred_i_28_n_0;
  wire ir0_inferred_i_29_n_0;
  wire ir0_inferred_i_30_n_0;
  wire ir0_inferred_i_31_n_0;
  wire ir0_inferred_i_32_n_0;
  wire \ir1_id_fl[20]_i_2_n_0 ;
  wire \ir1_id_fl[21]_i_2_n_0 ;
  wire ir1_inferred_i_17_n_0;
  wire ir1_inferred_i_18_n_0;
  wire ir1_inferred_i_19_n_0;
  wire ir1_inferred_i_20_n_0;
  wire ir1_inferred_i_21_n_0;
  wire ir1_inferred_i_22_n_0;
  wire ir1_inferred_i_23_n_0;
  wire ir1_inferred_i_24_n_0;
  wire ir1_inferred_i_25_n_0;
  wire ir1_inferred_i_26_n_0;
  wire ir1_inferred_i_27_n_0;
  wire ir1_inferred_i_28_n_0;
  wire ir1_inferred_i_29_n_0;
  wire ir1_inferred_i_30_n_0;
  wire ir1_inferred_i_31_n_0;
  wire ir1_inferred_i_32_n_0;
  wire ir1_inferred_i_33_n_0;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire \iv[15]_i_4_n_0 ;
  wire [5:4]\mem/bctl/ctl/p_0_in ;
  wire [1:1]\mem/bctl/ctl/stat_nx ;
  wire \mem/bctl/fch_term_fl ;
  wire \mem/mem_accslot ;
  wire [3:0]\mem/read_cyc ;
  wire \mul_a[15]_i_1__0_n_0 ;
  wire \mul_a[15]_i_1_n_0 ;
  wire \mul_a[16]_i_1__0_n_0 ;
  wire \mul_a[16]_i_1_n_0 ;
  wire \mul_a[31]_i_1__0_n_0 ;
  wire \mul_a[31]_i_1_n_0 ;
  wire \mul_a[32]_i_1__0_n_0 ;
  wire \mul_a[32]_i_1_n_0 ;
  wire \mul_b[31]_i_1__0_n_0 ;
  wire \mul_b[31]_i_1_n_0 ;
  wire \mul_b[32]_i_1__0_n_0 ;
  wire \mul_b[32]_i_1_n_0 ;
  wire \mulh[15]_i_1__0_n_0 ;
  wire \mulh[15]_i_1_n_0 ;
  wire \nir_id[12]_i_2_n_0 ;
  wire \nir_id[12]_i_3_n_0 ;
  wire \nir_id[12]_i_4_n_0 ;
  wire \nir_id[13]_i_2_n_0 ;
  wire \nir_id[13]_i_3_n_0 ;
  wire \nir_id[13]_i_4_n_0 ;
  wire \nir_id[13]_i_5_n_0 ;
  wire \nir_id[13]_i_6_n_0 ;
  wire \nir_id[13]_i_7_n_0 ;
  wire \nir_id[13]_i_8_n_0 ;
  wire \nir_id[13]_i_9_n_0 ;
  wire \nir_id[14]_i_10_n_0 ;
  wire \nir_id[14]_i_11_n_0 ;
  wire \nir_id[14]_i_12_n_0 ;
  wire \nir_id[14]_i_2_n_0 ;
  wire \nir_id[14]_i_3_n_0 ;
  wire \nir_id[14]_i_4_n_0 ;
  wire \nir_id[14]_i_5_n_0 ;
  wire \nir_id[14]_i_6_n_0 ;
  wire \nir_id[14]_i_7_n_0 ;
  wire \nir_id[14]_i_8_n_0 ;
  wire \nir_id[14]_i_9_n_0 ;
  wire \nir_id[15]_i_2_n_0 ;
  wire \nir_id[16]_i_2_n_0 ;
  wire \nir_id[16]_i_3_n_0 ;
  wire \nir_id[16]_i_4_n_0 ;
  wire \nir_id[16]_i_5_n_0 ;
  wire \nir_id[16]_i_6_n_0 ;
  wire \nir_id[17]_i_2_n_0 ;
  wire \nir_id[17]_i_3_n_0 ;
  wire \nir_id[17]_i_4_n_0 ;
  wire \nir_id[17]_i_5_n_0 ;
  wire \nir_id[17]_i_6_n_0 ;
  wire \nir_id[17]_i_7_n_0 ;
  wire \nir_id[18]_i_2_n_0 ;
  wire \nir_id[18]_i_3_n_0 ;
  wire \nir_id[18]_i_4_n_0 ;
  wire \nir_id[18]_i_5_n_0 ;
  wire \nir_id[18]_i_6_n_0 ;
  wire \nir_id[18]_i_7_n_0 ;
  wire \nir_id[19]_i_2_n_0 ;
  wire \nir_id[19]_i_3_n_0 ;
  wire \nir_id[19]_i_4_n_0 ;
  wire \nir_id[19]_i_5_n_0 ;
  wire \nir_id[19]_i_6_n_0 ;
  wire \nir_id[19]_i_7_n_0 ;
  wire \nir_id[20]_i_1_n_0 ;
  wire \nir_id[20]_i_2_n_0 ;
  wire \nir_id[20]_i_3_n_0 ;
  wire \nir_id[20]_i_4_n_0 ;
  wire \nir_id[20]_i_5_n_0 ;
  wire \nir_id[20]_i_6_n_0 ;
  wire \nir_id[20]_i_7_n_0 ;
  wire \nir_id[20]_i_8_n_0 ;
  wire \nir_id[21]_i_10_n_0 ;
  wire \nir_id[21]_i_2_n_0 ;
  wire \nir_id[21]_i_3_n_0 ;
  wire \nir_id[21]_i_4_n_0 ;
  wire \nir_id[21]_i_5_n_0 ;
  wire \nir_id[21]_i_6_n_0 ;
  wire \nir_id[21]_i_7_n_0 ;
  wire \nir_id[21]_i_8_n_0 ;
  wire \nir_id[21]_i_9_n_0 ;
  wire \nir_id[24]_i_11_n_0 ;
  wire \nir_id[24]_i_12_n_0 ;
  wire \nir_id[24]_i_13_n_0 ;
  wire \nir_id[24]_i_14_n_0 ;
  wire \nir_id[24]_i_15_n_0 ;
  wire \nir_id[24]_i_16_n_0 ;
  wire \nir_id[24]_i_17_n_0 ;
  wire \nir_id[24]_i_18_n_0 ;
  wire \nir_id[24]_i_19_n_0 ;
  wire \nir_id[24]_i_20_n_0 ;
  wire \nir_id[24]_i_21_n_0 ;
  wire \nir_id[24]_i_22_n_0 ;
  wire \nir_id[24]_i_23_n_0 ;
  wire \nir_id[24]_i_24_n_0 ;
  wire \nir_id[24]_i_25_n_0 ;
  wire \nir_id[24]_i_3_n_0 ;
  wire \nir_id[24]_i_4_n_0 ;
  wire \nir_id[24]_i_5_n_0 ;
  wire \nir_id[24]_i_6_n_0 ;
  wire \nir_id[24]_i_7_n_0 ;
  wire \nir_id[24]_i_8_n_0 ;
  wire [32:0]niss_dsp_a0;
  wire \niss_dsp_a0[15]_INST_0_i_1_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_10_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_11_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_12_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_13_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_14_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_15_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_16_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_1_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_2_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_3_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_4_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_5_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_6_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_7_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_8_n_0 ;
  wire \niss_dsp_a0[32]_INST_0_i_9_n_0 ;
  wire [32:0]niss_dsp_a1;
  wire \niss_dsp_a1[15]_INST_0_i_10_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_11_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_12_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_13_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_14_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_15_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_16_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_17_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_18_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_19_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_1_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_20_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_21_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_22_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_23_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_24_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_25_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_26_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_27_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_28_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_29_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_30_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_31_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_3_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_4_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_5_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_6_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_7_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_8_n_0 ;
  wire \niss_dsp_a1[15]_INST_0_i_9_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_10_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_11_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_12_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_13_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_14_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_15_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_16_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_17_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_18_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_19_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_1_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_20_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_21_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_22_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_23_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_24_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_25_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_26_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_27_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_28_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_29_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_2_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_30_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_31_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_32_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_33_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_34_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_35_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_36_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_37_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_38_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_39_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_3_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_40_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_41_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_42_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_43_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_44_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_45_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_46_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_47_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_48_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_49_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_4_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_5_n_0 ;
  wire \niss_dsp_a1[32]_INST_0_i_9_n_0 ;
  wire [32:0]niss_dsp_b0;
  wire \niss_dsp_b0[4]_INST_0_i_1_n_0 ;
  wire [32:0]niss_dsp_b1;
  wire \niss_dsp_b1[0]_INST_0_i_12_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_13_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_1_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_23_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_24_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_25_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_26_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_27_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_28_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_29_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_2_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_30_n_0 ;
  wire \niss_dsp_b1[0]_INST_0_i_8_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_12_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_13_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_1_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_23_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_24_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_25_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_26_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_27_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_28_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_29_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_2_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_30_n_0 ;
  wire \niss_dsp_b1[1]_INST_0_i_8_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_13_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_14_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_1_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_27_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_28_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_29_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_2_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_30_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_31_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_32_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_33_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_34_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_35_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_36_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_37_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_38_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_39_n_0 ;
  wire \niss_dsp_b1[2]_INST_0_i_8_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_1_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_20_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_21_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_22_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_23_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_24_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_25_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_26_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_27_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_28_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_29_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_2_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_30_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_31_n_0 ;
  wire \niss_dsp_b1[3]_INST_0_i_3_n_0 ;
  wire \niss_dsp_b1[4]_INST_0_i_1_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_1_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_25_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_26_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_28_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_2_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_30_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_31_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_33_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_35_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_37_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_38_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_3_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_40_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_42_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_45_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_46_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_48_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_49_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_50_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_51_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_52_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_53_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_54_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_55_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_56_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_57_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_58_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_59_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_60_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_61_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_62_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_63_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_64_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_65_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_66_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_67_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_68_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_69_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_70_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_71_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_72_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_73_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_74_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_75_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_76_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_77_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_78_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_79_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_80_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_81_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_82_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_83_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_84_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_85_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_86_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_87_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_88_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_89_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_8_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_90_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_91_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_92_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_93_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_94_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_95_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_96_n_0 ;
  wire \niss_dsp_b1[5]_INST_0_i_9_n_0 ;
  wire \niss_dsp_b1[6]_INST_0_i_1_n_0 ;
  wire \niss_dsp_b1[6]_INST_0_i_2_n_0 ;
  wire \niss_dsp_b1[6]_INST_0_i_5_n_0 ;
  wire \niss_dsp_b1[7]_INST_0_i_2_n_0 ;
  wire \niss_dsp_b1[7]_INST_0_i_5_n_0 ;
  wire [65:0]niss_dsp_c0;
  wire [65:0]niss_dsp_c1;
  wire [29:19]p_2_in;
  wire [15:0]p_2_in1_in;
  wire [15:0]p_2_in4_in;
  wire \pc0[10]_i_2_n_0 ;
  wire \pc0[10]_i_3_n_0 ;
  wire \pc0[11]_i_2_n_0 ;
  wire \pc0[11]_i_4_n_0 ;
  wire \pc0[12]_i_2_n_0 ;
  wire \pc0[12]_i_3_n_0 ;
  wire \pc0[13]_i_2_n_0 ;
  wire \pc0[13]_i_3_n_0 ;
  wire \pc0[14]_i_2_n_0 ;
  wire \pc0[14]_i_3_n_0 ;
  wire \pc0[15]_i_2_n_0 ;
  wire \pc0[15]_i_4_n_0 ;
  wire \pc0[15]_i_5_n_0 ;
  wire \pc0[15]_i_6_n_0 ;
  wire \pc0[15]_i_7_n_0 ;
  wire \pc0[15]_i_8_n_0 ;
  wire \pc0[1]_i_2_n_0 ;
  wire \pc0[1]_i_3_n_0 ;
  wire \pc0[2]_i_2_n_0 ;
  wire \pc0[2]_i_3_n_0 ;
  wire \pc0[3]_i_2_n_0 ;
  wire \pc0[3]_i_4_n_0 ;
  wire \pc0[3]_i_5_n_0 ;
  wire \pc0[3]_i_6_n_0 ;
  wire \pc0[4]_i_2_n_0 ;
  wire \pc0[4]_i_3_n_0 ;
  wire \pc0[5]_i_2_n_0 ;
  wire \pc0[5]_i_3_n_0 ;
  wire \pc0[6]_i_2_n_0 ;
  wire \pc0[6]_i_3_n_0 ;
  wire \pc0[7]_i_2_n_0 ;
  wire \pc0[7]_i_4_n_0 ;
  wire \pc0[8]_i_2_n_0 ;
  wire \pc0[8]_i_3_n_0 ;
  wire \pc0[9]_i_2_n_0 ;
  wire \pc0[9]_i_3_n_0 ;
  wire \pc0_reg[11]_i_3_n_0 ;
  wire \pc0_reg[11]_i_3_n_1 ;
  wire \pc0_reg[11]_i_3_n_2 ;
  wire \pc0_reg[11]_i_3_n_3 ;
  wire \pc0_reg[15]_i_3_n_1 ;
  wire \pc0_reg[15]_i_3_n_2 ;
  wire \pc0_reg[15]_i_3_n_3 ;
  wire \pc0_reg[3]_i_3_n_0 ;
  wire \pc0_reg[3]_i_3_n_1 ;
  wire \pc0_reg[3]_i_3_n_2 ;
  wire \pc0_reg[3]_i_3_n_3 ;
  wire \pc0_reg[7]_i_3_n_0 ;
  wire \pc0_reg[7]_i_3_n_1 ;
  wire \pc0_reg[7]_i_3_n_2 ;
  wire \pc0_reg[7]_i_3_n_3 ;
  wire \pc1[11]_i_2_n_0 ;
  wire \pc1[11]_i_3_n_0 ;
  wire \pc1[11]_i_4_n_0 ;
  wire \pc1[11]_i_5_n_0 ;
  wire \pc1[15]_i_2_n_0 ;
  wire \pc1[15]_i_3_n_0 ;
  wire \pc1[15]_i_4_n_0 ;
  wire \pc1[15]_i_5_n_0 ;
  wire \pc1[3]_i_2_n_0 ;
  wire \pc1[3]_i_3_n_0 ;
  wire \pc1[3]_i_4_n_0 ;
  wire \pc1[3]_i_5_n_0 ;
  wire \pc1[3]_i_6_n_0 ;
  wire \pc1[3]_i_7_n_0 ;
  wire \pc1[3]_i_8_n_0 ;
  wire \pc1[7]_i_2_n_0 ;
  wire \pc1[7]_i_3_n_0 ;
  wire \pc1[7]_i_4_n_0 ;
  wire \pc1[7]_i_5_n_0 ;
  wire \pc1_reg[11]_i_1_n_0 ;
  wire \pc1_reg[11]_i_1_n_1 ;
  wire \pc1_reg[11]_i_1_n_2 ;
  wire \pc1_reg[11]_i_1_n_3 ;
  wire \pc1_reg[11]_i_1_n_4 ;
  wire \pc1_reg[11]_i_1_n_5 ;
  wire \pc1_reg[11]_i_1_n_6 ;
  wire \pc1_reg[11]_i_1_n_7 ;
  wire \pc1_reg[15]_i_1_n_1 ;
  wire \pc1_reg[15]_i_1_n_2 ;
  wire \pc1_reg[15]_i_1_n_3 ;
  wire \pc1_reg[15]_i_1_n_4 ;
  wire \pc1_reg[15]_i_1_n_5 ;
  wire \pc1_reg[15]_i_1_n_6 ;
  wire \pc1_reg[15]_i_1_n_7 ;
  wire \pc1_reg[3]_i_1_n_0 ;
  wire \pc1_reg[3]_i_1_n_1 ;
  wire \pc1_reg[3]_i_1_n_2 ;
  wire \pc1_reg[3]_i_1_n_3 ;
  wire \pc1_reg[3]_i_1_n_4 ;
  wire \pc1_reg[3]_i_1_n_5 ;
  wire \pc1_reg[3]_i_1_n_6 ;
  wire \pc1_reg[3]_i_1_n_7 ;
  wire \pc1_reg[7]_i_1_n_0 ;
  wire \pc1_reg[7]_i_1_n_1 ;
  wire \pc1_reg[7]_i_1_n_2 ;
  wire \pc1_reg[7]_i_1_n_3 ;
  wire \pc1_reg[7]_i_1_n_4 ;
  wire \pc1_reg[7]_i_1_n_5 ;
  wire \pc1_reg[7]_i_1_n_6 ;
  wire \pc1_reg[7]_i_1_n_7 ;
  wire \pc[0]_i_3_n_0 ;
  wire \pc[10]_i_3_n_0 ;
  wire \pc[11]_i_3_n_0 ;
  wire \pc[12]_i_4_n_0 ;
  wire \pc[13]_i_4_n_0 ;
  wire \pc[14]_i_4_n_0 ;
  wire \pc[15]_i_11_n_0 ;
  wire \pc[15]_i_12_n_0 ;
  wire \pc[15]_i_7_n_0 ;
  wire \pc[1]_i_3_n_0 ;
  wire \pc[2]_i_4_n_0 ;
  wire \pc[3]_i_4_n_0 ;
  wire \pc[4]_i_10_n_0 ;
  wire \pc[4]_i_11_n_0 ;
  wire \pc[4]_i_12_n_0 ;
  wire \pc[4]_i_13_n_0 ;
  wire \pc[4]_i_4_n_0 ;
  wire \pc[4]_i_5_n_0 ;
  wire \pc[4]_i_6_n_0 ;
  wire \pc[4]_i_7_n_0 ;
  wire \pc[4]_i_8_n_0 ;
  wire \pc[4]_i_9_n_0 ;
  wire \pc[5]_i_10_n_0 ;
  wire \pc[5]_i_11_n_0 ;
  wire \pc[5]_i_12_n_0 ;
  wire \pc[5]_i_13_n_0 ;
  wire \pc[5]_i_14_n_0 ;
  wire \pc[5]_i_15_n_0 ;
  wire \pc[5]_i_4_n_0 ;
  wire \pc[5]_i_5_n_0 ;
  wire \pc[5]_i_6_n_0 ;
  wire \pc[5]_i_7_n_0 ;
  wire \pc[5]_i_8_n_0 ;
  wire \pc[5]_i_9_n_0 ;
  wire \pc[6]_i_3_n_0 ;
  wire \pc[7]_i_4_n_0 ;
  wire \pc[8]_i_3_n_0 ;
  wire \pc[9]_i_3_n_0 ;
  wire \quo[31]_i_1__0_n_0 ;
  wire \quo[31]_i_1_n_0 ;
  wire \quo[31]_i_3__0_n_0 ;
  wire \quo[31]_i_3_n_0 ;
  wire \quo[31]_i_4__0_n_0 ;
  wire \quo[31]_i_4_n_0 ;
  wire \quo[31]_i_5__0_n_0 ;
  wire \quo[31]_i_5_n_0 ;
  wire rem0_carry__0_i_1__0_n_0;
  wire rem0_carry__0_i_1_n_0;
  wire rem0_carry__0_i_2__0_n_0;
  wire rem0_carry__0_i_2_n_0;
  wire rem0_carry__0_i_3__0_n_0;
  wire rem0_carry__0_i_3_n_0;
  wire rem0_carry__0_i_4__0_n_0;
  wire rem0_carry__0_i_4_n_0;
  wire rem0_carry__1_i_1__0_n_0;
  wire rem0_carry__1_i_1_n_0;
  wire rem0_carry__1_i_2__0_n_0;
  wire rem0_carry__1_i_2_n_0;
  wire rem0_carry__1_i_3__0_n_0;
  wire rem0_carry__1_i_3_n_0;
  wire rem0_carry__1_i_4__0_n_0;
  wire rem0_carry__1_i_4_n_0;
  wire rem0_carry__2_i_1__0_n_0;
  wire rem0_carry__2_i_1_n_0;
  wire rem0_carry__2_i_2__0_n_0;
  wire rem0_carry__2_i_2_n_0;
  wire rem0_carry__2_i_3__0_n_0;
  wire rem0_carry__2_i_3_n_0;
  wire rem0_carry__2_i_4__0_n_0;
  wire rem0_carry__2_i_4_n_0;
  wire rem0_carry__3_i_1__0_n_0;
  wire rem0_carry__3_i_1_n_0;
  wire rem0_carry__3_i_2__0_n_0;
  wire rem0_carry__3_i_2_n_0;
  wire rem0_carry__3_i_3__0_n_0;
  wire rem0_carry__3_i_3_n_0;
  wire rem0_carry__3_i_4__0_n_0;
  wire rem0_carry__3_i_4_n_0;
  wire rem0_carry__4_i_1__0_n_0;
  wire rem0_carry__4_i_1_n_0;
  wire rem0_carry__4_i_2__0_n_0;
  wire rem0_carry__4_i_2_n_0;
  wire rem0_carry__4_i_3__0_n_0;
  wire rem0_carry__4_i_3_n_0;
  wire rem0_carry__4_i_4__0_n_0;
  wire rem0_carry__4_i_4_n_0;
  wire rem0_carry__5_i_1__0_n_0;
  wire rem0_carry__5_i_1_n_0;
  wire rem0_carry__5_i_2__0_n_0;
  wire rem0_carry__5_i_2_n_0;
  wire rem0_carry__5_i_3__0_n_0;
  wire rem0_carry__5_i_3_n_0;
  wire rem0_carry__5_i_4__0_n_0;
  wire rem0_carry__5_i_4_n_0;
  wire rem0_carry__6_i_1__0_n_0;
  wire rem0_carry__6_i_1_n_0;
  wire rem0_carry__6_i_2__0_n_0;
  wire rem0_carry__6_i_2_n_0;
  wire rem0_carry__6_i_3__0_n_0;
  wire rem0_carry__6_i_3_n_0;
  wire rem0_carry__6_i_4__0_n_0;
  wire rem0_carry__6_i_4_n_0;
  wire rem0_carry__7_i_1__0_n_0;
  wire rem0_carry__7_i_1_n_0;
  wire rem0_carry_i_1__0_n_0;
  wire rem0_carry_i_1_n_0;
  wire rem0_carry_i_2__0_n_0;
  wire rem0_carry_i_2_n_0;
  wire rem0_carry_i_3__0_n_0;
  wire rem0_carry_i_3_n_0;
  wire rem0_carry_i_4__0_n_0;
  wire rem0_carry_i_4_n_0;
  wire rem0_carry_i_5__0_n_0;
  wire rem0_carry_i_5_n_0;
  wire rem1_carry__0_i_1__0_n_0;
  wire rem1_carry__0_i_1_n_0;
  wire rem1_carry__0_i_2__0_n_0;
  wire rem1_carry__0_i_2_n_0;
  wire rem1_carry__0_i_3__0_n_0;
  wire rem1_carry__0_i_3_n_0;
  wire rem1_carry__0_i_4__0_n_0;
  wire rem1_carry__0_i_4_n_0;
  wire rem1_carry__1_i_1__0_n_0;
  wire rem1_carry__1_i_1_n_0;
  wire rem1_carry__1_i_2__0_n_0;
  wire rem1_carry__1_i_2_n_0;
  wire rem1_carry__1_i_3__0_n_0;
  wire rem1_carry__1_i_3_n_0;
  wire rem1_carry__1_i_4__0_n_0;
  wire rem1_carry__1_i_4_n_0;
  wire rem1_carry__2_i_1__0_n_0;
  wire rem1_carry__2_i_1_n_0;
  wire rem1_carry__2_i_2__0_n_0;
  wire rem1_carry__2_i_2_n_0;
  wire rem1_carry__2_i_3__0_n_0;
  wire rem1_carry__2_i_3_n_0;
  wire rem1_carry__2_i_4__0_n_0;
  wire rem1_carry__2_i_4_n_0;
  wire rem1_carry__3_i_1__0_n_0;
  wire rem1_carry__3_i_1_n_0;
  wire rem1_carry__3_i_2__0_n_0;
  wire rem1_carry__3_i_2_n_0;
  wire rem1_carry__3_i_3__0_n_0;
  wire rem1_carry__3_i_3_n_0;
  wire rem1_carry__3_i_4__0_n_0;
  wire rem1_carry__3_i_4_n_0;
  wire rem1_carry__4_i_1__0_n_0;
  wire rem1_carry__4_i_1_n_0;
  wire rem1_carry__4_i_2__0_n_0;
  wire rem1_carry__4_i_2_n_0;
  wire rem1_carry__4_i_3__0_n_0;
  wire rem1_carry__4_i_3_n_0;
  wire rem1_carry__4_i_4__0_n_0;
  wire rem1_carry__4_i_4_n_0;
  wire rem1_carry__5_i_1__0_n_0;
  wire rem1_carry__5_i_1_n_0;
  wire rem1_carry__5_i_2__0_n_0;
  wire rem1_carry__5_i_2_n_0;
  wire rem1_carry__5_i_3__0_n_0;
  wire rem1_carry__5_i_3_n_0;
  wire rem1_carry__5_i_4__0_n_0;
  wire rem1_carry__5_i_4_n_0;
  wire rem1_carry__6_i_1__0_n_0;
  wire rem1_carry__6_i_1_n_0;
  wire rem1_carry__6_i_2__0_n_0;
  wire rem1_carry__6_i_2_n_0;
  wire rem1_carry__6_i_3__0_n_0;
  wire rem1_carry__6_i_3_n_0;
  wire rem1_carry__6_i_4__0_n_0;
  wire rem1_carry__6_i_4_n_0;
  wire rem1_carry__7_i_1__0_n_0;
  wire rem1_carry__7_i_1_n_0;
  wire rem1_carry_i_1__0_n_0;
  wire rem1_carry_i_1_n_0;
  wire rem1_carry_i_2__0_n_0;
  wire rem1_carry_i_2_n_0;
  wire rem1_carry_i_3__0_n_0;
  wire rem1_carry_i_3_n_0;
  wire rem1_carry_i_4__0_n_0;
  wire rem1_carry_i_4_n_0;
  wire rem1_carry_i_5__0_n_0;
  wire rem1_carry_i_5_n_0;
  wire rem2_carry__0_i_1__0_n_0;
  wire rem2_carry__0_i_1_n_0;
  wire rem2_carry__0_i_2__0_n_0;
  wire rem2_carry__0_i_2_n_0;
  wire rem2_carry__0_i_3__0_n_0;
  wire rem2_carry__0_i_3_n_0;
  wire rem2_carry__0_i_4__0_n_0;
  wire rem2_carry__0_i_4_n_0;
  wire rem2_carry__1_i_1__0_n_0;
  wire rem2_carry__1_i_1_n_0;
  wire rem2_carry__1_i_2__0_n_0;
  wire rem2_carry__1_i_2_n_0;
  wire rem2_carry__1_i_3__0_n_0;
  wire rem2_carry__1_i_3_n_0;
  wire rem2_carry__1_i_4__0_n_0;
  wire rem2_carry__1_i_4_n_0;
  wire rem2_carry__2_i_1__0_n_0;
  wire rem2_carry__2_i_1_n_0;
  wire rem2_carry__2_i_2__0_n_0;
  wire rem2_carry__2_i_2_n_0;
  wire rem2_carry__2_i_3__0_n_0;
  wire rem2_carry__2_i_3_n_0;
  wire rem2_carry__2_i_4__0_n_0;
  wire rem2_carry__2_i_4_n_0;
  wire rem2_carry__3_i_1__0_n_0;
  wire rem2_carry__3_i_1_n_0;
  wire rem2_carry__3_i_2__0_n_0;
  wire rem2_carry__3_i_2_n_0;
  wire rem2_carry__3_i_3__0_n_0;
  wire rem2_carry__3_i_3_n_0;
  wire rem2_carry__3_i_4__0_n_0;
  wire rem2_carry__3_i_4_n_0;
  wire rem2_carry__4_i_1__0_n_0;
  wire rem2_carry__4_i_1_n_0;
  wire rem2_carry__4_i_2__0_n_0;
  wire rem2_carry__4_i_2_n_0;
  wire rem2_carry__4_i_3__0_n_0;
  wire rem2_carry__4_i_3_n_0;
  wire rem2_carry__4_i_4__0_n_0;
  wire rem2_carry__4_i_4_n_0;
  wire rem2_carry__5_i_1__0_n_0;
  wire rem2_carry__5_i_1_n_0;
  wire rem2_carry__5_i_2__0_n_0;
  wire rem2_carry__5_i_2_n_0;
  wire rem2_carry__5_i_3__0_n_0;
  wire rem2_carry__5_i_3_n_0;
  wire rem2_carry__5_i_4__0_n_0;
  wire rem2_carry__5_i_4_n_0;
  wire rem2_carry__6_i_1__0_n_0;
  wire rem2_carry__6_i_1_n_0;
  wire rem2_carry__6_i_2__0_n_0;
  wire rem2_carry__6_i_2_n_0;
  wire rem2_carry__6_i_3__0_n_0;
  wire rem2_carry__6_i_3_n_0;
  wire rem2_carry__6_i_4__0_n_0;
  wire rem2_carry__6_i_4_n_0;
  wire rem2_carry__7_i_1__0_n_0;
  wire rem2_carry__7_i_1_n_0;
  wire rem2_carry_i_2__0_n_0;
  wire rem2_carry_i_2_n_0;
  wire rem2_carry_i_3__0_n_0;
  wire rem2_carry_i_3_n_0;
  wire rem2_carry_i_4__0_n_0;
  wire rem2_carry_i_4_n_0;
  wire rem2_carry_i_5__0_n_0;
  wire rem2_carry_i_5_n_0;
  wire rem3_carry__0_i_1__0_n_0;
  wire rem3_carry__0_i_1_n_0;
  wire rem3_carry__0_i_2__0_n_0;
  wire rem3_carry__0_i_2_n_0;
  wire rem3_carry__0_i_3__0_n_0;
  wire rem3_carry__0_i_3_n_0;
  wire rem3_carry__0_i_4__0_n_0;
  wire rem3_carry__0_i_4_n_0;
  wire rem3_carry__1_i_1__0_n_0;
  wire rem3_carry__1_i_1_n_0;
  wire rem3_carry__1_i_2__0_n_0;
  wire rem3_carry__1_i_2_n_0;
  wire rem3_carry__1_i_3__0_n_0;
  wire rem3_carry__1_i_3_n_0;
  wire rem3_carry__1_i_4__0_n_0;
  wire rem3_carry__1_i_4_n_0;
  wire rem3_carry__2_i_1__0_n_0;
  wire rem3_carry__2_i_1_n_0;
  wire rem3_carry__2_i_2__0_n_0;
  wire rem3_carry__2_i_2_n_0;
  wire rem3_carry__2_i_3__0_n_0;
  wire rem3_carry__2_i_3_n_0;
  wire rem3_carry__2_i_4__0_n_0;
  wire rem3_carry__2_i_4_n_0;
  wire rem3_carry__3_i_1__0_n_0;
  wire rem3_carry__3_i_1_n_0;
  wire rem3_carry__3_i_2__0_n_0;
  wire rem3_carry__3_i_2_n_0;
  wire rem3_carry__3_i_3__0_n_0;
  wire rem3_carry__3_i_3_n_0;
  wire rem3_carry__3_i_4__0_n_0;
  wire rem3_carry__3_i_4_n_0;
  wire rem3_carry__4_i_1__0_n_0;
  wire rem3_carry__4_i_1_n_0;
  wire rem3_carry__4_i_2__0_n_0;
  wire rem3_carry__4_i_2_n_0;
  wire rem3_carry__4_i_3__0_n_0;
  wire rem3_carry__4_i_3_n_0;
  wire rem3_carry__4_i_4__0_n_0;
  wire rem3_carry__4_i_4_n_0;
  wire rem3_carry__5_i_1__0_n_0;
  wire rem3_carry__5_i_1_n_0;
  wire rem3_carry__5_i_2__0_n_0;
  wire rem3_carry__5_i_2_n_0;
  wire rem3_carry__5_i_3__0_n_0;
  wire rem3_carry__5_i_3_n_0;
  wire rem3_carry__5_i_4__0_n_0;
  wire rem3_carry__5_i_4_n_0;
  wire rem3_carry__6_i_1__0_n_0;
  wire rem3_carry__6_i_1_n_0;
  wire rem3_carry__6_i_2__0_n_0;
  wire rem3_carry__6_i_2_n_0;
  wire rem3_carry__6_i_3__0_n_0;
  wire rem3_carry__6_i_3_n_0;
  wire rem3_carry__6_i_4__0_n_0;
  wire rem3_carry__6_i_4_n_0;
  wire rem3_carry__7_i_1__0_n_0;
  wire rem3_carry__7_i_1_n_0;
  wire rem3_carry_i_2__0_n_0;
  wire rem3_carry_i_2_n_0;
  wire rem3_carry_i_3__0_n_0;
  wire rem3_carry_i_3_n_0;
  wire rem3_carry_i_4__0_n_0;
  wire rem3_carry_i_4_n_0;
  wire rem3_carry_i_5__0_n_0;
  wire rem3_carry_i_5_n_0;
  wire \rem[11]_i_2__0_n_0 ;
  wire \rem[11]_i_2_n_0 ;
  wire \rem[11]_i_3__0_n_0 ;
  wire \rem[11]_i_3_n_0 ;
  wire \rem[11]_i_4__0_n_0 ;
  wire \rem[11]_i_4_n_0 ;
  wire \rem[11]_i_5__0_n_0 ;
  wire \rem[11]_i_5_n_0 ;
  wire \rem[11]_i_6__0_n_0 ;
  wire \rem[11]_i_6_n_0 ;
  wire \rem[11]_i_7__0_n_0 ;
  wire \rem[11]_i_7_n_0 ;
  wire \rem[11]_i_8__0_n_0 ;
  wire \rem[11]_i_8_n_0 ;
  wire \rem[11]_i_9__0_n_0 ;
  wire \rem[11]_i_9_n_0 ;
  wire \rem[15]_i_2__0_n_0 ;
  wire \rem[15]_i_2_n_0 ;
  wire \rem[15]_i_3__0_n_0 ;
  wire \rem[15]_i_3_n_0 ;
  wire \rem[15]_i_4__0_n_0 ;
  wire \rem[15]_i_4_n_0 ;
  wire \rem[15]_i_5__0_n_0 ;
  wire \rem[15]_i_5_n_0 ;
  wire \rem[15]_i_6__0_n_0 ;
  wire \rem[15]_i_6_n_0 ;
  wire \rem[15]_i_7__0_n_0 ;
  wire \rem[15]_i_7_n_0 ;
  wire \rem[15]_i_8__0_n_0 ;
  wire \rem[15]_i_8_n_0 ;
  wire \rem[15]_i_9__0_n_0 ;
  wire \rem[15]_i_9_n_0 ;
  wire \rem[19]_i_2__0_n_0 ;
  wire \rem[19]_i_2_n_0 ;
  wire \rem[19]_i_3__0_n_0 ;
  wire \rem[19]_i_3_n_0 ;
  wire \rem[19]_i_4__0_n_0 ;
  wire \rem[19]_i_4_n_0 ;
  wire \rem[19]_i_5__0_n_0 ;
  wire \rem[19]_i_5_n_0 ;
  wire \rem[19]_i_6__0_n_0 ;
  wire \rem[19]_i_6_n_0 ;
  wire \rem[19]_i_7__0_n_0 ;
  wire \rem[19]_i_7_n_0 ;
  wire \rem[19]_i_8__0_n_0 ;
  wire \rem[19]_i_8_n_0 ;
  wire \rem[19]_i_9__0_n_0 ;
  wire \rem[19]_i_9_n_0 ;
  wire \rem[23]_i_2__0_n_0 ;
  wire \rem[23]_i_2_n_0 ;
  wire \rem[23]_i_3__0_n_0 ;
  wire \rem[23]_i_3_n_0 ;
  wire \rem[23]_i_4__0_n_0 ;
  wire \rem[23]_i_4_n_0 ;
  wire \rem[23]_i_5__0_n_0 ;
  wire \rem[23]_i_5_n_0 ;
  wire \rem[23]_i_6__0_n_0 ;
  wire \rem[23]_i_6_n_0 ;
  wire \rem[23]_i_7__0_n_0 ;
  wire \rem[23]_i_7_n_0 ;
  wire \rem[23]_i_8__0_n_0 ;
  wire \rem[23]_i_8_n_0 ;
  wire \rem[23]_i_9__0_n_0 ;
  wire \rem[23]_i_9_n_0 ;
  wire \rem[27]_i_2__0_n_0 ;
  wire \rem[27]_i_2_n_0 ;
  wire \rem[27]_i_3__0_n_0 ;
  wire \rem[27]_i_3_n_0 ;
  wire \rem[27]_i_4__0_n_0 ;
  wire \rem[27]_i_4_n_0 ;
  wire \rem[27]_i_5__0_n_0 ;
  wire \rem[27]_i_5_n_0 ;
  wire \rem[27]_i_6__0_n_0 ;
  wire \rem[27]_i_6_n_0 ;
  wire \rem[27]_i_7__0_n_0 ;
  wire \rem[27]_i_7_n_0 ;
  wire \rem[27]_i_8__0_n_0 ;
  wire \rem[27]_i_8_n_0 ;
  wire \rem[27]_i_9__0_n_0 ;
  wire \rem[27]_i_9_n_0 ;
  wire \rem[31]_i_10__0_n_0 ;
  wire \rem[31]_i_10_n_0 ;
  wire \rem[31]_i_11__0_n_0 ;
  wire \rem[31]_i_11_n_0 ;
  wire \rem[31]_i_1__0_n_0 ;
  wire \rem[31]_i_1_n_0 ;
  wire \rem[31]_i_3__0_n_0 ;
  wire \rem[31]_i_3_n_0 ;
  wire \rem[31]_i_4__0_n_0 ;
  wire \rem[31]_i_4_n_0 ;
  wire \rem[31]_i_5__0_n_0 ;
  wire \rem[31]_i_5_n_0 ;
  wire \rem[31]_i_6__0_n_0 ;
  wire \rem[31]_i_6_n_0 ;
  wire \rem[31]_i_7__0_n_0 ;
  wire \rem[31]_i_7_n_0 ;
  wire \rem[31]_i_8__0_n_0 ;
  wire \rem[31]_i_8_n_0 ;
  wire \rem[31]_i_9__0_n_0 ;
  wire \rem[31]_i_9_n_0 ;
  wire \rem[3]_i_2__0_n_0 ;
  wire \rem[3]_i_2_n_0 ;
  wire \rem[3]_i_3__0_n_0 ;
  wire \rem[3]_i_3_n_0 ;
  wire \rem[3]_i_4__0_n_0 ;
  wire \rem[3]_i_4_n_0 ;
  wire \rem[3]_i_5__0_n_0 ;
  wire \rem[3]_i_5_n_0 ;
  wire \rem[3]_i_6__0_n_0 ;
  wire \rem[3]_i_6_n_0 ;
  wire \rem[3]_i_7__0_n_0 ;
  wire \rem[3]_i_7_n_0 ;
  wire \rem[3]_i_8__0_n_0 ;
  wire \rem[3]_i_8_n_0 ;
  wire \rem[3]_i_9__0_n_0 ;
  wire \rem[3]_i_9_n_0 ;
  wire \rem[7]_i_2__0_n_0 ;
  wire \rem[7]_i_2_n_0 ;
  wire \rem[7]_i_3__0_n_0 ;
  wire \rem[7]_i_3_n_0 ;
  wire \rem[7]_i_4__0_n_0 ;
  wire \rem[7]_i_4_n_0 ;
  wire \rem[7]_i_5__0_n_0 ;
  wire \rem[7]_i_5_n_0 ;
  wire \rem[7]_i_6__0_n_0 ;
  wire \rem[7]_i_6_n_0 ;
  wire \rem[7]_i_7__0_n_0 ;
  wire \rem[7]_i_7_n_0 ;
  wire \rem[7]_i_8__0_n_0 ;
  wire \rem[7]_i_8_n_0 ;
  wire \rem[7]_i_9__0_n_0 ;
  wire \rem[7]_i_9_n_0 ;
  wire \rem_reg[11]_i_1__0_n_0 ;
  wire \rem_reg[11]_i_1__0_n_1 ;
  wire \rem_reg[11]_i_1__0_n_2 ;
  wire \rem_reg[11]_i_1__0_n_3 ;
  wire \rem_reg[11]_i_1__0_n_4 ;
  wire \rem_reg[11]_i_1__0_n_5 ;
  wire \rem_reg[11]_i_1__0_n_6 ;
  wire \rem_reg[11]_i_1__0_n_7 ;
  wire \rem_reg[11]_i_1_n_0 ;
  wire \rem_reg[11]_i_1_n_1 ;
  wire \rem_reg[11]_i_1_n_2 ;
  wire \rem_reg[11]_i_1_n_3 ;
  wire \rem_reg[11]_i_1_n_4 ;
  wire \rem_reg[11]_i_1_n_5 ;
  wire \rem_reg[11]_i_1_n_6 ;
  wire \rem_reg[11]_i_1_n_7 ;
  wire \rem_reg[15]_i_1__0_n_0 ;
  wire \rem_reg[15]_i_1__0_n_1 ;
  wire \rem_reg[15]_i_1__0_n_2 ;
  wire \rem_reg[15]_i_1__0_n_3 ;
  wire \rem_reg[15]_i_1__0_n_4 ;
  wire \rem_reg[15]_i_1__0_n_5 ;
  wire \rem_reg[15]_i_1__0_n_6 ;
  wire \rem_reg[15]_i_1__0_n_7 ;
  wire \rem_reg[15]_i_1_n_0 ;
  wire \rem_reg[15]_i_1_n_1 ;
  wire \rem_reg[15]_i_1_n_2 ;
  wire \rem_reg[15]_i_1_n_3 ;
  wire \rem_reg[15]_i_1_n_4 ;
  wire \rem_reg[15]_i_1_n_5 ;
  wire \rem_reg[15]_i_1_n_6 ;
  wire \rem_reg[15]_i_1_n_7 ;
  wire \rem_reg[19]_i_1__0_n_0 ;
  wire \rem_reg[19]_i_1__0_n_1 ;
  wire \rem_reg[19]_i_1__0_n_2 ;
  wire \rem_reg[19]_i_1__0_n_3 ;
  wire \rem_reg[19]_i_1__0_n_4 ;
  wire \rem_reg[19]_i_1__0_n_5 ;
  wire \rem_reg[19]_i_1__0_n_6 ;
  wire \rem_reg[19]_i_1__0_n_7 ;
  wire \rem_reg[19]_i_1_n_0 ;
  wire \rem_reg[19]_i_1_n_1 ;
  wire \rem_reg[19]_i_1_n_2 ;
  wire \rem_reg[19]_i_1_n_3 ;
  wire \rem_reg[19]_i_1_n_4 ;
  wire \rem_reg[19]_i_1_n_5 ;
  wire \rem_reg[19]_i_1_n_6 ;
  wire \rem_reg[19]_i_1_n_7 ;
  wire \rem_reg[23]_i_1__0_n_0 ;
  wire \rem_reg[23]_i_1__0_n_1 ;
  wire \rem_reg[23]_i_1__0_n_2 ;
  wire \rem_reg[23]_i_1__0_n_3 ;
  wire \rem_reg[23]_i_1__0_n_4 ;
  wire \rem_reg[23]_i_1__0_n_5 ;
  wire \rem_reg[23]_i_1__0_n_6 ;
  wire \rem_reg[23]_i_1__0_n_7 ;
  wire \rem_reg[23]_i_1_n_0 ;
  wire \rem_reg[23]_i_1_n_1 ;
  wire \rem_reg[23]_i_1_n_2 ;
  wire \rem_reg[23]_i_1_n_3 ;
  wire \rem_reg[23]_i_1_n_4 ;
  wire \rem_reg[23]_i_1_n_5 ;
  wire \rem_reg[23]_i_1_n_6 ;
  wire \rem_reg[23]_i_1_n_7 ;
  wire \rem_reg[27]_i_1__0_n_0 ;
  wire \rem_reg[27]_i_1__0_n_1 ;
  wire \rem_reg[27]_i_1__0_n_2 ;
  wire \rem_reg[27]_i_1__0_n_3 ;
  wire \rem_reg[27]_i_1__0_n_4 ;
  wire \rem_reg[27]_i_1__0_n_5 ;
  wire \rem_reg[27]_i_1__0_n_6 ;
  wire \rem_reg[27]_i_1__0_n_7 ;
  wire \rem_reg[27]_i_1_n_0 ;
  wire \rem_reg[27]_i_1_n_1 ;
  wire \rem_reg[27]_i_1_n_2 ;
  wire \rem_reg[27]_i_1_n_3 ;
  wire \rem_reg[27]_i_1_n_4 ;
  wire \rem_reg[27]_i_1_n_5 ;
  wire \rem_reg[27]_i_1_n_6 ;
  wire \rem_reg[27]_i_1_n_7 ;
  wire \rem_reg[31]_i_2__0_n_1 ;
  wire \rem_reg[31]_i_2__0_n_2 ;
  wire \rem_reg[31]_i_2__0_n_3 ;
  wire \rem_reg[31]_i_2__0_n_4 ;
  wire \rem_reg[31]_i_2__0_n_5 ;
  wire \rem_reg[31]_i_2__0_n_6 ;
  wire \rem_reg[31]_i_2__0_n_7 ;
  wire \rem_reg[31]_i_2_n_1 ;
  wire \rem_reg[31]_i_2_n_2 ;
  wire \rem_reg[31]_i_2_n_3 ;
  wire \rem_reg[31]_i_2_n_4 ;
  wire \rem_reg[31]_i_2_n_5 ;
  wire \rem_reg[31]_i_2_n_6 ;
  wire \rem_reg[31]_i_2_n_7 ;
  wire \rem_reg[3]_i_1__0_n_0 ;
  wire \rem_reg[3]_i_1__0_n_1 ;
  wire \rem_reg[3]_i_1__0_n_2 ;
  wire \rem_reg[3]_i_1__0_n_3 ;
  wire \rem_reg[3]_i_1__0_n_4 ;
  wire \rem_reg[3]_i_1__0_n_5 ;
  wire \rem_reg[3]_i_1__0_n_6 ;
  wire \rem_reg[3]_i_1__0_n_7 ;
  wire \rem_reg[3]_i_1_n_0 ;
  wire \rem_reg[3]_i_1_n_1 ;
  wire \rem_reg[3]_i_1_n_2 ;
  wire \rem_reg[3]_i_1_n_3 ;
  wire \rem_reg[3]_i_1_n_4 ;
  wire \rem_reg[3]_i_1_n_5 ;
  wire \rem_reg[3]_i_1_n_6 ;
  wire \rem_reg[3]_i_1_n_7 ;
  wire \rem_reg[7]_i_1__0_n_0 ;
  wire \rem_reg[7]_i_1__0_n_1 ;
  wire \rem_reg[7]_i_1__0_n_2 ;
  wire \rem_reg[7]_i_1__0_n_3 ;
  wire \rem_reg[7]_i_1__0_n_4 ;
  wire \rem_reg[7]_i_1__0_n_5 ;
  wire \rem_reg[7]_i_1__0_n_6 ;
  wire \rem_reg[7]_i_1__0_n_7 ;
  wire \rem_reg[7]_i_1_n_0 ;
  wire \rem_reg[7]_i_1_n_1 ;
  wire \rem_reg[7]_i_1_n_2 ;
  wire \rem_reg[7]_i_1_n_3 ;
  wire \rem_reg[7]_i_1_n_4 ;
  wire \rem_reg[7]_i_1_n_5 ;
  wire \rem_reg[7]_i_1_n_6 ;
  wire \rem_reg[7]_i_1_n_7 ;
  wire \remden[0]_i_1__0_n_0 ;
  wire \remden[0]_i_1_n_0 ;
  wire \remden[10]_i_1__0_n_0 ;
  wire \remden[10]_i_1_n_0 ;
  wire \remden[11]_i_1__0_n_0 ;
  wire \remden[11]_i_1_n_0 ;
  wire \remden[12]_i_1__0_n_0 ;
  wire \remden[12]_i_1_n_0 ;
  wire \remden[13]_i_1__0_n_0 ;
  wire \remden[13]_i_1_n_0 ;
  wire \remden[14]_i_1__0_n_0 ;
  wire \remden[14]_i_1_n_0 ;
  wire \remden[15]_i_1__0_n_0 ;
  wire \remden[15]_i_1_n_0 ;
  wire \remden[16]_i_1__0_n_0 ;
  wire \remden[16]_i_1_n_0 ;
  wire \remden[16]_i_2__0_n_0 ;
  wire \remden[16]_i_2_n_0 ;
  wire \remden[17]_i_1__0_n_0 ;
  wire \remden[17]_i_1_n_0 ;
  wire \remden[17]_i_2__0_n_0 ;
  wire \remden[17]_i_2_n_0 ;
  wire \remden[18]_i_1__0_n_0 ;
  wire \remden[18]_i_1_n_0 ;
  wire \remden[18]_i_2__0_n_0 ;
  wire \remden[18]_i_2_n_0 ;
  wire \remden[19]_i_1__0_n_0 ;
  wire \remden[19]_i_1_n_0 ;
  wire \remden[19]_i_2__0_n_0 ;
  wire \remden[19]_i_2_n_0 ;
  wire \remden[1]_i_1__0_n_0 ;
  wire \remden[1]_i_1_n_0 ;
  wire \remden[20]_i_1__0_n_0 ;
  wire \remden[20]_i_1_n_0 ;
  wire \remden[20]_i_2__0_n_0 ;
  wire \remden[20]_i_2_n_0 ;
  wire \remden[21]_i_1__0_n_0 ;
  wire \remden[21]_i_1_n_0 ;
  wire \remden[21]_i_2__0_n_0 ;
  wire \remden[21]_i_2_n_0 ;
  wire \remden[22]_i_1__0_n_0 ;
  wire \remden[22]_i_1_n_0 ;
  wire \remden[22]_i_2__0_n_0 ;
  wire \remden[22]_i_2_n_0 ;
  wire \remden[23]_i_1__0_n_0 ;
  wire \remden[23]_i_1_n_0 ;
  wire \remden[23]_i_2__0_n_0 ;
  wire \remden[23]_i_2_n_0 ;
  wire \remden[24]_i_1__0_n_0 ;
  wire \remden[24]_i_1_n_0 ;
  wire \remden[24]_i_2__0_n_0 ;
  wire \remden[24]_i_2_n_0 ;
  wire \remden[25]_i_1__0_n_0 ;
  wire \remden[25]_i_1_n_0 ;
  wire \remden[25]_i_2__0_n_0 ;
  wire \remden[25]_i_2_n_0 ;
  wire \remden[26]_i_1__0_n_0 ;
  wire \remden[26]_i_1_n_0 ;
  wire \remden[26]_i_2__0_n_0 ;
  wire \remden[26]_i_2_n_0 ;
  wire \remden[27]_i_1__0_n_0 ;
  wire \remden[27]_i_1_n_0 ;
  wire \remden[27]_i_2__0_n_0 ;
  wire \remden[27]_i_2_n_0 ;
  wire \remden[28]_i_1__0_n_0 ;
  wire \remden[28]_i_1_n_0 ;
  wire \remden[28]_i_2__0_n_0 ;
  wire \remden[28]_i_2_n_0 ;
  wire \remden[29]_i_1__0_n_0 ;
  wire \remden[29]_i_1_n_0 ;
  wire \remden[29]_i_2__0_n_0 ;
  wire \remden[29]_i_2_n_0 ;
  wire \remden[2]_i_1__0_n_0 ;
  wire \remden[2]_i_1_n_0 ;
  wire \remden[30]_i_1__0_n_0 ;
  wire \remden[30]_i_1_n_0 ;
  wire \remden[30]_i_2__0_n_0 ;
  wire \remden[30]_i_2_n_0 ;
  wire \remden[31]_i_1__0_n_0 ;
  wire \remden[31]_i_1_n_0 ;
  wire \remden[31]_i_2__0_n_0 ;
  wire \remden[31]_i_2_n_0 ;
  wire \remden[31]_i_3_n_0 ;
  wire \remden[32]_i_1__0_n_0 ;
  wire \remden[32]_i_1_n_0 ;
  wire \remden[33]_i_1__0_n_0 ;
  wire \remden[33]_i_1_n_0 ;
  wire \remden[34]_i_1__0_n_0 ;
  wire \remden[34]_i_1_n_0 ;
  wire \remden[35]_i_1__0_n_0 ;
  wire \remden[35]_i_1_n_0 ;
  wire \remden[36]_i_1__0_n_0 ;
  wire \remden[36]_i_1_n_0 ;
  wire \remden[37]_i_1__0_n_0 ;
  wire \remden[37]_i_1_n_0 ;
  wire \remden[38]_i_1__0_n_0 ;
  wire \remden[38]_i_1_n_0 ;
  wire \remden[39]_i_1__0_n_0 ;
  wire \remden[39]_i_1_n_0 ;
  wire \remden[3]_i_1__0_n_0 ;
  wire \remden[3]_i_1_n_0 ;
  wire \remden[40]_i_1__0_n_0 ;
  wire \remden[40]_i_1_n_0 ;
  wire \remden[41]_i_1__0_n_0 ;
  wire \remden[41]_i_1_n_0 ;
  wire \remden[42]_i_1__0_n_0 ;
  wire \remden[42]_i_1_n_0 ;
  wire \remden[43]_i_1__0_n_0 ;
  wire \remden[43]_i_1_n_0 ;
  wire \remden[44]_i_1__0_n_0 ;
  wire \remden[44]_i_1_n_0 ;
  wire \remden[45]_i_1__0_n_0 ;
  wire \remden[45]_i_1_n_0 ;
  wire \remden[46]_i_1__0_n_0 ;
  wire \remden[46]_i_1_n_0 ;
  wire \remden[47]_i_1__0_n_0 ;
  wire \remden[47]_i_1_n_0 ;
  wire \remden[48]_i_1__0_n_0 ;
  wire \remden[48]_i_1_n_0 ;
  wire \remden[49]_i_1__0_n_0 ;
  wire \remden[49]_i_1_n_0 ;
  wire \remden[4]_i_1__0_n_0 ;
  wire \remden[4]_i_1_n_0 ;
  wire \remden[50]_i_1__0_n_0 ;
  wire \remden[50]_i_1_n_0 ;
  wire \remden[51]_i_1__0_n_0 ;
  wire \remden[51]_i_1_n_0 ;
  wire \remden[52]_i_1__0_n_0 ;
  wire \remden[52]_i_1_n_0 ;
  wire \remden[53]_i_1__0_n_0 ;
  wire \remden[53]_i_1_n_0 ;
  wire \remden[54]_i_1__0_n_0 ;
  wire \remden[54]_i_1_n_0 ;
  wire \remden[55]_i_1__0_n_0 ;
  wire \remden[55]_i_1_n_0 ;
  wire \remden[56]_i_1__0_n_0 ;
  wire \remden[56]_i_1_n_0 ;
  wire \remden[57]_i_1__0_n_0 ;
  wire \remden[57]_i_1_n_0 ;
  wire \remden[58]_i_1__0_n_0 ;
  wire \remden[58]_i_1_n_0 ;
  wire \remden[59]_i_1__0_n_0 ;
  wire \remden[59]_i_1_n_0 ;
  wire \remden[5]_i_1__0_n_0 ;
  wire \remden[5]_i_1_n_0 ;
  wire \remden[60]_i_1__0_n_0 ;
  wire \remden[60]_i_1_n_0 ;
  wire \remden[61]_i_1__0_n_0 ;
  wire \remden[61]_i_1_n_0 ;
  wire \remden[62]_i_1__0_n_0 ;
  wire \remden[62]_i_1_n_0 ;
  wire \remden[63]_i_1__0_n_0 ;
  wire \remden[63]_i_1_n_0 ;
  wire \remden[64]_i_1__0_n_0 ;
  wire \remden[64]_i_1_n_0 ;
  wire \remden[64]_i_2__0_n_0 ;
  wire \remden[64]_i_2_n_0 ;
  wire \remden[64]_i_3__0_n_0 ;
  wire \remden[64]_i_3_n_0 ;
  wire \remden[64]_i_4__0_n_0 ;
  wire \remden[64]_i_4_n_0 ;
  wire \remden[64]_i_5__0_n_0 ;
  wire \remden[64]_i_5_n_0 ;
  wire \remden[64]_i_6__0_n_0 ;
  wire \remden[64]_i_6_n_0 ;
  wire \remden[6]_i_1__0_n_0 ;
  wire \remden[6]_i_1_n_0 ;
  wire \remden[7]_i_1__0_n_0 ;
  wire \remden[7]_i_1_n_0 ;
  wire \remden[8]_i_1__0_n_0 ;
  wire \remden[8]_i_1_n_0 ;
  wire \remden[9]_i_1__0_n_0 ;
  wire \remden[9]_i_1_n_0 ;
  wire [15:0]\rgf/a0bus_b13 ;
  wire \rgf/a0bus_out/badr[0]_INST_0_i_12_n_0 ;
  wire \rgf/a0bus_out/badr[10]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[11]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[12]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[13]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[14]_INST_0_i_12_n_0 ;
  wire \rgf/a0bus_out/badr[15]_INST_0_i_13_n_0 ;
  wire \rgf/a0bus_out/badr[1]_INST_0_i_12_n_0 ;
  wire \rgf/a0bus_out/badr[2]_INST_0_i_12_n_0 ;
  wire \rgf/a0bus_out/badr[3]_INST_0_i_12_n_0 ;
  wire \rgf/a0bus_out/badr[4]_INST_0_i_12_n_0 ;
  wire \rgf/a0bus_out/badr[5]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[6]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[7]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[8]_INST_0_i_14_n_0 ;
  wire \rgf/a0bus_out/badr[9]_INST_0_i_14_n_0 ;
  wire [5:1]\rgf/a0bus_sel_cr ;
  wire [31:16]\rgf/a0bus_sp ;
  wire [15:0]\rgf/a0bus_sr ;
  wire [15:0]\rgf/a1bus_b02 ;
  wire [15:0]\rgf/a1bus_b13 ;
  wire \rgf/a1bus_out/badr[0]_INST_0_i_6_n_0 ;
  wire \rgf/a1bus_out/badr[10]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[11]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[12]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[13]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[14]_INST_0_i_3_n_0 ;
  wire \rgf/a1bus_out/badr[14]_INST_0_i_6_n_0 ;
  wire \rgf/a1bus_out/badr[15]_INST_0_i_3_n_0 ;
  wire \rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ;
  wire \rgf/a1bus_out/badr[1]_INST_0_i_3_n_0 ;
  wire \rgf/a1bus_out/badr[1]_INST_0_i_6_n_0 ;
  wire \rgf/a1bus_out/badr[2]_INST_0_i_3_n_0 ;
  wire \rgf/a1bus_out/badr[2]_INST_0_i_6_n_0 ;
  wire \rgf/a1bus_out/badr[3]_INST_0_i_3_n_0 ;
  wire \rgf/a1bus_out/badr[3]_INST_0_i_6_n_0 ;
  wire \rgf/a1bus_out/badr[4]_INST_0_i_3_n_0 ;
  wire \rgf/a1bus_out/badr[4]_INST_0_i_6_n_0 ;
  wire \rgf/a1bus_out/badr[5]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[6]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[7]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[8]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/badr[9]_INST_0_i_8_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[10]_i_32_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[10]_i_33_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[19]_i_39_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_45_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_46_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_47_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_48_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_49_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_50_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_51_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[28]_i_52_n_0 ;
  wire \rgf/a1bus_out/rgf_c1bus_wb[4]_i_28_n_0 ;
  wire [5:0]\rgf/a1bus_sel_cr ;
  wire [31:16]\rgf/a1bus_sp ;
  wire [15:0]\rgf/a1bus_sr ;
  wire \rgf/b0bus_out/bbus_o[0]_INST_0_i_17_n_0 ;
  wire \rgf/b0bus_out/bbus_o[0]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bbus_o[1]_INST_0_i_11_n_0 ;
  wire \rgf/b0bus_out/bbus_o[1]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[1]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[1]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bbus_o[2]_INST_0_i_11_n_0 ;
  wire \rgf/b0bus_out/bbus_o[2]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[2]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[2]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bbus_o[3]_INST_0_i_12_n_0 ;
  wire \rgf/b0bus_out/bbus_o[3]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[3]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[3]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bbus_o[4]_INST_0_i_11_n_0 ;
  wire \rgf/b0bus_out/bbus_o[4]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[4]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[4]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bbus_o[5]_INST_0_i_18_n_0 ;
  wire \rgf/b0bus_out/bbus_o[5]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[5]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bbus_o[5]_INST_0_i_6_n_0 ;
  wire \rgf/b0bus_out/bbus_o[6]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[6]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[6]_INST_0_i_8_n_0 ;
  wire \rgf/b0bus_out/bbus_o[7]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bbus_o[7]_INST_0_i_8_n_0 ;
  wire \rgf/b0bus_out/bdatw[10]_INST_0_i_10_n_0 ;
  wire \rgf/b0bus_out/bdatw[10]_INST_0_i_11_n_0 ;
  wire \rgf/b0bus_out/bdatw[10]_INST_0_i_22_n_0 ;
  wire \rgf/b0bus_out/bdatw[11]_INST_0_i_10_n_0 ;
  wire \rgf/b0bus_out/bdatw[11]_INST_0_i_11_n_0 ;
  wire \rgf/b0bus_out/bdatw[11]_INST_0_i_22_n_0 ;
  wire \rgf/b0bus_out/bdatw[12]_INST_0_i_10_n_0 ;
  wire \rgf/b0bus_out/bdatw[12]_INST_0_i_26_n_0 ;
  wire \rgf/b0bus_out/bdatw[12]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/bdatw[13]_INST_0_i_17_n_0 ;
  wire \rgf/b0bus_out/bdatw[13]_INST_0_i_8_n_0 ;
  wire \rgf/b0bus_out/bdatw[13]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/bdatw[14]_INST_0_i_10_n_0 ;
  wire \rgf/b0bus_out/bdatw[14]_INST_0_i_18_n_0 ;
  wire \rgf/b0bus_out/bdatw[14]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/bdatw[15]_INST_0_i_12_n_0 ;
  wire \rgf/b0bus_out/bdatw[15]_INST_0_i_13_n_0 ;
  wire \rgf/b0bus_out/bdatw[15]_INST_0_i_26_n_0 ;
  wire \rgf/b0bus_out/bdatw[16]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[16]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[17]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[17]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[18]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[18]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[19]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[19]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[20]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[20]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[21]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[21]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[22]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[22]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[23]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[23]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[24]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[24]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[25]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[25]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[26]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[26]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[27]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[27]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[28]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[28]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[29]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[29]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[30]_INST_0_i_3_n_0 ;
  wire \rgf/b0bus_out/bdatw[30]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[31]_INST_0_i_4_n_0 ;
  wire \rgf/b0bus_out/bdatw[31]_INST_0_i_5_n_0 ;
  wire \rgf/b0bus_out/bdatw[8]_INST_0_i_18_n_0 ;
  wire \rgf/b0bus_out/bdatw[8]_INST_0_i_7_n_0 ;
  wire \rgf/b0bus_out/bdatw[8]_INST_0_i_8_n_0 ;
  wire \rgf/b0bus_out/bdatw[9]_INST_0_i_20_n_0 ;
  wire \rgf/b0bus_out/bdatw[9]_INST_0_i_8_n_0 ;
  wire \rgf/b0bus_out/bdatw[9]_INST_0_i_9_n_0 ;
  wire \rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ;
  wire [7:0]\rgf/b0bus_sel_0 ;
  wire [5:0]\rgf/b0bus_sel_cr ;
  wire [0:0]\rgf/b0bus_sr ;
  wire [5:3]\rgf/b1bus_b02 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_14_n_0 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_7_n_0 ;
  wire \rgf/b1bus_out/bdatw[10]_INST_0_i_8_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_13_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_7_n_0 ;
  wire \rgf/b1bus_out/bdatw[11]_INST_0_i_8_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_12_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_15_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_19_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_38_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[12]_INST_0_i_7_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_12_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[13]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_11_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[14]_INST_0_i_7_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_10_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_15_n_0 ;
  wire \rgf/b1bus_out/bdatw[15]_INST_0_i_9_n_0 ;
  wire \rgf/b1bus_out/bdatw[16]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[16]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[17]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[17]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[18]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[18]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[19]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[19]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[20]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[20]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[21]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[21]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[22]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[22]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[23]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[23]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[24]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[24]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[25]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[25]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[26]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[26]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[27]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[27]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[28]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[28]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[29]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[29]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[30]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[30]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[31]_INST_0_i_10_n_0 ;
  wire \rgf/b1bus_out/bdatw[31]_INST_0_i_9_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_13_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[8]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_14_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/bdatw[9]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_17_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_3_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_17_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_3_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_19_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_3_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_6_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_7_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_8_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_10_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_5_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_7_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_3_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_4_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_8_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_3_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_4_n_0 ;
  wire \rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_8_n_0 ;
  wire \rgf/b1bus_out/rgf_c1bus_wb[31]_i_68_n_0 ;
  wire [7:0]\rgf/b1bus_sel_0 ;
  wire [5:0]\rgf/b1bus_sel_cr ;
  wire [5:0]\rgf/b1bus_sr ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_38_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_55_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso/i_/rgf_c1bus_wb[10]_i_34_n_0 ;
  wire \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_53_n_0 ;
  wire \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_55_n_0 ;
  wire \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_58_n_0 ;
  wire \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_62_n_0 ;
  wire \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_65_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_6_n_0 ;
  wire \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_62_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_54_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_55_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_73_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_50_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_53_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_79_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_81_n_0 ;
  wire \rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_84_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_8_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_33_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_34_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_52_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_53_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_72_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_41_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_49_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_76_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_80_n_0 ;
  wire \rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_83_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_31_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_32_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_46_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_47_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_69_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_22_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_27_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_28_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_71_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_40_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_4_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_9_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_13_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_7_n_0 ;
  wire \rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_80_n_0 ;
  wire \rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_81_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_29_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_30_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_35_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_37_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_44_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_68_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_10_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_36_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_25_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_26_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_42_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_70_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_39_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_14_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_15_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_16_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_5_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_17_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_18_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_20_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_21_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_6_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_11_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_12_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_19_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_6_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_79_n_0 ;
  wire \rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_82_n_0 ;
  wire \rgf/bank02/bank_sel00_out ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr00 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr01 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr02 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr03 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr04 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr05 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr06 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr07 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr20 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr21 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr22 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr23 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr24 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr25 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr26 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank02/gr27 ;
  wire \rgf/bank02/grn00/grn1__0 ;
  wire \rgf/bank02/grn01/grn1__0 ;
  wire \rgf/bank02/grn02/grn1__0 ;
  wire \rgf/bank02/grn03/grn1__0 ;
  wire \rgf/bank02/grn04/grn1__0 ;
  wire \rgf/bank02/grn05/grn1__0 ;
  wire \rgf/bank02/grn06/grn1__0 ;
  wire \rgf/bank02/grn07/grn1__0 ;
  wire \rgf/bank02/grn20/grn1__0 ;
  wire \rgf/bank02/grn21/grn1__0 ;
  wire \rgf/bank02/grn22/grn1__0 ;
  wire \rgf/bank02/grn23/grn1__0 ;
  wire \rgf/bank02/grn24/grn1__0 ;
  wire \rgf/bank02/grn25/grn1__0 ;
  wire \rgf/bank02/grn26/grn1__0 ;
  wire \rgf/bank02/grn27/grn1__0 ;
  wire [15:0]\rgf/bank02/p_0_in ;
  wire [13:5]\rgf/bank02/p_0_in0_in ;
  wire [15:0]\rgf/bank02/p_0_in2_in ;
  wire [15:0]\rgf/bank02/p_1_in ;
  wire [13:5]\rgf/bank02/p_1_in1_in ;
  wire [15:0]\rgf/bank02/p_1_in3_in ;
  wire \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_45_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_69_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_36_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[19]_i_43_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_57_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_59_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_64_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_66_n_0 ;
  wire \rgf/bank13/a1buso/i_/rgf_c1bus_wb[4]_i_29_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_6_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_7_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_8_n_0 ;
  wire \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_45_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_76_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_45_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_54_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_60_n_0 ;
  wire \rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_67_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_56_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_57_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_74_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_32_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_33_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_54_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_57_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_84_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_45_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_45_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_58_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_59_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_75_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_43_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_36_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_44_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_58_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_61_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_89_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_46_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_46_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_40_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_48_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_49_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_70_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_25_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_31_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_34_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_66_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_19_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_10_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_9_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_28_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_41_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_50_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_51_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_71_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_26_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_27_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_39_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_24_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_35_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_38_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_69_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_15_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_16_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_30_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_42_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_20_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_21_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_23_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_11_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_12_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_13_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_14_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_10_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_10_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_17_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_18_n_0 ;
  wire \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_22_n_0 ;
  wire \rgf/bank13/bank_sel00_out ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr00 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr01 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr02 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr03 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr04 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr05 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr06 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr07 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr20 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr21 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr22 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr23 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr24 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr25 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr26 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/bank13/gr27 ;
  wire \rgf/bank13/grn00/grn1__0 ;
  wire \rgf/bank13/grn01/grn1__0 ;
  wire \rgf/bank13/grn02/grn1__0 ;
  wire \rgf/bank13/grn03/grn1__0 ;
  wire \rgf/bank13/grn04/grn1__0 ;
  wire \rgf/bank13/grn05/grn1__0 ;
  wire \rgf/bank13/grn06/grn1__0 ;
  wire \rgf/bank13/grn07/grn1__0 ;
  wire \rgf/bank13/grn20/grn1__0 ;
  wire \rgf/bank13/grn21/grn1__0 ;
  wire \rgf/bank13/grn22/grn1__0 ;
  wire \rgf/bank13/grn23/grn1__0 ;
  wire \rgf/bank13/grn24/grn1__0 ;
  wire \rgf/bank13/grn25/grn1__0 ;
  wire \rgf/bank13/grn26/grn1__0 ;
  wire \rgf/bank13/grn27/grn1__0 ;
  wire [15:6]\rgf/bank13/p_0_in2_in ;
  wire [15:6]\rgf/bank13/p_1_in3_in ;
  wire [2:0]\rgf/bank_sel ;
  wire [15:15]\rgf/c0bus_bk2 ;
  wire [7:1]\rgf/c0bus_sel_0 ;
  wire [5:0]\rgf/c0bus_sel_cr ;
  wire [5:0]\rgf/c1bus_sel_cr ;
  (* DONT_TOUCH *) wire [15:0]\rgf/ivec/iv ;
  wire [15:0]\rgf/ivec/p_1_in ;
  wire [15:0]\rgf/p_2_in ;
  wire [15:0]\rgf/pcnt/p_1_in ;
  (* DONT_TOUCH *) wire [15:0]\rgf/pcnt/pc ;
  wire [4:0]\rgf/rctl/p_0_in ;
  wire \rgf/rctl/p_2_in ;
  wire [31:0]\rgf/rctl/rgf_c0bus_wb ;
  wire [31:0]\rgf/rctl/rgf_c1bus_wb ;
  wire [2:0]\rgf/rctl/rgf_selc0_rn_wb ;
  wire \rgf/rctl/rgf_selc0_stat ;
  wire [1:0]\rgf/rctl/rgf_selc0_wb ;
  wire [1:0]\rgf/rctl/rgf_selc1 ;
  wire [2:0]\rgf/rctl/rgf_selc1_rn ;
  wire [2:0]\rgf/rctl/rgf_selc1_rn_wb ;
  wire \rgf/rctl/rgf_selc1_stat ;
  wire [1:0]\rgf/rctl/rgf_selc1_wb ;
  wire [31:0]\rgf/rgf_c0bus_0 ;
  wire [31:0]\rgf/rgf_c1bus_0 ;
  wire \rgf/sptr/ctl_sp_id4 ;
  wire [31:0]\rgf/sptr/data2 ;
  wire [31:1]\rgf/sptr/data3 ;
  (* DONT_TOUCH *) wire [31:0]\rgf/sptr/sp ;
  wire [15:0]\rgf/sreg/p_0_in__0 ;
  (* DONT_TOUCH *) wire [15:0]\rgf/sreg/sr ;
  wire [31:0]\rgf/treg/p_1_in ;
  (* DONT_TOUCH *) wire [31:0]\rgf/treg/tr ;
  wire \rgf_c0bus_wb[0]_i_10_n_0 ;
  wire \rgf_c0bus_wb[0]_i_11_n_0 ;
  wire \rgf_c0bus_wb[0]_i_12_n_0 ;
  wire \rgf_c0bus_wb[0]_i_13_n_0 ;
  wire \rgf_c0bus_wb[0]_i_14_n_0 ;
  wire \rgf_c0bus_wb[0]_i_15_n_0 ;
  wire \rgf_c0bus_wb[0]_i_16_n_0 ;
  wire \rgf_c0bus_wb[0]_i_17_n_0 ;
  wire \rgf_c0bus_wb[0]_i_18_n_0 ;
  wire \rgf_c0bus_wb[0]_i_19_n_0 ;
  wire \rgf_c0bus_wb[0]_i_20_n_0 ;
  wire \rgf_c0bus_wb[0]_i_21_n_0 ;
  wire \rgf_c0bus_wb[0]_i_22_n_0 ;
  wire \rgf_c0bus_wb[0]_i_23_n_0 ;
  wire \rgf_c0bus_wb[0]_i_2_n_0 ;
  wire \rgf_c0bus_wb[0]_i_3_n_0 ;
  wire \rgf_c0bus_wb[0]_i_4_n_0 ;
  wire \rgf_c0bus_wb[0]_i_5_n_0 ;
  wire \rgf_c0bus_wb[0]_i_6_n_0 ;
  wire \rgf_c0bus_wb[0]_i_7_n_0 ;
  wire \rgf_c0bus_wb[0]_i_8_n_0 ;
  wire \rgf_c0bus_wb[0]_i_9_n_0 ;
  wire \rgf_c0bus_wb[10]_i_10_n_0 ;
  wire \rgf_c0bus_wb[10]_i_11_n_0 ;
  wire \rgf_c0bus_wb[10]_i_12_n_0 ;
  wire \rgf_c0bus_wb[10]_i_13_n_0 ;
  wire \rgf_c0bus_wb[10]_i_14_n_0 ;
  wire \rgf_c0bus_wb[10]_i_15_n_0 ;
  wire \rgf_c0bus_wb[10]_i_16_n_0 ;
  wire \rgf_c0bus_wb[10]_i_17_n_0 ;
  wire \rgf_c0bus_wb[10]_i_18_n_0 ;
  wire \rgf_c0bus_wb[10]_i_20_n_0 ;
  wire \rgf_c0bus_wb[10]_i_21_n_0 ;
  wire \rgf_c0bus_wb[10]_i_22_n_0 ;
  wire \rgf_c0bus_wb[10]_i_23_n_0 ;
  wire \rgf_c0bus_wb[10]_i_24_n_0 ;
  wire \rgf_c0bus_wb[10]_i_25_n_0 ;
  wire \rgf_c0bus_wb[10]_i_26_n_0 ;
  wire \rgf_c0bus_wb[10]_i_27_n_0 ;
  wire \rgf_c0bus_wb[10]_i_28_n_0 ;
  wire \rgf_c0bus_wb[10]_i_2_n_0 ;
  wire \rgf_c0bus_wb[10]_i_3_n_0 ;
  wire \rgf_c0bus_wb[10]_i_4_n_0 ;
  wire \rgf_c0bus_wb[10]_i_5_n_0 ;
  wire \rgf_c0bus_wb[10]_i_6_n_0 ;
  wire \rgf_c0bus_wb[10]_i_7_n_0 ;
  wire \rgf_c0bus_wb[10]_i_8_n_0 ;
  wire \rgf_c0bus_wb[10]_i_9_n_0 ;
  wire \rgf_c0bus_wb[11]_i_10_n_0 ;
  wire \rgf_c0bus_wb[11]_i_11_n_0 ;
  wire \rgf_c0bus_wb[11]_i_12_n_0 ;
  wire \rgf_c0bus_wb[11]_i_13_n_0 ;
  wire \rgf_c0bus_wb[11]_i_14_n_0 ;
  wire \rgf_c0bus_wb[11]_i_15_n_0 ;
  wire \rgf_c0bus_wb[11]_i_16_n_0 ;
  wire \rgf_c0bus_wb[11]_i_17_n_0 ;
  wire \rgf_c0bus_wb[11]_i_18_n_0 ;
  wire \rgf_c0bus_wb[11]_i_19_n_0 ;
  wire \rgf_c0bus_wb[11]_i_21_n_0 ;
  wire \rgf_c0bus_wb[11]_i_22_n_0 ;
  wire \rgf_c0bus_wb[11]_i_23_n_0 ;
  wire \rgf_c0bus_wb[11]_i_24_n_0 ;
  wire \rgf_c0bus_wb[11]_i_25_n_0 ;
  wire \rgf_c0bus_wb[11]_i_26_n_0 ;
  wire \rgf_c0bus_wb[11]_i_27_n_0 ;
  wire \rgf_c0bus_wb[11]_i_28_n_0 ;
  wire \rgf_c0bus_wb[11]_i_2_n_0 ;
  wire \rgf_c0bus_wb[11]_i_33_n_0 ;
  wire \rgf_c0bus_wb[11]_i_34_n_0 ;
  wire \rgf_c0bus_wb[11]_i_36_n_0 ;
  wire \rgf_c0bus_wb[11]_i_3_n_0 ;
  wire \rgf_c0bus_wb[11]_i_4_n_0 ;
  wire \rgf_c0bus_wb[11]_i_5_n_0 ;
  wire \rgf_c0bus_wb[11]_i_6_n_0 ;
  wire \rgf_c0bus_wb[11]_i_7_n_0 ;
  wire \rgf_c0bus_wb[11]_i_8_n_0 ;
  wire \rgf_c0bus_wb[11]_i_9_n_0 ;
  wire \rgf_c0bus_wb[12]_i_10_n_0 ;
  wire \rgf_c0bus_wb[12]_i_11_n_0 ;
  wire \rgf_c0bus_wb[12]_i_12_n_0 ;
  wire \rgf_c0bus_wb[12]_i_13_n_0 ;
  wire \rgf_c0bus_wb[12]_i_14_n_0 ;
  wire \rgf_c0bus_wb[12]_i_15_n_0 ;
  wire \rgf_c0bus_wb[12]_i_16_n_0 ;
  wire \rgf_c0bus_wb[12]_i_17_n_0 ;
  wire \rgf_c0bus_wb[12]_i_18_n_0 ;
  wire \rgf_c0bus_wb[12]_i_19_n_0 ;
  wire \rgf_c0bus_wb[12]_i_20_n_0 ;
  wire \rgf_c0bus_wb[12]_i_21_n_0 ;
  wire \rgf_c0bus_wb[12]_i_22_n_0 ;
  wire \rgf_c0bus_wb[12]_i_24_n_0 ;
  wire \rgf_c0bus_wb[12]_i_25_n_0 ;
  wire \rgf_c0bus_wb[12]_i_26_n_0 ;
  wire \rgf_c0bus_wb[12]_i_27_n_0 ;
  wire \rgf_c0bus_wb[12]_i_28_n_0 ;
  wire \rgf_c0bus_wb[12]_i_29_n_0 ;
  wire \rgf_c0bus_wb[12]_i_2_n_0 ;
  wire \rgf_c0bus_wb[12]_i_30_n_0 ;
  wire \rgf_c0bus_wb[12]_i_31_n_0 ;
  wire \rgf_c0bus_wb[12]_i_3_n_0 ;
  wire \rgf_c0bus_wb[12]_i_4_n_0 ;
  wire \rgf_c0bus_wb[12]_i_5_n_0 ;
  wire \rgf_c0bus_wb[12]_i_6_n_0 ;
  wire \rgf_c0bus_wb[12]_i_7_n_0 ;
  wire \rgf_c0bus_wb[12]_i_8_n_0 ;
  wire \rgf_c0bus_wb[12]_i_9_n_0 ;
  wire \rgf_c0bus_wb[13]_i_10_n_0 ;
  wire \rgf_c0bus_wb[13]_i_11_n_0 ;
  wire \rgf_c0bus_wb[13]_i_12_n_0 ;
  wire \rgf_c0bus_wb[13]_i_13_n_0 ;
  wire \rgf_c0bus_wb[13]_i_14_n_0 ;
  wire \rgf_c0bus_wb[13]_i_15_n_0 ;
  wire \rgf_c0bus_wb[13]_i_16_n_0 ;
  wire \rgf_c0bus_wb[13]_i_17_n_0 ;
  wire \rgf_c0bus_wb[13]_i_18_n_0 ;
  wire \rgf_c0bus_wb[13]_i_19_n_0 ;
  wire \rgf_c0bus_wb[13]_i_20_n_0 ;
  wire \rgf_c0bus_wb[13]_i_21_n_0 ;
  wire \rgf_c0bus_wb[13]_i_22_n_0 ;
  wire \rgf_c0bus_wb[13]_i_23_n_0 ;
  wire \rgf_c0bus_wb[13]_i_24_n_0 ;
  wire \rgf_c0bus_wb[13]_i_25_n_0 ;
  wire \rgf_c0bus_wb[13]_i_26_n_0 ;
  wire \rgf_c0bus_wb[13]_i_27_n_0 ;
  wire \rgf_c0bus_wb[13]_i_28_n_0 ;
  wire \rgf_c0bus_wb[13]_i_29_n_0 ;
  wire \rgf_c0bus_wb[13]_i_2_n_0 ;
  wire \rgf_c0bus_wb[13]_i_30_n_0 ;
  wire \rgf_c0bus_wb[13]_i_31_n_0 ;
  wire \rgf_c0bus_wb[13]_i_3_n_0 ;
  wire \rgf_c0bus_wb[13]_i_4_n_0 ;
  wire \rgf_c0bus_wb[13]_i_5_n_0 ;
  wire \rgf_c0bus_wb[13]_i_6_n_0 ;
  wire \rgf_c0bus_wb[13]_i_7_n_0 ;
  wire \rgf_c0bus_wb[13]_i_8_n_0 ;
  wire \rgf_c0bus_wb[13]_i_9_n_0 ;
  wire \rgf_c0bus_wb[14]_i_10_n_0 ;
  wire \rgf_c0bus_wb[14]_i_11_n_0 ;
  wire \rgf_c0bus_wb[14]_i_12_n_0 ;
  wire \rgf_c0bus_wb[14]_i_13_n_0 ;
  wire \rgf_c0bus_wb[14]_i_14_n_0 ;
  wire \rgf_c0bus_wb[14]_i_15_n_0 ;
  wire \rgf_c0bus_wb[14]_i_16_n_0 ;
  wire \rgf_c0bus_wb[14]_i_17_n_0 ;
  wire \rgf_c0bus_wb[14]_i_18_n_0 ;
  wire \rgf_c0bus_wb[14]_i_19_n_0 ;
  wire \rgf_c0bus_wb[14]_i_20_n_0 ;
  wire \rgf_c0bus_wb[14]_i_21_n_0 ;
  wire \rgf_c0bus_wb[14]_i_22_n_0 ;
  wire \rgf_c0bus_wb[14]_i_23_n_0 ;
  wire \rgf_c0bus_wb[14]_i_24_n_0 ;
  wire \rgf_c0bus_wb[14]_i_25_n_0 ;
  wire \rgf_c0bus_wb[14]_i_26_n_0 ;
  wire \rgf_c0bus_wb[14]_i_27_n_0 ;
  wire \rgf_c0bus_wb[14]_i_2_n_0 ;
  wire \rgf_c0bus_wb[14]_i_3_n_0 ;
  wire \rgf_c0bus_wb[14]_i_4_n_0 ;
  wire \rgf_c0bus_wb[14]_i_5_n_0 ;
  wire \rgf_c0bus_wb[14]_i_6_n_0 ;
  wire \rgf_c0bus_wb[14]_i_7_n_0 ;
  wire \rgf_c0bus_wb[14]_i_8_n_0 ;
  wire \rgf_c0bus_wb[14]_i_9_n_0 ;
  wire \rgf_c0bus_wb[15]_i_10_n_0 ;
  wire \rgf_c0bus_wb[15]_i_11_n_0 ;
  wire \rgf_c0bus_wb[15]_i_12_n_0 ;
  wire \rgf_c0bus_wb[15]_i_13_n_0 ;
  wire \rgf_c0bus_wb[15]_i_14_n_0 ;
  wire \rgf_c0bus_wb[15]_i_15_n_0 ;
  wire \rgf_c0bus_wb[15]_i_16_n_0 ;
  wire \rgf_c0bus_wb[15]_i_17_n_0 ;
  wire \rgf_c0bus_wb[15]_i_18_n_0 ;
  wire \rgf_c0bus_wb[15]_i_20_n_0 ;
  wire \rgf_c0bus_wb[15]_i_21_n_0 ;
  wire \rgf_c0bus_wb[15]_i_22_n_0 ;
  wire \rgf_c0bus_wb[15]_i_23_n_0 ;
  wire \rgf_c0bus_wb[15]_i_24_n_0 ;
  wire \rgf_c0bus_wb[15]_i_25_n_0 ;
  wire \rgf_c0bus_wb[15]_i_26_n_0 ;
  wire \rgf_c0bus_wb[15]_i_27_n_0 ;
  wire \rgf_c0bus_wb[15]_i_28_n_0 ;
  wire \rgf_c0bus_wb[15]_i_2_n_0 ;
  wire \rgf_c0bus_wb[15]_i_33_n_0 ;
  wire \rgf_c0bus_wb[15]_i_34_n_0 ;
  wire \rgf_c0bus_wb[15]_i_35_n_0 ;
  wire \rgf_c0bus_wb[15]_i_36_n_0 ;
  wire \rgf_c0bus_wb[15]_i_3_n_0 ;
  wire \rgf_c0bus_wb[15]_i_4_n_0 ;
  wire \rgf_c0bus_wb[15]_i_5_n_0 ;
  wire \rgf_c0bus_wb[15]_i_6_n_0 ;
  wire \rgf_c0bus_wb[15]_i_7_n_0 ;
  wire \rgf_c0bus_wb[15]_i_8_n_0 ;
  wire \rgf_c0bus_wb[15]_i_9_n_0 ;
  wire \rgf_c0bus_wb[16]_i_10_n_0 ;
  wire \rgf_c0bus_wb[16]_i_11_n_0 ;
  wire \rgf_c0bus_wb[16]_i_12_n_0 ;
  wire \rgf_c0bus_wb[16]_i_13_n_0 ;
  wire \rgf_c0bus_wb[16]_i_14_n_0 ;
  wire \rgf_c0bus_wb[16]_i_15_n_0 ;
  wire \rgf_c0bus_wb[16]_i_16_n_0 ;
  wire \rgf_c0bus_wb[16]_i_17_n_0 ;
  wire \rgf_c0bus_wb[16]_i_18_n_0 ;
  wire \rgf_c0bus_wb[16]_i_19_n_0 ;
  wire \rgf_c0bus_wb[16]_i_20_n_0 ;
  wire \rgf_c0bus_wb[16]_i_21_n_0 ;
  wire \rgf_c0bus_wb[16]_i_22_n_0 ;
  wire \rgf_c0bus_wb[16]_i_23_n_0 ;
  wire \rgf_c0bus_wb[16]_i_24_n_0 ;
  wire \rgf_c0bus_wb[16]_i_25_n_0 ;
  wire \rgf_c0bus_wb[16]_i_26_n_0 ;
  wire \rgf_c0bus_wb[16]_i_27_n_0 ;
  wire \rgf_c0bus_wb[16]_i_28_n_0 ;
  wire \rgf_c0bus_wb[16]_i_29_n_0 ;
  wire \rgf_c0bus_wb[16]_i_2_n_0 ;
  wire \rgf_c0bus_wb[16]_i_30_n_0 ;
  wire \rgf_c0bus_wb[16]_i_31_n_0 ;
  wire \rgf_c0bus_wb[16]_i_32_n_0 ;
  wire \rgf_c0bus_wb[16]_i_33_n_0 ;
  wire \rgf_c0bus_wb[16]_i_34_n_0 ;
  wire \rgf_c0bus_wb[16]_i_35_n_0 ;
  wire \rgf_c0bus_wb[16]_i_36_n_0 ;
  wire \rgf_c0bus_wb[16]_i_37_n_0 ;
  wire \rgf_c0bus_wb[16]_i_38_n_0 ;
  wire \rgf_c0bus_wb[16]_i_39_n_0 ;
  wire \rgf_c0bus_wb[16]_i_3_n_0 ;
  wire \rgf_c0bus_wb[16]_i_40_n_0 ;
  wire \rgf_c0bus_wb[16]_i_4_n_0 ;
  wire \rgf_c0bus_wb[16]_i_5_n_0 ;
  wire \rgf_c0bus_wb[16]_i_6_n_0 ;
  wire \rgf_c0bus_wb[16]_i_7_n_0 ;
  wire \rgf_c0bus_wb[16]_i_8_n_0 ;
  wire \rgf_c0bus_wb[16]_i_9_n_0 ;
  wire \rgf_c0bus_wb[17]_i_10_n_0 ;
  wire \rgf_c0bus_wb[17]_i_11_n_0 ;
  wire \rgf_c0bus_wb[17]_i_12_n_0 ;
  wire \rgf_c0bus_wb[17]_i_13_n_0 ;
  wire \rgf_c0bus_wb[17]_i_14_n_0 ;
  wire \rgf_c0bus_wb[17]_i_15_n_0 ;
  wire \rgf_c0bus_wb[17]_i_16_n_0 ;
  wire \rgf_c0bus_wb[17]_i_17_n_0 ;
  wire \rgf_c0bus_wb[17]_i_18_n_0 ;
  wire \rgf_c0bus_wb[17]_i_19_n_0 ;
  wire \rgf_c0bus_wb[17]_i_20_n_0 ;
  wire \rgf_c0bus_wb[17]_i_21_n_0 ;
  wire \rgf_c0bus_wb[17]_i_22_n_0 ;
  wire \rgf_c0bus_wb[17]_i_23_n_0 ;
  wire \rgf_c0bus_wb[17]_i_24_n_0 ;
  wire \rgf_c0bus_wb[17]_i_25_n_0 ;
  wire \rgf_c0bus_wb[17]_i_26_n_0 ;
  wire \rgf_c0bus_wb[17]_i_27_n_0 ;
  wire \rgf_c0bus_wb[17]_i_28_n_0 ;
  wire \rgf_c0bus_wb[17]_i_29_n_0 ;
  wire \rgf_c0bus_wb[17]_i_2_n_0 ;
  wire \rgf_c0bus_wb[17]_i_30_n_0 ;
  wire \rgf_c0bus_wb[17]_i_31_n_0 ;
  wire \rgf_c0bus_wb[17]_i_32_n_0 ;
  wire \rgf_c0bus_wb[17]_i_3_n_0 ;
  wire \rgf_c0bus_wb[17]_i_4_n_0 ;
  wire \rgf_c0bus_wb[17]_i_5_n_0 ;
  wire \rgf_c0bus_wb[17]_i_6_n_0 ;
  wire \rgf_c0bus_wb[17]_i_7_n_0 ;
  wire \rgf_c0bus_wb[17]_i_8_n_0 ;
  wire \rgf_c0bus_wb[17]_i_9_n_0 ;
  wire \rgf_c0bus_wb[18]_i_10_n_0 ;
  wire \rgf_c0bus_wb[18]_i_11_n_0 ;
  wire \rgf_c0bus_wb[18]_i_12_n_0 ;
  wire \rgf_c0bus_wb[18]_i_13_n_0 ;
  wire \rgf_c0bus_wb[18]_i_14_n_0 ;
  wire \rgf_c0bus_wb[18]_i_15_n_0 ;
  wire \rgf_c0bus_wb[18]_i_16_n_0 ;
  wire \rgf_c0bus_wb[18]_i_17_n_0 ;
  wire \rgf_c0bus_wb[18]_i_18_n_0 ;
  wire \rgf_c0bus_wb[18]_i_19_n_0 ;
  wire \rgf_c0bus_wb[18]_i_20_n_0 ;
  wire \rgf_c0bus_wb[18]_i_21_n_0 ;
  wire \rgf_c0bus_wb[18]_i_22_n_0 ;
  wire \rgf_c0bus_wb[18]_i_23_n_0 ;
  wire \rgf_c0bus_wb[18]_i_24_n_0 ;
  wire \rgf_c0bus_wb[18]_i_25_n_0 ;
  wire \rgf_c0bus_wb[18]_i_26_n_0 ;
  wire \rgf_c0bus_wb[18]_i_27_n_0 ;
  wire \rgf_c0bus_wb[18]_i_28_n_0 ;
  wire \rgf_c0bus_wb[18]_i_29_n_0 ;
  wire \rgf_c0bus_wb[18]_i_2_n_0 ;
  wire \rgf_c0bus_wb[18]_i_30_n_0 ;
  wire \rgf_c0bus_wb[18]_i_31_n_0 ;
  wire \rgf_c0bus_wb[18]_i_32_n_0 ;
  wire \rgf_c0bus_wb[18]_i_33_n_0 ;
  wire \rgf_c0bus_wb[18]_i_34_n_0 ;
  wire \rgf_c0bus_wb[18]_i_35_n_0 ;
  wire \rgf_c0bus_wb[18]_i_36_n_0 ;
  wire \rgf_c0bus_wb[18]_i_37_n_0 ;
  wire \rgf_c0bus_wb[18]_i_38_n_0 ;
  wire \rgf_c0bus_wb[18]_i_39_n_0 ;
  wire \rgf_c0bus_wb[18]_i_3_n_0 ;
  wire \rgf_c0bus_wb[18]_i_4_n_0 ;
  wire \rgf_c0bus_wb[18]_i_5_n_0 ;
  wire \rgf_c0bus_wb[18]_i_6_n_0 ;
  wire \rgf_c0bus_wb[18]_i_7_n_0 ;
  wire \rgf_c0bus_wb[18]_i_8_n_0 ;
  wire \rgf_c0bus_wb[18]_i_9_n_0 ;
  wire \rgf_c0bus_wb[19]_i_10_n_0 ;
  wire \rgf_c0bus_wb[19]_i_12_n_0 ;
  wire \rgf_c0bus_wb[19]_i_13_n_0 ;
  wire \rgf_c0bus_wb[19]_i_14_n_0 ;
  wire \rgf_c0bus_wb[19]_i_15_n_0 ;
  wire \rgf_c0bus_wb[19]_i_16_n_0 ;
  wire \rgf_c0bus_wb[19]_i_17_n_0 ;
  wire \rgf_c0bus_wb[19]_i_18_n_0 ;
  wire \rgf_c0bus_wb[19]_i_19_n_0 ;
  wire \rgf_c0bus_wb[19]_i_20_n_0 ;
  wire \rgf_c0bus_wb[19]_i_21_n_0 ;
  wire \rgf_c0bus_wb[19]_i_22_n_0 ;
  wire \rgf_c0bus_wb[19]_i_23_n_0 ;
  wire \rgf_c0bus_wb[19]_i_24_n_0 ;
  wire \rgf_c0bus_wb[19]_i_25_n_0 ;
  wire \rgf_c0bus_wb[19]_i_26_n_0 ;
  wire \rgf_c0bus_wb[19]_i_27_n_0 ;
  wire \rgf_c0bus_wb[19]_i_31_n_0 ;
  wire \rgf_c0bus_wb[19]_i_32_n_0 ;
  wire \rgf_c0bus_wb[19]_i_33_n_0 ;
  wire \rgf_c0bus_wb[19]_i_34_n_0 ;
  wire \rgf_c0bus_wb[19]_i_3_n_0 ;
  wire \rgf_c0bus_wb[19]_i_4_n_0 ;
  wire \rgf_c0bus_wb[19]_i_5_n_0 ;
  wire \rgf_c0bus_wb[19]_i_6_n_0 ;
  wire \rgf_c0bus_wb[19]_i_7_n_0 ;
  wire \rgf_c0bus_wb[19]_i_8_n_0 ;
  wire \rgf_c0bus_wb[19]_i_9_n_0 ;
  wire \rgf_c0bus_wb[1]_i_10_n_0 ;
  wire \rgf_c0bus_wb[1]_i_11_n_0 ;
  wire \rgf_c0bus_wb[1]_i_12_n_0 ;
  wire \rgf_c0bus_wb[1]_i_13_n_0 ;
  wire \rgf_c0bus_wb[1]_i_14_n_0 ;
  wire \rgf_c0bus_wb[1]_i_15_n_0 ;
  wire \rgf_c0bus_wb[1]_i_16_n_0 ;
  wire \rgf_c0bus_wb[1]_i_17_n_0 ;
  wire \rgf_c0bus_wb[1]_i_18_n_0 ;
  wire \rgf_c0bus_wb[1]_i_19_n_0 ;
  wire \rgf_c0bus_wb[1]_i_20_n_0 ;
  wire \rgf_c0bus_wb[1]_i_21_n_0 ;
  wire \rgf_c0bus_wb[1]_i_22_n_0 ;
  wire \rgf_c0bus_wb[1]_i_23_n_0 ;
  wire \rgf_c0bus_wb[1]_i_24_n_0 ;
  wire \rgf_c0bus_wb[1]_i_2_n_0 ;
  wire \rgf_c0bus_wb[1]_i_3_n_0 ;
  wire \rgf_c0bus_wb[1]_i_4_n_0 ;
  wire \rgf_c0bus_wb[1]_i_5_n_0 ;
  wire \rgf_c0bus_wb[1]_i_6_n_0 ;
  wire \rgf_c0bus_wb[1]_i_7_n_0 ;
  wire \rgf_c0bus_wb[1]_i_8_n_0 ;
  wire \rgf_c0bus_wb[1]_i_9_n_0 ;
  wire \rgf_c0bus_wb[20]_i_10_n_0 ;
  wire \rgf_c0bus_wb[20]_i_11_n_0 ;
  wire \rgf_c0bus_wb[20]_i_12_n_0 ;
  wire \rgf_c0bus_wb[20]_i_13_n_0 ;
  wire \rgf_c0bus_wb[20]_i_14_n_0 ;
  wire \rgf_c0bus_wb[20]_i_15_n_0 ;
  wire \rgf_c0bus_wb[20]_i_16_n_0 ;
  wire \rgf_c0bus_wb[20]_i_17_n_0 ;
  wire \rgf_c0bus_wb[20]_i_18_n_0 ;
  wire \rgf_c0bus_wb[20]_i_19_n_0 ;
  wire \rgf_c0bus_wb[20]_i_20_n_0 ;
  wire \rgf_c0bus_wb[20]_i_21_n_0 ;
  wire \rgf_c0bus_wb[20]_i_22_n_0 ;
  wire \rgf_c0bus_wb[20]_i_23_n_0 ;
  wire \rgf_c0bus_wb[20]_i_24_n_0 ;
  wire \rgf_c0bus_wb[20]_i_25_n_0 ;
  wire \rgf_c0bus_wb[20]_i_26_n_0 ;
  wire \rgf_c0bus_wb[20]_i_27_n_0 ;
  wire \rgf_c0bus_wb[20]_i_28_n_0 ;
  wire \rgf_c0bus_wb[20]_i_29_n_0 ;
  wire \rgf_c0bus_wb[20]_i_2_n_0 ;
  wire \rgf_c0bus_wb[20]_i_30_n_0 ;
  wire \rgf_c0bus_wb[20]_i_31_n_0 ;
  wire \rgf_c0bus_wb[20]_i_32_n_0 ;
  wire \rgf_c0bus_wb[20]_i_33_n_0 ;
  wire \rgf_c0bus_wb[20]_i_34_n_0 ;
  wire \rgf_c0bus_wb[20]_i_3_n_0 ;
  wire \rgf_c0bus_wb[20]_i_4_n_0 ;
  wire \rgf_c0bus_wb[20]_i_5_n_0 ;
  wire \rgf_c0bus_wb[20]_i_6_n_0 ;
  wire \rgf_c0bus_wb[20]_i_7_n_0 ;
  wire \rgf_c0bus_wb[20]_i_8_n_0 ;
  wire \rgf_c0bus_wb[20]_i_9_n_0 ;
  wire \rgf_c0bus_wb[21]_i_10_n_0 ;
  wire \rgf_c0bus_wb[21]_i_11_n_0 ;
  wire \rgf_c0bus_wb[21]_i_12_n_0 ;
  wire \rgf_c0bus_wb[21]_i_13_n_0 ;
  wire \rgf_c0bus_wb[21]_i_14_n_0 ;
  wire \rgf_c0bus_wb[21]_i_15_n_0 ;
  wire \rgf_c0bus_wb[21]_i_16_n_0 ;
  wire \rgf_c0bus_wb[21]_i_17_n_0 ;
  wire \rgf_c0bus_wb[21]_i_18_n_0 ;
  wire \rgf_c0bus_wb[21]_i_19_n_0 ;
  wire \rgf_c0bus_wb[21]_i_20_n_0 ;
  wire \rgf_c0bus_wb[21]_i_21_n_0 ;
  wire \rgf_c0bus_wb[21]_i_22_n_0 ;
  wire \rgf_c0bus_wb[21]_i_23_n_0 ;
  wire \rgf_c0bus_wb[21]_i_24_n_0 ;
  wire \rgf_c0bus_wb[21]_i_25_n_0 ;
  wire \rgf_c0bus_wb[21]_i_26_n_0 ;
  wire \rgf_c0bus_wb[21]_i_27_n_0 ;
  wire \rgf_c0bus_wb[21]_i_28_n_0 ;
  wire \rgf_c0bus_wb[21]_i_29_n_0 ;
  wire \rgf_c0bus_wb[21]_i_2_n_0 ;
  wire \rgf_c0bus_wb[21]_i_30_n_0 ;
  wire \rgf_c0bus_wb[21]_i_31_n_0 ;
  wire \rgf_c0bus_wb[21]_i_32_n_0 ;
  wire \rgf_c0bus_wb[21]_i_33_n_0 ;
  wire \rgf_c0bus_wb[21]_i_34_n_0 ;
  wire \rgf_c0bus_wb[21]_i_35_n_0 ;
  wire \rgf_c0bus_wb[21]_i_36_n_0 ;
  wire \rgf_c0bus_wb[21]_i_37_n_0 ;
  wire \rgf_c0bus_wb[21]_i_38_n_0 ;
  wire \rgf_c0bus_wb[21]_i_39_n_0 ;
  wire \rgf_c0bus_wb[21]_i_3_n_0 ;
  wire \rgf_c0bus_wb[21]_i_4_n_0 ;
  wire \rgf_c0bus_wb[21]_i_5_n_0 ;
  wire \rgf_c0bus_wb[21]_i_6_n_0 ;
  wire \rgf_c0bus_wb[21]_i_7_n_0 ;
  wire \rgf_c0bus_wb[21]_i_8_n_0 ;
  wire \rgf_c0bus_wb[21]_i_9_n_0 ;
  wire \rgf_c0bus_wb[22]_i_10_n_0 ;
  wire \rgf_c0bus_wb[22]_i_11_n_0 ;
  wire \rgf_c0bus_wb[22]_i_12_n_0 ;
  wire \rgf_c0bus_wb[22]_i_13_n_0 ;
  wire \rgf_c0bus_wb[22]_i_14_n_0 ;
  wire \rgf_c0bus_wb[22]_i_15_n_0 ;
  wire \rgf_c0bus_wb[22]_i_16_n_0 ;
  wire \rgf_c0bus_wb[22]_i_17_n_0 ;
  wire \rgf_c0bus_wb[22]_i_18_n_0 ;
  wire \rgf_c0bus_wb[22]_i_19_n_0 ;
  wire \rgf_c0bus_wb[22]_i_20_n_0 ;
  wire \rgf_c0bus_wb[22]_i_21_n_0 ;
  wire \rgf_c0bus_wb[22]_i_22_n_0 ;
  wire \rgf_c0bus_wb[22]_i_23_n_0 ;
  wire \rgf_c0bus_wb[22]_i_24_n_0 ;
  wire \rgf_c0bus_wb[22]_i_25_n_0 ;
  wire \rgf_c0bus_wb[22]_i_26_n_0 ;
  wire \rgf_c0bus_wb[22]_i_27_n_0 ;
  wire \rgf_c0bus_wb[22]_i_28_n_0 ;
  wire \rgf_c0bus_wb[22]_i_29_n_0 ;
  wire \rgf_c0bus_wb[22]_i_2_n_0 ;
  wire \rgf_c0bus_wb[22]_i_30_n_0 ;
  wire \rgf_c0bus_wb[22]_i_31_n_0 ;
  wire \rgf_c0bus_wb[22]_i_32_n_0 ;
  wire \rgf_c0bus_wb[22]_i_33_n_0 ;
  wire \rgf_c0bus_wb[22]_i_34_n_0 ;
  wire \rgf_c0bus_wb[22]_i_3_n_0 ;
  wire \rgf_c0bus_wb[22]_i_4_n_0 ;
  wire \rgf_c0bus_wb[22]_i_5_n_0 ;
  wire \rgf_c0bus_wb[22]_i_6_n_0 ;
  wire \rgf_c0bus_wb[22]_i_7_n_0 ;
  wire \rgf_c0bus_wb[22]_i_8_n_0 ;
  wire \rgf_c0bus_wb[22]_i_9_n_0 ;
  wire \rgf_c0bus_wb[23]_i_10_n_0 ;
  wire \rgf_c0bus_wb[23]_i_11_n_0 ;
  wire \rgf_c0bus_wb[23]_i_12_n_0 ;
  wire \rgf_c0bus_wb[23]_i_13_n_0 ;
  wire \rgf_c0bus_wb[23]_i_14_n_0 ;
  wire \rgf_c0bus_wb[23]_i_15_n_0 ;
  wire \rgf_c0bus_wb[23]_i_16_n_0 ;
  wire \rgf_c0bus_wb[23]_i_17_n_0 ;
  wire \rgf_c0bus_wb[23]_i_18_n_0 ;
  wire \rgf_c0bus_wb[23]_i_19_n_0 ;
  wire \rgf_c0bus_wb[23]_i_20_n_0 ;
  wire \rgf_c0bus_wb[23]_i_21_n_0 ;
  wire \rgf_c0bus_wb[23]_i_22_n_0 ;
  wire \rgf_c0bus_wb[23]_i_23_n_0 ;
  wire \rgf_c0bus_wb[23]_i_25_n_0 ;
  wire \rgf_c0bus_wb[23]_i_26_n_0 ;
  wire \rgf_c0bus_wb[23]_i_27_n_0 ;
  wire \rgf_c0bus_wb[23]_i_28_n_0 ;
  wire \rgf_c0bus_wb[23]_i_29_n_0 ;
  wire \rgf_c0bus_wb[23]_i_2_n_0 ;
  wire \rgf_c0bus_wb[23]_i_30_n_0 ;
  wire \rgf_c0bus_wb[23]_i_31_n_0 ;
  wire \rgf_c0bus_wb[23]_i_32_n_0 ;
  wire \rgf_c0bus_wb[23]_i_33_n_0 ;
  wire \rgf_c0bus_wb[23]_i_34_n_0 ;
  wire \rgf_c0bus_wb[23]_i_35_n_0 ;
  wire \rgf_c0bus_wb[23]_i_36_n_0 ;
  wire \rgf_c0bus_wb[23]_i_37_n_0 ;
  wire \rgf_c0bus_wb[23]_i_3_n_0 ;
  wire \rgf_c0bus_wb[23]_i_40_n_0 ;
  wire \rgf_c0bus_wb[23]_i_41_n_0 ;
  wire \rgf_c0bus_wb[23]_i_4_n_0 ;
  wire \rgf_c0bus_wb[23]_i_5_n_0 ;
  wire \rgf_c0bus_wb[23]_i_6_n_0 ;
  wire \rgf_c0bus_wb[23]_i_7_n_0 ;
  wire \rgf_c0bus_wb[23]_i_8_n_0 ;
  wire \rgf_c0bus_wb[23]_i_9_n_0 ;
  wire \rgf_c0bus_wb[24]_i_10_n_0 ;
  wire \rgf_c0bus_wb[24]_i_11_n_0 ;
  wire \rgf_c0bus_wb[24]_i_12_n_0 ;
  wire \rgf_c0bus_wb[24]_i_13_n_0 ;
  wire \rgf_c0bus_wb[24]_i_14_n_0 ;
  wire \rgf_c0bus_wb[24]_i_15_n_0 ;
  wire \rgf_c0bus_wb[24]_i_16_n_0 ;
  wire \rgf_c0bus_wb[24]_i_17_n_0 ;
  wire \rgf_c0bus_wb[24]_i_18_n_0 ;
  wire \rgf_c0bus_wb[24]_i_19_n_0 ;
  wire \rgf_c0bus_wb[24]_i_20_n_0 ;
  wire \rgf_c0bus_wb[24]_i_21_n_0 ;
  wire \rgf_c0bus_wb[24]_i_22_n_0 ;
  wire \rgf_c0bus_wb[24]_i_23_n_0 ;
  wire \rgf_c0bus_wb[24]_i_24_n_0 ;
  wire \rgf_c0bus_wb[24]_i_25_n_0 ;
  wire \rgf_c0bus_wb[24]_i_26_n_0 ;
  wire \rgf_c0bus_wb[24]_i_27_n_0 ;
  wire \rgf_c0bus_wb[24]_i_28_n_0 ;
  wire \rgf_c0bus_wb[24]_i_29_n_0 ;
  wire \rgf_c0bus_wb[24]_i_30_n_0 ;
  wire \rgf_c0bus_wb[24]_i_3_n_0 ;
  wire \rgf_c0bus_wb[24]_i_4_n_0 ;
  wire \rgf_c0bus_wb[24]_i_5_n_0 ;
  wire \rgf_c0bus_wb[24]_i_6_n_0 ;
  wire \rgf_c0bus_wb[24]_i_7_n_0 ;
  wire \rgf_c0bus_wb[24]_i_8_n_0 ;
  wire \rgf_c0bus_wb[24]_i_9_n_0 ;
  wire \rgf_c0bus_wb[25]_i_10_n_0 ;
  wire \rgf_c0bus_wb[25]_i_11_n_0 ;
  wire \rgf_c0bus_wb[25]_i_12_n_0 ;
  wire \rgf_c0bus_wb[25]_i_13_n_0 ;
  wire \rgf_c0bus_wb[25]_i_14_n_0 ;
  wire \rgf_c0bus_wb[25]_i_15_n_0 ;
  wire \rgf_c0bus_wb[25]_i_16_n_0 ;
  wire \rgf_c0bus_wb[25]_i_17_n_0 ;
  wire \rgf_c0bus_wb[25]_i_18_n_0 ;
  wire \rgf_c0bus_wb[25]_i_19_n_0 ;
  wire \rgf_c0bus_wb[25]_i_20_n_0 ;
  wire \rgf_c0bus_wb[25]_i_21_n_0 ;
  wire \rgf_c0bus_wb[25]_i_22_n_0 ;
  wire \rgf_c0bus_wb[25]_i_23_n_0 ;
  wire \rgf_c0bus_wb[25]_i_24_n_0 ;
  wire \rgf_c0bus_wb[25]_i_25_n_0 ;
  wire \rgf_c0bus_wb[25]_i_26_n_0 ;
  wire \rgf_c0bus_wb[25]_i_27_n_0 ;
  wire \rgf_c0bus_wb[25]_i_28_n_0 ;
  wire \rgf_c0bus_wb[25]_i_29_n_0 ;
  wire \rgf_c0bus_wb[25]_i_2_n_0 ;
  wire \rgf_c0bus_wb[25]_i_30_n_0 ;
  wire \rgf_c0bus_wb[25]_i_31_n_0 ;
  wire \rgf_c0bus_wb[25]_i_32_n_0 ;
  wire \rgf_c0bus_wb[25]_i_33_n_0 ;
  wire \rgf_c0bus_wb[25]_i_34_n_0 ;
  wire \rgf_c0bus_wb[25]_i_35_n_0 ;
  wire \rgf_c0bus_wb[25]_i_36_n_0 ;
  wire \rgf_c0bus_wb[25]_i_37_n_0 ;
  wire \rgf_c0bus_wb[25]_i_38_n_0 ;
  wire \rgf_c0bus_wb[25]_i_39_n_0 ;
  wire \rgf_c0bus_wb[25]_i_3_n_0 ;
  wire \rgf_c0bus_wb[25]_i_40_n_0 ;
  wire \rgf_c0bus_wb[25]_i_41_n_0 ;
  wire \rgf_c0bus_wb[25]_i_42_n_0 ;
  wire \rgf_c0bus_wb[25]_i_43_n_0 ;
  wire \rgf_c0bus_wb[25]_i_44_n_0 ;
  wire \rgf_c0bus_wb[25]_i_4_n_0 ;
  wire \rgf_c0bus_wb[25]_i_5_n_0 ;
  wire \rgf_c0bus_wb[25]_i_6_n_0 ;
  wire \rgf_c0bus_wb[25]_i_7_n_0 ;
  wire \rgf_c0bus_wb[25]_i_8_n_0 ;
  wire \rgf_c0bus_wb[25]_i_9_n_0 ;
  wire \rgf_c0bus_wb[26]_i_10_n_0 ;
  wire \rgf_c0bus_wb[26]_i_11_n_0 ;
  wire \rgf_c0bus_wb[26]_i_12_n_0 ;
  wire \rgf_c0bus_wb[26]_i_13_n_0 ;
  wire \rgf_c0bus_wb[26]_i_14_n_0 ;
  wire \rgf_c0bus_wb[26]_i_15_n_0 ;
  wire \rgf_c0bus_wb[26]_i_16_n_0 ;
  wire \rgf_c0bus_wb[26]_i_17_n_0 ;
  wire \rgf_c0bus_wb[26]_i_18_n_0 ;
  wire \rgf_c0bus_wb[26]_i_19_n_0 ;
  wire \rgf_c0bus_wb[26]_i_20_n_0 ;
  wire \rgf_c0bus_wb[26]_i_21_n_0 ;
  wire \rgf_c0bus_wb[26]_i_22_n_0 ;
  wire \rgf_c0bus_wb[26]_i_23_n_0 ;
  wire \rgf_c0bus_wb[26]_i_24_n_0 ;
  wire \rgf_c0bus_wb[26]_i_3_n_0 ;
  wire \rgf_c0bus_wb[26]_i_4_n_0 ;
  wire \rgf_c0bus_wb[26]_i_5_n_0 ;
  wire \rgf_c0bus_wb[26]_i_6_n_0 ;
  wire \rgf_c0bus_wb[26]_i_7_n_0 ;
  wire \rgf_c0bus_wb[26]_i_8_n_0 ;
  wire \rgf_c0bus_wb[26]_i_9_n_0 ;
  wire \rgf_c0bus_wb[27]_i_10_n_0 ;
  wire \rgf_c0bus_wb[27]_i_11_n_0 ;
  wire \rgf_c0bus_wb[27]_i_12_n_0 ;
  wire \rgf_c0bus_wb[27]_i_13_n_0 ;
  wire \rgf_c0bus_wb[27]_i_14_n_0 ;
  wire \rgf_c0bus_wb[27]_i_15_n_0 ;
  wire \rgf_c0bus_wb[27]_i_16_n_0 ;
  wire \rgf_c0bus_wb[27]_i_17_n_0 ;
  wire \rgf_c0bus_wb[27]_i_18_n_0 ;
  wire \rgf_c0bus_wb[27]_i_19_n_0 ;
  wire \rgf_c0bus_wb[27]_i_20_n_0 ;
  wire \rgf_c0bus_wb[27]_i_21_n_0 ;
  wire \rgf_c0bus_wb[27]_i_22_n_0 ;
  wire \rgf_c0bus_wb[27]_i_24_n_0 ;
  wire \rgf_c0bus_wb[27]_i_25_n_0 ;
  wire \rgf_c0bus_wb[27]_i_26_n_0 ;
  wire \rgf_c0bus_wb[27]_i_27_n_0 ;
  wire \rgf_c0bus_wb[27]_i_28_n_0 ;
  wire \rgf_c0bus_wb[27]_i_29_n_0 ;
  wire \rgf_c0bus_wb[27]_i_2_n_0 ;
  wire \rgf_c0bus_wb[27]_i_30_n_0 ;
  wire \rgf_c0bus_wb[27]_i_31_n_0 ;
  wire \rgf_c0bus_wb[27]_i_32_n_0 ;
  wire \rgf_c0bus_wb[27]_i_33_n_0 ;
  wire \rgf_c0bus_wb[27]_i_34_n_0 ;
  wire \rgf_c0bus_wb[27]_i_35_n_0 ;
  wire \rgf_c0bus_wb[27]_i_36_n_0 ;
  wire \rgf_c0bus_wb[27]_i_37_n_0 ;
  wire \rgf_c0bus_wb[27]_i_38_n_0 ;
  wire \rgf_c0bus_wb[27]_i_39_n_0 ;
  wire \rgf_c0bus_wb[27]_i_3_n_0 ;
  wire \rgf_c0bus_wb[27]_i_42_n_0 ;
  wire \rgf_c0bus_wb[27]_i_43_n_0 ;
  wire \rgf_c0bus_wb[27]_i_44_n_0 ;
  wire \rgf_c0bus_wb[27]_i_45_n_0 ;
  wire \rgf_c0bus_wb[27]_i_46_n_0 ;
  wire \rgf_c0bus_wb[27]_i_4_n_0 ;
  wire \rgf_c0bus_wb[27]_i_5_n_0 ;
  wire \rgf_c0bus_wb[27]_i_6_n_0 ;
  wire \rgf_c0bus_wb[27]_i_7_n_0 ;
  wire \rgf_c0bus_wb[27]_i_8_n_0 ;
  wire \rgf_c0bus_wb[27]_i_9_n_0 ;
  wire \rgf_c0bus_wb[28]_i_10_n_0 ;
  wire \rgf_c0bus_wb[28]_i_11_n_0 ;
  wire \rgf_c0bus_wb[28]_i_12_n_0 ;
  wire \rgf_c0bus_wb[28]_i_13_n_0 ;
  wire \rgf_c0bus_wb[28]_i_14_n_0 ;
  wire \rgf_c0bus_wb[28]_i_15_n_0 ;
  wire \rgf_c0bus_wb[28]_i_16_n_0 ;
  wire \rgf_c0bus_wb[28]_i_17_n_0 ;
  wire \rgf_c0bus_wb[28]_i_18_n_0 ;
  wire \rgf_c0bus_wb[28]_i_19_n_0 ;
  wire \rgf_c0bus_wb[28]_i_20_n_0 ;
  wire \rgf_c0bus_wb[28]_i_21_n_0 ;
  wire \rgf_c0bus_wb[28]_i_22_n_0 ;
  wire \rgf_c0bus_wb[28]_i_23_n_0 ;
  wire \rgf_c0bus_wb[28]_i_24_n_0 ;
  wire \rgf_c0bus_wb[28]_i_25_n_0 ;
  wire \rgf_c0bus_wb[28]_i_26_n_0 ;
  wire \rgf_c0bus_wb[28]_i_27_n_0 ;
  wire \rgf_c0bus_wb[28]_i_28_n_0 ;
  wire \rgf_c0bus_wb[28]_i_29_n_0 ;
  wire \rgf_c0bus_wb[28]_i_2_n_0 ;
  wire \rgf_c0bus_wb[28]_i_30_n_0 ;
  wire \rgf_c0bus_wb[28]_i_31_n_0 ;
  wire \rgf_c0bus_wb[28]_i_32_n_0 ;
  wire \rgf_c0bus_wb[28]_i_33_n_0 ;
  wire \rgf_c0bus_wb[28]_i_34_n_0 ;
  wire \rgf_c0bus_wb[28]_i_35_n_0 ;
  wire \rgf_c0bus_wb[28]_i_36_n_0 ;
  wire \rgf_c0bus_wb[28]_i_37_n_0 ;
  wire \rgf_c0bus_wb[28]_i_38_n_0 ;
  wire \rgf_c0bus_wb[28]_i_39_n_0 ;
  wire \rgf_c0bus_wb[28]_i_3_n_0 ;
  wire \rgf_c0bus_wb[28]_i_40_n_0 ;
  wire \rgf_c0bus_wb[28]_i_41_n_0 ;
  wire \rgf_c0bus_wb[28]_i_42_n_0 ;
  wire \rgf_c0bus_wb[28]_i_43_n_0 ;
  wire \rgf_c0bus_wb[28]_i_44_n_0 ;
  wire \rgf_c0bus_wb[28]_i_4_n_0 ;
  wire \rgf_c0bus_wb[28]_i_5_n_0 ;
  wire \rgf_c0bus_wb[28]_i_6_n_0 ;
  wire \rgf_c0bus_wb[28]_i_7_n_0 ;
  wire \rgf_c0bus_wb[28]_i_8_n_0 ;
  wire \rgf_c0bus_wb[28]_i_9_n_0 ;
  wire \rgf_c0bus_wb[29]_i_10_n_0 ;
  wire \rgf_c0bus_wb[29]_i_12_n_0 ;
  wire \rgf_c0bus_wb[29]_i_13_n_0 ;
  wire \rgf_c0bus_wb[29]_i_14_n_0 ;
  wire \rgf_c0bus_wb[29]_i_15_n_0 ;
  wire \rgf_c0bus_wb[29]_i_16_n_0 ;
  wire \rgf_c0bus_wb[29]_i_17_n_0 ;
  wire \rgf_c0bus_wb[29]_i_18_n_0 ;
  wire \rgf_c0bus_wb[29]_i_19_n_0 ;
  wire \rgf_c0bus_wb[29]_i_20_n_0 ;
  wire \rgf_c0bus_wb[29]_i_21_n_0 ;
  wire \rgf_c0bus_wb[29]_i_22_n_0 ;
  wire \rgf_c0bus_wb[29]_i_23_n_0 ;
  wire \rgf_c0bus_wb[29]_i_24_n_0 ;
  wire \rgf_c0bus_wb[29]_i_25_n_0 ;
  wire \rgf_c0bus_wb[29]_i_26_n_0 ;
  wire \rgf_c0bus_wb[29]_i_27_n_0 ;
  wire \rgf_c0bus_wb[29]_i_28_n_0 ;
  wire \rgf_c0bus_wb[29]_i_31_n_0 ;
  wire \rgf_c0bus_wb[29]_i_32_n_0 ;
  wire \rgf_c0bus_wb[29]_i_33_n_0 ;
  wire \rgf_c0bus_wb[29]_i_34_n_0 ;
  wire \rgf_c0bus_wb[29]_i_3_n_0 ;
  wire \rgf_c0bus_wb[29]_i_4_n_0 ;
  wire \rgf_c0bus_wb[29]_i_5_n_0 ;
  wire \rgf_c0bus_wb[29]_i_6_n_0 ;
  wire \rgf_c0bus_wb[29]_i_7_n_0 ;
  wire \rgf_c0bus_wb[29]_i_8_n_0 ;
  wire \rgf_c0bus_wb[29]_i_9_n_0 ;
  wire \rgf_c0bus_wb[2]_i_10_n_0 ;
  wire \rgf_c0bus_wb[2]_i_11_n_0 ;
  wire \rgf_c0bus_wb[2]_i_12_n_0 ;
  wire \rgf_c0bus_wb[2]_i_13_n_0 ;
  wire \rgf_c0bus_wb[2]_i_14_n_0 ;
  wire \rgf_c0bus_wb[2]_i_15_n_0 ;
  wire \rgf_c0bus_wb[2]_i_16_n_0 ;
  wire \rgf_c0bus_wb[2]_i_17_n_0 ;
  wire \rgf_c0bus_wb[2]_i_18_n_0 ;
  wire \rgf_c0bus_wb[2]_i_19_n_0 ;
  wire \rgf_c0bus_wb[2]_i_20_n_0 ;
  wire \rgf_c0bus_wb[2]_i_21_n_0 ;
  wire \rgf_c0bus_wb[2]_i_22_n_0 ;
  wire \rgf_c0bus_wb[2]_i_23_n_0 ;
  wire \rgf_c0bus_wb[2]_i_24_n_0 ;
  wire \rgf_c0bus_wb[2]_i_25_n_0 ;
  wire \rgf_c0bus_wb[2]_i_26_n_0 ;
  wire \rgf_c0bus_wb[2]_i_27_n_0 ;
  wire \rgf_c0bus_wb[2]_i_28_n_0 ;
  wire \rgf_c0bus_wb[2]_i_29_n_0 ;
  wire \rgf_c0bus_wb[2]_i_2_n_0 ;
  wire \rgf_c0bus_wb[2]_i_30_n_0 ;
  wire \rgf_c0bus_wb[2]_i_31_n_0 ;
  wire \rgf_c0bus_wb[2]_i_32_n_0 ;
  wire \rgf_c0bus_wb[2]_i_33_n_0 ;
  wire \rgf_c0bus_wb[2]_i_34_n_0 ;
  wire \rgf_c0bus_wb[2]_i_35_n_0 ;
  wire \rgf_c0bus_wb[2]_i_36_n_0 ;
  wire \rgf_c0bus_wb[2]_i_37_n_0 ;
  wire \rgf_c0bus_wb[2]_i_38_n_0 ;
  wire \rgf_c0bus_wb[2]_i_3_n_0 ;
  wire \rgf_c0bus_wb[2]_i_4_n_0 ;
  wire \rgf_c0bus_wb[2]_i_5_n_0 ;
  wire \rgf_c0bus_wb[2]_i_6_n_0 ;
  wire \rgf_c0bus_wb[2]_i_7_n_0 ;
  wire \rgf_c0bus_wb[2]_i_8_n_0 ;
  wire \rgf_c0bus_wb[2]_i_9_n_0 ;
  wire \rgf_c0bus_wb[30]_i_10_n_0 ;
  wire \rgf_c0bus_wb[30]_i_11_n_0 ;
  wire \rgf_c0bus_wb[30]_i_12_n_0 ;
  wire \rgf_c0bus_wb[30]_i_13_n_0 ;
  wire \rgf_c0bus_wb[30]_i_14_n_0 ;
  wire \rgf_c0bus_wb[30]_i_15_n_0 ;
  wire \rgf_c0bus_wb[30]_i_16_n_0 ;
  wire \rgf_c0bus_wb[30]_i_17_n_0 ;
  wire \rgf_c0bus_wb[30]_i_18_n_0 ;
  wire \rgf_c0bus_wb[30]_i_19_n_0 ;
  wire \rgf_c0bus_wb[30]_i_20_n_0 ;
  wire \rgf_c0bus_wb[30]_i_21_n_0 ;
  wire \rgf_c0bus_wb[30]_i_22_n_0 ;
  wire \rgf_c0bus_wb[30]_i_23_n_0 ;
  wire \rgf_c0bus_wb[30]_i_24_n_0 ;
  wire \rgf_c0bus_wb[30]_i_25_n_0 ;
  wire \rgf_c0bus_wb[30]_i_26_n_0 ;
  wire \rgf_c0bus_wb[30]_i_27_n_0 ;
  wire \rgf_c0bus_wb[30]_i_28_n_0 ;
  wire \rgf_c0bus_wb[30]_i_29_n_0 ;
  wire \rgf_c0bus_wb[30]_i_2_n_0 ;
  wire \rgf_c0bus_wb[30]_i_30_n_0 ;
  wire \rgf_c0bus_wb[30]_i_31_n_0 ;
  wire \rgf_c0bus_wb[30]_i_32_n_0 ;
  wire \rgf_c0bus_wb[30]_i_33_n_0 ;
  wire \rgf_c0bus_wb[30]_i_34_n_0 ;
  wire \rgf_c0bus_wb[30]_i_35_n_0 ;
  wire \rgf_c0bus_wb[30]_i_36_n_0 ;
  wire \rgf_c0bus_wb[30]_i_37_n_0 ;
  wire \rgf_c0bus_wb[30]_i_38_n_0 ;
  wire \rgf_c0bus_wb[30]_i_39_n_0 ;
  wire \rgf_c0bus_wb[30]_i_3_n_0 ;
  wire \rgf_c0bus_wb[30]_i_40_n_0 ;
  wire \rgf_c0bus_wb[30]_i_41_n_0 ;
  wire \rgf_c0bus_wb[30]_i_42_n_0 ;
  wire \rgf_c0bus_wb[30]_i_43_n_0 ;
  wire \rgf_c0bus_wb[30]_i_44_n_0 ;
  wire \rgf_c0bus_wb[30]_i_45_n_0 ;
  wire \rgf_c0bus_wb[30]_i_46_n_0 ;
  wire \rgf_c0bus_wb[30]_i_47_n_0 ;
  wire \rgf_c0bus_wb[30]_i_48_n_0 ;
  wire \rgf_c0bus_wb[30]_i_49_n_0 ;
  wire \rgf_c0bus_wb[30]_i_4_n_0 ;
  wire \rgf_c0bus_wb[30]_i_50_n_0 ;
  wire \rgf_c0bus_wb[30]_i_51_n_0 ;
  wire \rgf_c0bus_wb[30]_i_52_n_0 ;
  wire \rgf_c0bus_wb[30]_i_53_n_0 ;
  wire \rgf_c0bus_wb[30]_i_54_n_0 ;
  wire \rgf_c0bus_wb[30]_i_55_n_0 ;
  wire \rgf_c0bus_wb[30]_i_56_n_0 ;
  wire \rgf_c0bus_wb[30]_i_57_n_0 ;
  wire \rgf_c0bus_wb[30]_i_58_n_0 ;
  wire \rgf_c0bus_wb[30]_i_59_n_0 ;
  wire \rgf_c0bus_wb[30]_i_5_n_0 ;
  wire \rgf_c0bus_wb[30]_i_60_n_0 ;
  wire \rgf_c0bus_wb[30]_i_61_n_0 ;
  wire \rgf_c0bus_wb[30]_i_62_n_0 ;
  wire \rgf_c0bus_wb[30]_i_63_n_0 ;
  wire \rgf_c0bus_wb[30]_i_64_n_0 ;
  wire \rgf_c0bus_wb[30]_i_6_n_0 ;
  wire \rgf_c0bus_wb[30]_i_7_n_0 ;
  wire \rgf_c0bus_wb[30]_i_8_n_0 ;
  wire \rgf_c0bus_wb[30]_i_9_n_0 ;
  wire \rgf_c0bus_wb[31]_i_10_n_0 ;
  wire \rgf_c0bus_wb[31]_i_11_n_0 ;
  wire \rgf_c0bus_wb[31]_i_12_n_0 ;
  wire \rgf_c0bus_wb[31]_i_13_n_0 ;
  wire \rgf_c0bus_wb[31]_i_14_n_0 ;
  wire \rgf_c0bus_wb[31]_i_15_n_0 ;
  wire \rgf_c0bus_wb[31]_i_16_n_0 ;
  wire \rgf_c0bus_wb[31]_i_17_n_0 ;
  wire \rgf_c0bus_wb[31]_i_18_n_0 ;
  wire \rgf_c0bus_wb[31]_i_19_n_0 ;
  wire \rgf_c0bus_wb[31]_i_20_n_0 ;
  wire \rgf_c0bus_wb[31]_i_21_n_0 ;
  wire \rgf_c0bus_wb[31]_i_22_n_0 ;
  wire \rgf_c0bus_wb[31]_i_23_n_0 ;
  wire \rgf_c0bus_wb[31]_i_24_n_0 ;
  wire \rgf_c0bus_wb[31]_i_25_n_0 ;
  wire \rgf_c0bus_wb[31]_i_26_n_0 ;
  wire \rgf_c0bus_wb[31]_i_27_n_0 ;
  wire \rgf_c0bus_wb[31]_i_28_n_0 ;
  wire \rgf_c0bus_wb[31]_i_29_n_0 ;
  wire \rgf_c0bus_wb[31]_i_2_n_0 ;
  wire \rgf_c0bus_wb[31]_i_30_n_0 ;
  wire \rgf_c0bus_wb[31]_i_31_n_0 ;
  wire \rgf_c0bus_wb[31]_i_32_n_0 ;
  wire \rgf_c0bus_wb[31]_i_33_n_0 ;
  wire \rgf_c0bus_wb[31]_i_34_n_0 ;
  wire \rgf_c0bus_wb[31]_i_35_n_0 ;
  wire \rgf_c0bus_wb[31]_i_36_n_0 ;
  wire \rgf_c0bus_wb[31]_i_37_n_0 ;
  wire \rgf_c0bus_wb[31]_i_38_n_0 ;
  wire \rgf_c0bus_wb[31]_i_39_n_0 ;
  wire \rgf_c0bus_wb[31]_i_3_n_0 ;
  wire \rgf_c0bus_wb[31]_i_40_n_0 ;
  wire \rgf_c0bus_wb[31]_i_41_n_0 ;
  wire \rgf_c0bus_wb[31]_i_42_n_0 ;
  wire \rgf_c0bus_wb[31]_i_43_n_0 ;
  wire \rgf_c0bus_wb[31]_i_44_n_0 ;
  wire \rgf_c0bus_wb[31]_i_45_n_0 ;
  wire \rgf_c0bus_wb[31]_i_46_n_0 ;
  wire \rgf_c0bus_wb[31]_i_47_n_0 ;
  wire \rgf_c0bus_wb[31]_i_48_n_0 ;
  wire \rgf_c0bus_wb[31]_i_49_n_0 ;
  wire \rgf_c0bus_wb[31]_i_4_n_0 ;
  wire \rgf_c0bus_wb[31]_i_50_n_0 ;
  wire \rgf_c0bus_wb[31]_i_51_n_0 ;
  wire \rgf_c0bus_wb[31]_i_52_n_0 ;
  wire \rgf_c0bus_wb[31]_i_53_n_0 ;
  wire \rgf_c0bus_wb[31]_i_54_n_0 ;
  wire \rgf_c0bus_wb[31]_i_55_n_0 ;
  wire \rgf_c0bus_wb[31]_i_56_n_0 ;
  wire \rgf_c0bus_wb[31]_i_57_n_0 ;
  wire \rgf_c0bus_wb[31]_i_58_n_0 ;
  wire \rgf_c0bus_wb[31]_i_59_n_0 ;
  wire \rgf_c0bus_wb[31]_i_5_n_0 ;
  wire \rgf_c0bus_wb[31]_i_60_n_0 ;
  wire \rgf_c0bus_wb[31]_i_61_n_0 ;
  wire \rgf_c0bus_wb[31]_i_62_n_0 ;
  wire \rgf_c0bus_wb[31]_i_63_n_0 ;
  wire \rgf_c0bus_wb[31]_i_64_n_0 ;
  wire \rgf_c0bus_wb[31]_i_65_n_0 ;
  wire \rgf_c0bus_wb[31]_i_66_n_0 ;
  wire \rgf_c0bus_wb[31]_i_67_n_0 ;
  wire \rgf_c0bus_wb[31]_i_68_n_0 ;
  wire \rgf_c0bus_wb[31]_i_69_n_0 ;
  wire \rgf_c0bus_wb[31]_i_6_n_0 ;
  wire \rgf_c0bus_wb[31]_i_70_n_0 ;
  wire \rgf_c0bus_wb[31]_i_71_n_0 ;
  wire \rgf_c0bus_wb[31]_i_72_n_0 ;
  wire \rgf_c0bus_wb[31]_i_73_n_0 ;
  wire \rgf_c0bus_wb[31]_i_74_n_0 ;
  wire \rgf_c0bus_wb[31]_i_75_n_0 ;
  wire \rgf_c0bus_wb[31]_i_76_n_0 ;
  wire \rgf_c0bus_wb[31]_i_78_n_0 ;
  wire \rgf_c0bus_wb[31]_i_7_n_0 ;
  wire \rgf_c0bus_wb[31]_i_82_n_0 ;
  wire \rgf_c0bus_wb[31]_i_8_n_0 ;
  wire \rgf_c0bus_wb[31]_i_9_n_0 ;
  wire \rgf_c0bus_wb[3]_i_10_n_0 ;
  wire \rgf_c0bus_wb[3]_i_12_n_0 ;
  wire \rgf_c0bus_wb[3]_i_13_n_0 ;
  wire \rgf_c0bus_wb[3]_i_14_n_0 ;
  wire \rgf_c0bus_wb[3]_i_15_n_0 ;
  wire \rgf_c0bus_wb[3]_i_16_n_0 ;
  wire \rgf_c0bus_wb[3]_i_17_n_0 ;
  wire \rgf_c0bus_wb[3]_i_18_n_0 ;
  wire \rgf_c0bus_wb[3]_i_19_n_0 ;
  wire \rgf_c0bus_wb[3]_i_20_n_0 ;
  wire \rgf_c0bus_wb[3]_i_21_n_0 ;
  wire \rgf_c0bus_wb[3]_i_22_n_0 ;
  wire \rgf_c0bus_wb[3]_i_27_n_0 ;
  wire \rgf_c0bus_wb[3]_i_28_n_0 ;
  wire \rgf_c0bus_wb[3]_i_29_n_0 ;
  wire \rgf_c0bus_wb[3]_i_2_n_0 ;
  wire \rgf_c0bus_wb[3]_i_30_n_0 ;
  wire \rgf_c0bus_wb[3]_i_31_n_0 ;
  wire \rgf_c0bus_wb[3]_i_3_n_0 ;
  wire \rgf_c0bus_wb[3]_i_4_n_0 ;
  wire \rgf_c0bus_wb[3]_i_5_n_0 ;
  wire \rgf_c0bus_wb[3]_i_6_n_0 ;
  wire \rgf_c0bus_wb[3]_i_7_n_0 ;
  wire \rgf_c0bus_wb[3]_i_8_n_0 ;
  wire \rgf_c0bus_wb[3]_i_9_n_0 ;
  wire \rgf_c0bus_wb[4]_i_10_n_0 ;
  wire \rgf_c0bus_wb[4]_i_11_n_0 ;
  wire \rgf_c0bus_wb[4]_i_12_n_0 ;
  wire \rgf_c0bus_wb[4]_i_13_n_0 ;
  wire \rgf_c0bus_wb[4]_i_14_n_0 ;
  wire \rgf_c0bus_wb[4]_i_15_n_0 ;
  wire \rgf_c0bus_wb[4]_i_16_n_0 ;
  wire \rgf_c0bus_wb[4]_i_17_n_0 ;
  wire \rgf_c0bus_wb[4]_i_18_n_0 ;
  wire \rgf_c0bus_wb[4]_i_19_n_0 ;
  wire \rgf_c0bus_wb[4]_i_20_n_0 ;
  wire \rgf_c0bus_wb[4]_i_21_n_0 ;
  wire \rgf_c0bus_wb[4]_i_22_n_0 ;
  wire \rgf_c0bus_wb[4]_i_23_n_0 ;
  wire \rgf_c0bus_wb[4]_i_24_n_0 ;
  wire \rgf_c0bus_wb[4]_i_25_n_0 ;
  wire \rgf_c0bus_wb[4]_i_2_n_0 ;
  wire \rgf_c0bus_wb[4]_i_3_n_0 ;
  wire \rgf_c0bus_wb[4]_i_4_n_0 ;
  wire \rgf_c0bus_wb[4]_i_5_n_0 ;
  wire \rgf_c0bus_wb[4]_i_6_n_0 ;
  wire \rgf_c0bus_wb[4]_i_7_n_0 ;
  wire \rgf_c0bus_wb[4]_i_8_n_0 ;
  wire \rgf_c0bus_wb[4]_i_9_n_0 ;
  wire \rgf_c0bus_wb[5]_i_10_n_0 ;
  wire \rgf_c0bus_wb[5]_i_11_n_0 ;
  wire \rgf_c0bus_wb[5]_i_12_n_0 ;
  wire \rgf_c0bus_wb[5]_i_13_n_0 ;
  wire \rgf_c0bus_wb[5]_i_14_n_0 ;
  wire \rgf_c0bus_wb[5]_i_15_n_0 ;
  wire \rgf_c0bus_wb[5]_i_16_n_0 ;
  wire \rgf_c0bus_wb[5]_i_17_n_0 ;
  wire \rgf_c0bus_wb[5]_i_18_n_0 ;
  wire \rgf_c0bus_wb[5]_i_19_n_0 ;
  wire \rgf_c0bus_wb[5]_i_20_n_0 ;
  wire \rgf_c0bus_wb[5]_i_21_n_0 ;
  wire \rgf_c0bus_wb[5]_i_22_n_0 ;
  wire \rgf_c0bus_wb[5]_i_23_n_0 ;
  wire \rgf_c0bus_wb[5]_i_24_n_0 ;
  wire \rgf_c0bus_wb[5]_i_25_n_0 ;
  wire \rgf_c0bus_wb[5]_i_26_n_0 ;
  wire \rgf_c0bus_wb[5]_i_27_n_0 ;
  wire \rgf_c0bus_wb[5]_i_28_n_0 ;
  wire \rgf_c0bus_wb[5]_i_2_n_0 ;
  wire \rgf_c0bus_wb[5]_i_3_n_0 ;
  wire \rgf_c0bus_wb[5]_i_4_n_0 ;
  wire \rgf_c0bus_wb[5]_i_5_n_0 ;
  wire \rgf_c0bus_wb[5]_i_6_n_0 ;
  wire \rgf_c0bus_wb[5]_i_7_n_0 ;
  wire \rgf_c0bus_wb[5]_i_8_n_0 ;
  wire \rgf_c0bus_wb[5]_i_9_n_0 ;
  wire \rgf_c0bus_wb[6]_i_10_n_0 ;
  wire \rgf_c0bus_wb[6]_i_11_n_0 ;
  wire \rgf_c0bus_wb[6]_i_12_n_0 ;
  wire \rgf_c0bus_wb[6]_i_13_n_0 ;
  wire \rgf_c0bus_wb[6]_i_14_n_0 ;
  wire \rgf_c0bus_wb[6]_i_15_n_0 ;
  wire \rgf_c0bus_wb[6]_i_16_n_0 ;
  wire \rgf_c0bus_wb[6]_i_17_n_0 ;
  wire \rgf_c0bus_wb[6]_i_18_n_0 ;
  wire \rgf_c0bus_wb[6]_i_19_n_0 ;
  wire \rgf_c0bus_wb[6]_i_20_n_0 ;
  wire \rgf_c0bus_wb[6]_i_21_n_0 ;
  wire \rgf_c0bus_wb[6]_i_22_n_0 ;
  wire \rgf_c0bus_wb[6]_i_23_n_0 ;
  wire \rgf_c0bus_wb[6]_i_24_n_0 ;
  wire \rgf_c0bus_wb[6]_i_25_n_0 ;
  wire \rgf_c0bus_wb[6]_i_26_n_0 ;
  wire \rgf_c0bus_wb[6]_i_2_n_0 ;
  wire \rgf_c0bus_wb[6]_i_3_n_0 ;
  wire \rgf_c0bus_wb[6]_i_4_n_0 ;
  wire \rgf_c0bus_wb[6]_i_5_n_0 ;
  wire \rgf_c0bus_wb[6]_i_6_n_0 ;
  wire \rgf_c0bus_wb[6]_i_7_n_0 ;
  wire \rgf_c0bus_wb[6]_i_8_n_0 ;
  wire \rgf_c0bus_wb[6]_i_9_n_0 ;
  wire \rgf_c0bus_wb[7]_i_10_n_0 ;
  wire \rgf_c0bus_wb[7]_i_11_n_0 ;
  wire \rgf_c0bus_wb[7]_i_13_n_0 ;
  wire \rgf_c0bus_wb[7]_i_14_n_0 ;
  wire \rgf_c0bus_wb[7]_i_15_n_0 ;
  wire \rgf_c0bus_wb[7]_i_16_n_0 ;
  wire \rgf_c0bus_wb[7]_i_17_n_0 ;
  wire \rgf_c0bus_wb[7]_i_18_n_0 ;
  wire \rgf_c0bus_wb[7]_i_19_n_0 ;
  wire \rgf_c0bus_wb[7]_i_20_n_0 ;
  wire \rgf_c0bus_wb[7]_i_21_n_0 ;
  wire \rgf_c0bus_wb[7]_i_22_n_0 ;
  wire \rgf_c0bus_wb[7]_i_23_n_0 ;
  wire \rgf_c0bus_wb[7]_i_24_n_0 ;
  wire \rgf_c0bus_wb[7]_i_25_n_0 ;
  wire \rgf_c0bus_wb[7]_i_26_n_0 ;
  wire \rgf_c0bus_wb[7]_i_27_n_0 ;
  wire \rgf_c0bus_wb[7]_i_28_n_0 ;
  wire \rgf_c0bus_wb[7]_i_29_n_0 ;
  wire \rgf_c0bus_wb[7]_i_2_n_0 ;
  wire \rgf_c0bus_wb[7]_i_34_n_0 ;
  wire \rgf_c0bus_wb[7]_i_35_n_0 ;
  wire \rgf_c0bus_wb[7]_i_36_n_0 ;
  wire \rgf_c0bus_wb[7]_i_37_n_0 ;
  wire \rgf_c0bus_wb[7]_i_38_n_0 ;
  wire \rgf_c0bus_wb[7]_i_3_n_0 ;
  wire \rgf_c0bus_wb[7]_i_4_n_0 ;
  wire \rgf_c0bus_wb[7]_i_5_n_0 ;
  wire \rgf_c0bus_wb[7]_i_6_n_0 ;
  wire \rgf_c0bus_wb[7]_i_7_n_0 ;
  wire \rgf_c0bus_wb[7]_i_8_n_0 ;
  wire \rgf_c0bus_wb[7]_i_9_n_0 ;
  wire \rgf_c0bus_wb[8]_i_10_n_0 ;
  wire \rgf_c0bus_wb[8]_i_11_n_0 ;
  wire \rgf_c0bus_wb[8]_i_12_n_0 ;
  wire \rgf_c0bus_wb[8]_i_13_n_0 ;
  wire \rgf_c0bus_wb[8]_i_14_n_0 ;
  wire \rgf_c0bus_wb[8]_i_15_n_0 ;
  wire \rgf_c0bus_wb[8]_i_16_n_0 ;
  wire \rgf_c0bus_wb[8]_i_17_n_0 ;
  wire \rgf_c0bus_wb[8]_i_18_n_0 ;
  wire \rgf_c0bus_wb[8]_i_20_n_0 ;
  wire \rgf_c0bus_wb[8]_i_21_n_0 ;
  wire \rgf_c0bus_wb[8]_i_22_n_0 ;
  wire \rgf_c0bus_wb[8]_i_23_n_0 ;
  wire \rgf_c0bus_wb[8]_i_24_n_0 ;
  wire \rgf_c0bus_wb[8]_i_25_n_0 ;
  wire \rgf_c0bus_wb[8]_i_26_n_0 ;
  wire \rgf_c0bus_wb[8]_i_2_n_0 ;
  wire \rgf_c0bus_wb[8]_i_3_n_0 ;
  wire \rgf_c0bus_wb[8]_i_4_n_0 ;
  wire \rgf_c0bus_wb[8]_i_5_n_0 ;
  wire \rgf_c0bus_wb[8]_i_6_n_0 ;
  wire \rgf_c0bus_wb[8]_i_7_n_0 ;
  wire \rgf_c0bus_wb[8]_i_8_n_0 ;
  wire \rgf_c0bus_wb[8]_i_9_n_0 ;
  wire \rgf_c0bus_wb[9]_i_10_n_0 ;
  wire \rgf_c0bus_wb[9]_i_11_n_0 ;
  wire \rgf_c0bus_wb[9]_i_12_n_0 ;
  wire \rgf_c0bus_wb[9]_i_13_n_0 ;
  wire \rgf_c0bus_wb[9]_i_14_n_0 ;
  wire \rgf_c0bus_wb[9]_i_15_n_0 ;
  wire \rgf_c0bus_wb[9]_i_16_n_0 ;
  wire \rgf_c0bus_wb[9]_i_17_n_0 ;
  wire \rgf_c0bus_wb[9]_i_18_n_0 ;
  wire \rgf_c0bus_wb[9]_i_19_n_0 ;
  wire \rgf_c0bus_wb[9]_i_20_n_0 ;
  wire \rgf_c0bus_wb[9]_i_21_n_0 ;
  wire \rgf_c0bus_wb[9]_i_22_n_0 ;
  wire \rgf_c0bus_wb[9]_i_23_n_0 ;
  wire \rgf_c0bus_wb[9]_i_24_n_0 ;
  wire \rgf_c0bus_wb[9]_i_25_n_0 ;
  wire \rgf_c0bus_wb[9]_i_26_n_0 ;
  wire \rgf_c0bus_wb[9]_i_27_n_0 ;
  wire \rgf_c0bus_wb[9]_i_28_n_0 ;
  wire \rgf_c0bus_wb[9]_i_29_n_0 ;
  wire \rgf_c0bus_wb[9]_i_2_n_0 ;
  wire \rgf_c0bus_wb[9]_i_31_n_0 ;
  wire \rgf_c0bus_wb[9]_i_3_n_0 ;
  wire \rgf_c0bus_wb[9]_i_4_n_0 ;
  wire \rgf_c0bus_wb[9]_i_5_n_0 ;
  wire \rgf_c0bus_wb[9]_i_6_n_0 ;
  wire \rgf_c0bus_wb[9]_i_7_n_0 ;
  wire \rgf_c0bus_wb[9]_i_8_n_0 ;
  wire \rgf_c0bus_wb[9]_i_9_n_0 ;
  wire \rgf_c0bus_wb_reg[10]_i_19_n_0 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_0 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_1 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_2 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_3 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_4 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_5 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_6 ;
  wire \rgf_c0bus_wb_reg[11]_i_20_n_7 ;
  wire \rgf_c0bus_wb_reg[12]_i_23_n_0 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_0 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_1 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_2 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_3 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_4 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_5 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_6 ;
  wire \rgf_c0bus_wb_reg[15]_i_19_n_7 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_0 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_1 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_2 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_3 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_4 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_5 ;
  wire \rgf_c0bus_wb_reg[19]_i_11_n_7 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_0 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_1 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_2 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_3 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_4 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_5 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_6 ;
  wire \rgf_c0bus_wb_reg[23]_i_24_n_7 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_0 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_1 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_2 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_3 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_4 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_5 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_6 ;
  wire \rgf_c0bus_wb_reg[27]_i_23_n_7 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_0 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_1 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_2 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_3 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_4 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_5 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_6 ;
  wire \rgf_c0bus_wb_reg[29]_i_11_n_7 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_0 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_1 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_2 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_3 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_4 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_5 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_6 ;
  wire \rgf_c0bus_wb_reg[3]_i_11_n_7 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_0 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_1 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_2 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_3 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_4 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_5 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_6 ;
  wire \rgf_c0bus_wb_reg[7]_i_12_n_7 ;
  wire \rgf_c0bus_wb_reg[8]_i_19_n_0 ;
  wire \rgf_c1bus_wb[0]_i_10_n_0 ;
  wire \rgf_c1bus_wb[0]_i_11_n_0 ;
  wire \rgf_c1bus_wb[0]_i_12_n_0 ;
  wire \rgf_c1bus_wb[0]_i_13_n_0 ;
  wire \rgf_c1bus_wb[0]_i_14_n_0 ;
  wire \rgf_c1bus_wb[0]_i_15_n_0 ;
  wire \rgf_c1bus_wb[0]_i_16_n_0 ;
  wire \rgf_c1bus_wb[0]_i_17_n_0 ;
  wire \rgf_c1bus_wb[0]_i_18_n_0 ;
  wire \rgf_c1bus_wb[0]_i_19_n_0 ;
  wire \rgf_c1bus_wb[0]_i_20_n_0 ;
  wire \rgf_c1bus_wb[0]_i_21_n_0 ;
  wire \rgf_c1bus_wb[0]_i_2_n_0 ;
  wire \rgf_c1bus_wb[0]_i_3_n_0 ;
  wire \rgf_c1bus_wb[0]_i_4_n_0 ;
  wire \rgf_c1bus_wb[0]_i_5_n_0 ;
  wire \rgf_c1bus_wb[0]_i_6_n_0 ;
  wire \rgf_c1bus_wb[0]_i_7_n_0 ;
  wire \rgf_c1bus_wb[0]_i_8_n_0 ;
  wire \rgf_c1bus_wb[0]_i_9_n_0 ;
  wire \rgf_c1bus_wb[10]_i_10_n_0 ;
  wire \rgf_c1bus_wb[10]_i_11_n_0 ;
  wire \rgf_c1bus_wb[10]_i_12_n_0 ;
  wire \rgf_c1bus_wb[10]_i_13_n_0 ;
  wire \rgf_c1bus_wb[10]_i_14_n_0 ;
  wire \rgf_c1bus_wb[10]_i_15_n_0 ;
  wire \rgf_c1bus_wb[10]_i_16_n_0 ;
  wire \rgf_c1bus_wb[10]_i_17_n_0 ;
  wire \rgf_c1bus_wb[10]_i_18_n_0 ;
  wire \rgf_c1bus_wb[10]_i_19_n_0 ;
  wire \rgf_c1bus_wb[10]_i_20_n_0 ;
  wire \rgf_c1bus_wb[10]_i_21_n_0 ;
  wire \rgf_c1bus_wb[10]_i_22_n_0 ;
  wire \rgf_c1bus_wb[10]_i_23_n_0 ;
  wire \rgf_c1bus_wb[10]_i_24_n_0 ;
  wire \rgf_c1bus_wb[10]_i_25_n_0 ;
  wire \rgf_c1bus_wb[10]_i_26_n_0 ;
  wire \rgf_c1bus_wb[10]_i_27_n_0 ;
  wire \rgf_c1bus_wb[10]_i_28_n_0 ;
  wire \rgf_c1bus_wb[10]_i_29_n_0 ;
  wire \rgf_c1bus_wb[10]_i_2_n_0 ;
  wire \rgf_c1bus_wb[10]_i_30_n_0 ;
  wire \rgf_c1bus_wb[10]_i_31_n_0 ;
  wire \rgf_c1bus_wb[10]_i_37_n_0 ;
  wire \rgf_c1bus_wb[10]_i_38_n_0 ;
  wire \rgf_c1bus_wb[10]_i_39_n_0 ;
  wire \rgf_c1bus_wb[10]_i_3_n_0 ;
  wire \rgf_c1bus_wb[10]_i_40_n_0 ;
  wire \rgf_c1bus_wb[10]_i_4_n_0 ;
  wire \rgf_c1bus_wb[10]_i_5_n_0 ;
  wire \rgf_c1bus_wb[10]_i_6_n_0 ;
  wire \rgf_c1bus_wb[10]_i_7_n_0 ;
  wire \rgf_c1bus_wb[10]_i_8_n_0 ;
  wire \rgf_c1bus_wb[10]_i_9_n_0 ;
  wire \rgf_c1bus_wb[11]_i_11_n_0 ;
  wire \rgf_c1bus_wb[11]_i_12_n_0 ;
  wire \rgf_c1bus_wb[11]_i_13_n_0 ;
  wire \rgf_c1bus_wb[11]_i_14_n_0 ;
  wire \rgf_c1bus_wb[11]_i_15_n_0 ;
  wire \rgf_c1bus_wb[11]_i_16_n_0 ;
  wire \rgf_c1bus_wb[11]_i_17_n_0 ;
  wire \rgf_c1bus_wb[11]_i_18_n_0 ;
  wire \rgf_c1bus_wb[11]_i_19_n_0 ;
  wire \rgf_c1bus_wb[11]_i_20_n_0 ;
  wire \rgf_c1bus_wb[11]_i_21_n_0 ;
  wire \rgf_c1bus_wb[11]_i_22_n_0 ;
  wire \rgf_c1bus_wb[11]_i_23_n_0 ;
  wire \rgf_c1bus_wb[11]_i_24_n_0 ;
  wire \rgf_c1bus_wb[11]_i_25_n_0 ;
  wire \rgf_c1bus_wb[11]_i_2_n_0 ;
  wire \rgf_c1bus_wb[11]_i_30_n_0 ;
  wire \rgf_c1bus_wb[11]_i_31_n_0 ;
  wire \rgf_c1bus_wb[11]_i_32_n_0 ;
  wire \rgf_c1bus_wb[11]_i_33_n_0 ;
  wire \rgf_c1bus_wb[11]_i_34_n_0 ;
  wire \rgf_c1bus_wb[11]_i_35_n_0 ;
  wire \rgf_c1bus_wb[11]_i_36_n_0 ;
  wire \rgf_c1bus_wb[11]_i_37_n_0 ;
  wire \rgf_c1bus_wb[11]_i_3_n_0 ;
  wire \rgf_c1bus_wb[11]_i_4_n_0 ;
  wire \rgf_c1bus_wb[11]_i_5_n_0 ;
  wire \rgf_c1bus_wb[11]_i_6_n_0 ;
  wire \rgf_c1bus_wb[11]_i_7_n_0 ;
  wire \rgf_c1bus_wb[11]_i_8_n_0 ;
  wire \rgf_c1bus_wb[11]_i_9_n_0 ;
  wire \rgf_c1bus_wb[12]_i_10_n_0 ;
  wire \rgf_c1bus_wb[12]_i_11_n_0 ;
  wire \rgf_c1bus_wb[12]_i_12_n_0 ;
  wire \rgf_c1bus_wb[12]_i_13_n_0 ;
  wire \rgf_c1bus_wb[12]_i_14_n_0 ;
  wire \rgf_c1bus_wb[12]_i_15_n_0 ;
  wire \rgf_c1bus_wb[12]_i_16_n_0 ;
  wire \rgf_c1bus_wb[12]_i_17_n_0 ;
  wire \rgf_c1bus_wb[12]_i_18_n_0 ;
  wire \rgf_c1bus_wb[12]_i_19_n_0 ;
  wire \rgf_c1bus_wb[12]_i_20_n_0 ;
  wire \rgf_c1bus_wb[12]_i_21_n_0 ;
  wire \rgf_c1bus_wb[12]_i_22_n_0 ;
  wire \rgf_c1bus_wb[12]_i_23_n_0 ;
  wire \rgf_c1bus_wb[12]_i_24_n_0 ;
  wire \rgf_c1bus_wb[12]_i_25_n_0 ;
  wire \rgf_c1bus_wb[12]_i_26_n_0 ;
  wire \rgf_c1bus_wb[12]_i_27_n_0 ;
  wire \rgf_c1bus_wb[12]_i_28_n_0 ;
  wire \rgf_c1bus_wb[12]_i_29_n_0 ;
  wire \rgf_c1bus_wb[12]_i_2_n_0 ;
  wire \rgf_c1bus_wb[12]_i_30_n_0 ;
  wire \rgf_c1bus_wb[12]_i_3_n_0 ;
  wire \rgf_c1bus_wb[12]_i_4_n_0 ;
  wire \rgf_c1bus_wb[12]_i_5_n_0 ;
  wire \rgf_c1bus_wb[12]_i_6_n_0 ;
  wire \rgf_c1bus_wb[12]_i_7_n_0 ;
  wire \rgf_c1bus_wb[12]_i_8_n_0 ;
  wire \rgf_c1bus_wb[12]_i_9_n_0 ;
  wire \rgf_c1bus_wb[13]_i_10_n_0 ;
  wire \rgf_c1bus_wb[13]_i_11_n_0 ;
  wire \rgf_c1bus_wb[13]_i_12_n_0 ;
  wire \rgf_c1bus_wb[13]_i_13_n_0 ;
  wire \rgf_c1bus_wb[13]_i_14_n_0 ;
  wire \rgf_c1bus_wb[13]_i_15_n_0 ;
  wire \rgf_c1bus_wb[13]_i_16_n_0 ;
  wire \rgf_c1bus_wb[13]_i_17_n_0 ;
  wire \rgf_c1bus_wb[13]_i_18_n_0 ;
  wire \rgf_c1bus_wb[13]_i_19_n_0 ;
  wire \rgf_c1bus_wb[13]_i_20_n_0 ;
  wire \rgf_c1bus_wb[13]_i_21_n_0 ;
  wire \rgf_c1bus_wb[13]_i_22_n_0 ;
  wire \rgf_c1bus_wb[13]_i_23_n_0 ;
  wire \rgf_c1bus_wb[13]_i_24_n_0 ;
  wire \rgf_c1bus_wb[13]_i_25_n_0 ;
  wire \rgf_c1bus_wb[13]_i_26_n_0 ;
  wire \rgf_c1bus_wb[13]_i_27_n_0 ;
  wire \rgf_c1bus_wb[13]_i_28_n_0 ;
  wire \rgf_c1bus_wb[13]_i_29_n_0 ;
  wire \rgf_c1bus_wb[13]_i_2_n_0 ;
  wire \rgf_c1bus_wb[13]_i_30_n_0 ;
  wire \rgf_c1bus_wb[13]_i_31_n_0 ;
  wire \rgf_c1bus_wb[13]_i_32_n_0 ;
  wire \rgf_c1bus_wb[13]_i_33_n_0 ;
  wire \rgf_c1bus_wb[13]_i_34_n_0 ;
  wire \rgf_c1bus_wb[13]_i_35_n_0 ;
  wire \rgf_c1bus_wb[13]_i_3_n_0 ;
  wire \rgf_c1bus_wb[13]_i_4_n_0 ;
  wire \rgf_c1bus_wb[13]_i_5_n_0 ;
  wire \rgf_c1bus_wb[13]_i_6_n_0 ;
  wire \rgf_c1bus_wb[13]_i_7_n_0 ;
  wire \rgf_c1bus_wb[13]_i_8_n_0 ;
  wire \rgf_c1bus_wb[13]_i_9_n_0 ;
  wire \rgf_c1bus_wb[14]_i_10_n_0 ;
  wire \rgf_c1bus_wb[14]_i_11_n_0 ;
  wire \rgf_c1bus_wb[14]_i_12_n_0 ;
  wire \rgf_c1bus_wb[14]_i_13_n_0 ;
  wire \rgf_c1bus_wb[14]_i_14_n_0 ;
  wire \rgf_c1bus_wb[14]_i_15_n_0 ;
  wire \rgf_c1bus_wb[14]_i_16_n_0 ;
  wire \rgf_c1bus_wb[14]_i_17_n_0 ;
  wire \rgf_c1bus_wb[14]_i_18_n_0 ;
  wire \rgf_c1bus_wb[14]_i_19_n_0 ;
  wire \rgf_c1bus_wb[14]_i_20_n_0 ;
  wire \rgf_c1bus_wb[14]_i_21_n_0 ;
  wire \rgf_c1bus_wb[14]_i_22_n_0 ;
  wire \rgf_c1bus_wb[14]_i_23_n_0 ;
  wire \rgf_c1bus_wb[14]_i_24_n_0 ;
  wire \rgf_c1bus_wb[14]_i_25_n_0 ;
  wire \rgf_c1bus_wb[14]_i_26_n_0 ;
  wire \rgf_c1bus_wb[14]_i_27_n_0 ;
  wire \rgf_c1bus_wb[14]_i_28_n_0 ;
  wire \rgf_c1bus_wb[14]_i_29_n_0 ;
  wire \rgf_c1bus_wb[14]_i_2_n_0 ;
  wire \rgf_c1bus_wb[14]_i_30_n_0 ;
  wire \rgf_c1bus_wb[14]_i_31_n_0 ;
  wire \rgf_c1bus_wb[14]_i_32_n_0 ;
  wire \rgf_c1bus_wb[14]_i_33_n_0 ;
  wire \rgf_c1bus_wb[14]_i_34_n_0 ;
  wire \rgf_c1bus_wb[14]_i_3_n_0 ;
  wire \rgf_c1bus_wb[14]_i_4_n_0 ;
  wire \rgf_c1bus_wb[14]_i_5_n_0 ;
  wire \rgf_c1bus_wb[14]_i_6_n_0 ;
  wire \rgf_c1bus_wb[14]_i_7_n_0 ;
  wire \rgf_c1bus_wb[14]_i_8_n_0 ;
  wire \rgf_c1bus_wb[14]_i_9_n_0 ;
  wire \rgf_c1bus_wb[15]_i_10_n_0 ;
  wire \rgf_c1bus_wb[15]_i_11_n_0 ;
  wire \rgf_c1bus_wb[15]_i_12_n_0 ;
  wire \rgf_c1bus_wb[15]_i_13_n_0 ;
  wire \rgf_c1bus_wb[15]_i_14_n_0 ;
  wire \rgf_c1bus_wb[15]_i_15_n_0 ;
  wire \rgf_c1bus_wb[15]_i_16_n_0 ;
  wire \rgf_c1bus_wb[15]_i_17_n_0 ;
  wire \rgf_c1bus_wb[15]_i_18_n_0 ;
  wire \rgf_c1bus_wb[15]_i_19_n_0 ;
  wire \rgf_c1bus_wb[15]_i_20_n_0 ;
  wire \rgf_c1bus_wb[15]_i_21_n_0 ;
  wire \rgf_c1bus_wb[15]_i_22_n_0 ;
  wire \rgf_c1bus_wb[15]_i_23_n_0 ;
  wire \rgf_c1bus_wb[15]_i_24_n_0 ;
  wire \rgf_c1bus_wb[15]_i_25_n_0 ;
  wire \rgf_c1bus_wb[15]_i_26_n_0 ;
  wire \rgf_c1bus_wb[15]_i_27_n_0 ;
  wire \rgf_c1bus_wb[15]_i_28_n_0 ;
  wire \rgf_c1bus_wb[15]_i_29_n_0 ;
  wire \rgf_c1bus_wb[15]_i_2_n_0 ;
  wire \rgf_c1bus_wb[15]_i_30_n_0 ;
  wire \rgf_c1bus_wb[15]_i_31_n_0 ;
  wire \rgf_c1bus_wb[15]_i_32_n_0 ;
  wire \rgf_c1bus_wb[15]_i_33_n_0 ;
  wire \rgf_c1bus_wb[15]_i_3_n_0 ;
  wire \rgf_c1bus_wb[15]_i_4_n_0 ;
  wire \rgf_c1bus_wb[15]_i_5_n_0 ;
  wire \rgf_c1bus_wb[15]_i_6_n_0 ;
  wire \rgf_c1bus_wb[15]_i_7_n_0 ;
  wire \rgf_c1bus_wb[15]_i_8_n_0 ;
  wire \rgf_c1bus_wb[15]_i_9_n_0 ;
  wire \rgf_c1bus_wb[16]_i_10_n_0 ;
  wire \rgf_c1bus_wb[16]_i_11_n_0 ;
  wire \rgf_c1bus_wb[16]_i_12_n_0 ;
  wire \rgf_c1bus_wb[16]_i_13_n_0 ;
  wire \rgf_c1bus_wb[16]_i_14_n_0 ;
  wire \rgf_c1bus_wb[16]_i_15_n_0 ;
  wire \rgf_c1bus_wb[16]_i_16_n_0 ;
  wire \rgf_c1bus_wb[16]_i_17_n_0 ;
  wire \rgf_c1bus_wb[16]_i_18_n_0 ;
  wire \rgf_c1bus_wb[16]_i_19_n_0 ;
  wire \rgf_c1bus_wb[16]_i_20_n_0 ;
  wire \rgf_c1bus_wb[16]_i_21_n_0 ;
  wire \rgf_c1bus_wb[16]_i_22_n_0 ;
  wire \rgf_c1bus_wb[16]_i_23_n_0 ;
  wire \rgf_c1bus_wb[16]_i_24_n_0 ;
  wire \rgf_c1bus_wb[16]_i_25_n_0 ;
  wire \rgf_c1bus_wb[16]_i_26_n_0 ;
  wire \rgf_c1bus_wb[16]_i_27_n_0 ;
  wire \rgf_c1bus_wb[16]_i_28_n_0 ;
  wire \rgf_c1bus_wb[16]_i_29_n_0 ;
  wire \rgf_c1bus_wb[16]_i_2_n_0 ;
  wire \rgf_c1bus_wb[16]_i_30_n_0 ;
  wire \rgf_c1bus_wb[16]_i_31_n_0 ;
  wire \rgf_c1bus_wb[16]_i_32_n_0 ;
  wire \rgf_c1bus_wb[16]_i_33_n_0 ;
  wire \rgf_c1bus_wb[16]_i_34_n_0 ;
  wire \rgf_c1bus_wb[16]_i_35_n_0 ;
  wire \rgf_c1bus_wb[16]_i_36_n_0 ;
  wire \rgf_c1bus_wb[16]_i_37_n_0 ;
  wire \rgf_c1bus_wb[16]_i_38_n_0 ;
  wire \rgf_c1bus_wb[16]_i_39_n_0 ;
  wire \rgf_c1bus_wb[16]_i_3_n_0 ;
  wire \rgf_c1bus_wb[16]_i_40_n_0 ;
  wire \rgf_c1bus_wb[16]_i_41_n_0 ;
  wire \rgf_c1bus_wb[16]_i_42_n_0 ;
  wire \rgf_c1bus_wb[16]_i_43_n_0 ;
  wire \rgf_c1bus_wb[16]_i_4_n_0 ;
  wire \rgf_c1bus_wb[16]_i_5_n_0 ;
  wire \rgf_c1bus_wb[16]_i_6_n_0 ;
  wire \rgf_c1bus_wb[16]_i_7_n_0 ;
  wire \rgf_c1bus_wb[16]_i_8_n_0 ;
  wire \rgf_c1bus_wb[16]_i_9_n_0 ;
  wire \rgf_c1bus_wb[17]_i_10_n_0 ;
  wire \rgf_c1bus_wb[17]_i_11_n_0 ;
  wire \rgf_c1bus_wb[17]_i_12_n_0 ;
  wire \rgf_c1bus_wb[17]_i_13_n_0 ;
  wire \rgf_c1bus_wb[17]_i_14_n_0 ;
  wire \rgf_c1bus_wb[17]_i_15_n_0 ;
  wire \rgf_c1bus_wb[17]_i_16_n_0 ;
  wire \rgf_c1bus_wb[17]_i_17_n_0 ;
  wire \rgf_c1bus_wb[17]_i_18_n_0 ;
  wire \rgf_c1bus_wb[17]_i_19_n_0 ;
  wire \rgf_c1bus_wb[17]_i_20_n_0 ;
  wire \rgf_c1bus_wb[17]_i_21_n_0 ;
  wire \rgf_c1bus_wb[17]_i_22_n_0 ;
  wire \rgf_c1bus_wb[17]_i_23_n_0 ;
  wire \rgf_c1bus_wb[17]_i_24_n_0 ;
  wire \rgf_c1bus_wb[17]_i_25_n_0 ;
  wire \rgf_c1bus_wb[17]_i_26_n_0 ;
  wire \rgf_c1bus_wb[17]_i_27_n_0 ;
  wire \rgf_c1bus_wb[17]_i_2_n_0 ;
  wire \rgf_c1bus_wb[17]_i_3_n_0 ;
  wire \rgf_c1bus_wb[17]_i_4_n_0 ;
  wire \rgf_c1bus_wb[17]_i_5_n_0 ;
  wire \rgf_c1bus_wb[17]_i_6_n_0 ;
  wire \rgf_c1bus_wb[17]_i_7_n_0 ;
  wire \rgf_c1bus_wb[17]_i_8_n_0 ;
  wire \rgf_c1bus_wb[17]_i_9_n_0 ;
  wire \rgf_c1bus_wb[18]_i_10_n_0 ;
  wire \rgf_c1bus_wb[18]_i_11_n_0 ;
  wire \rgf_c1bus_wb[18]_i_12_n_0 ;
  wire \rgf_c1bus_wb[18]_i_13_n_0 ;
  wire \rgf_c1bus_wb[18]_i_14_n_0 ;
  wire \rgf_c1bus_wb[18]_i_15_n_0 ;
  wire \rgf_c1bus_wb[18]_i_16_n_0 ;
  wire \rgf_c1bus_wb[18]_i_17_n_0 ;
  wire \rgf_c1bus_wb[18]_i_18_n_0 ;
  wire \rgf_c1bus_wb[18]_i_19_n_0 ;
  wire \rgf_c1bus_wb[18]_i_20_n_0 ;
  wire \rgf_c1bus_wb[18]_i_21_n_0 ;
  wire \rgf_c1bus_wb[18]_i_22_n_0 ;
  wire \rgf_c1bus_wb[18]_i_23_n_0 ;
  wire \rgf_c1bus_wb[18]_i_24_n_0 ;
  wire \rgf_c1bus_wb[18]_i_25_n_0 ;
  wire \rgf_c1bus_wb[18]_i_26_n_0 ;
  wire \rgf_c1bus_wb[18]_i_27_n_0 ;
  wire \rgf_c1bus_wb[18]_i_28_n_0 ;
  wire \rgf_c1bus_wb[18]_i_29_n_0 ;
  wire \rgf_c1bus_wb[18]_i_2_n_0 ;
  wire \rgf_c1bus_wb[18]_i_3_n_0 ;
  wire \rgf_c1bus_wb[18]_i_4_n_0 ;
  wire \rgf_c1bus_wb[18]_i_5_n_0 ;
  wire \rgf_c1bus_wb[18]_i_6_n_0 ;
  wire \rgf_c1bus_wb[18]_i_7_n_0 ;
  wire \rgf_c1bus_wb[18]_i_8_n_0 ;
  wire \rgf_c1bus_wb[18]_i_9_n_0 ;
  wire \rgf_c1bus_wb[19]_i_11_n_0 ;
  wire \rgf_c1bus_wb[19]_i_12_n_0 ;
  wire \rgf_c1bus_wb[19]_i_13_n_0 ;
  wire \rgf_c1bus_wb[19]_i_14_n_0 ;
  wire \rgf_c1bus_wb[19]_i_15_n_0 ;
  wire \rgf_c1bus_wb[19]_i_16_n_0 ;
  wire \rgf_c1bus_wb[19]_i_17_n_0 ;
  wire \rgf_c1bus_wb[19]_i_19_n_0 ;
  wire \rgf_c1bus_wb[19]_i_20_n_0 ;
  wire \rgf_c1bus_wb[19]_i_21_n_0 ;
  wire \rgf_c1bus_wb[19]_i_27_n_0 ;
  wire \rgf_c1bus_wb[19]_i_28_n_0 ;
  wire \rgf_c1bus_wb[19]_i_29_n_0 ;
  wire \rgf_c1bus_wb[19]_i_2_n_0 ;
  wire \rgf_c1bus_wb[19]_i_30_n_0 ;
  wire \rgf_c1bus_wb[19]_i_31_n_0 ;
  wire \rgf_c1bus_wb[19]_i_32_n_0 ;
  wire \rgf_c1bus_wb[19]_i_33_n_0 ;
  wire \rgf_c1bus_wb[19]_i_34_n_0 ;
  wire \rgf_c1bus_wb[19]_i_3_n_0 ;
  wire \rgf_c1bus_wb[19]_i_41_n_0 ;
  wire \rgf_c1bus_wb[19]_i_42_n_0 ;
  wire \rgf_c1bus_wb[19]_i_44_n_0 ;
  wire \rgf_c1bus_wb[19]_i_45_n_0 ;
  wire \rgf_c1bus_wb[19]_i_46_n_0 ;
  wire \rgf_c1bus_wb[19]_i_4_n_0 ;
  wire \rgf_c1bus_wb[19]_i_5_n_0 ;
  wire \rgf_c1bus_wb[19]_i_6_n_0 ;
  wire \rgf_c1bus_wb[19]_i_7_n_0 ;
  wire \rgf_c1bus_wb[19]_i_8_n_0 ;
  wire \rgf_c1bus_wb[19]_i_9_n_0 ;
  wire \rgf_c1bus_wb[1]_i_10_n_0 ;
  wire \rgf_c1bus_wb[1]_i_11_n_0 ;
  wire \rgf_c1bus_wb[1]_i_12_n_0 ;
  wire \rgf_c1bus_wb[1]_i_13_n_0 ;
  wire \rgf_c1bus_wb[1]_i_14_n_0 ;
  wire \rgf_c1bus_wb[1]_i_15_n_0 ;
  wire \rgf_c1bus_wb[1]_i_16_n_0 ;
  wire \rgf_c1bus_wb[1]_i_17_n_0 ;
  wire \rgf_c1bus_wb[1]_i_18_n_0 ;
  wire \rgf_c1bus_wb[1]_i_19_n_0 ;
  wire \rgf_c1bus_wb[1]_i_20_n_0 ;
  wire \rgf_c1bus_wb[1]_i_21_n_0 ;
  wire \rgf_c1bus_wb[1]_i_22_n_0 ;
  wire \rgf_c1bus_wb[1]_i_23_n_0 ;
  wire \rgf_c1bus_wb[1]_i_24_n_0 ;
  wire \rgf_c1bus_wb[1]_i_25_n_0 ;
  wire \rgf_c1bus_wb[1]_i_2_n_0 ;
  wire \rgf_c1bus_wb[1]_i_3_n_0 ;
  wire \rgf_c1bus_wb[1]_i_4_n_0 ;
  wire \rgf_c1bus_wb[1]_i_5_n_0 ;
  wire \rgf_c1bus_wb[1]_i_6_n_0 ;
  wire \rgf_c1bus_wb[1]_i_7_n_0 ;
  wire \rgf_c1bus_wb[1]_i_8_n_0 ;
  wire \rgf_c1bus_wb[1]_i_9_n_0 ;
  wire \rgf_c1bus_wb[20]_i_10_n_0 ;
  wire \rgf_c1bus_wb[20]_i_11_n_0 ;
  wire \rgf_c1bus_wb[20]_i_12_n_0 ;
  wire \rgf_c1bus_wb[20]_i_13_n_0 ;
  wire \rgf_c1bus_wb[20]_i_14_n_0 ;
  wire \rgf_c1bus_wb[20]_i_15_n_0 ;
  wire \rgf_c1bus_wb[20]_i_16_n_0 ;
  wire \rgf_c1bus_wb[20]_i_17_n_0 ;
  wire \rgf_c1bus_wb[20]_i_18_n_0 ;
  wire \rgf_c1bus_wb[20]_i_19_n_0 ;
  wire \rgf_c1bus_wb[20]_i_20_n_0 ;
  wire \rgf_c1bus_wb[20]_i_21_n_0 ;
  wire \rgf_c1bus_wb[20]_i_22_n_0 ;
  wire \rgf_c1bus_wb[20]_i_23_n_0 ;
  wire \rgf_c1bus_wb[20]_i_24_n_0 ;
  wire \rgf_c1bus_wb[20]_i_25_n_0 ;
  wire \rgf_c1bus_wb[20]_i_26_n_0 ;
  wire \rgf_c1bus_wb[20]_i_2_n_0 ;
  wire \rgf_c1bus_wb[20]_i_3_n_0 ;
  wire \rgf_c1bus_wb[20]_i_4_n_0 ;
  wire \rgf_c1bus_wb[20]_i_5_n_0 ;
  wire \rgf_c1bus_wb[20]_i_6_n_0 ;
  wire \rgf_c1bus_wb[20]_i_7_n_0 ;
  wire \rgf_c1bus_wb[20]_i_8_n_0 ;
  wire \rgf_c1bus_wb[20]_i_9_n_0 ;
  wire \rgf_c1bus_wb[21]_i_10_n_0 ;
  wire \rgf_c1bus_wb[21]_i_11_n_0 ;
  wire \rgf_c1bus_wb[21]_i_12_n_0 ;
  wire \rgf_c1bus_wb[21]_i_13_n_0 ;
  wire \rgf_c1bus_wb[21]_i_14_n_0 ;
  wire \rgf_c1bus_wb[21]_i_15_n_0 ;
  wire \rgf_c1bus_wb[21]_i_16_n_0 ;
  wire \rgf_c1bus_wb[21]_i_17_n_0 ;
  wire \rgf_c1bus_wb[21]_i_18_n_0 ;
  wire \rgf_c1bus_wb[21]_i_19_n_0 ;
  wire \rgf_c1bus_wb[21]_i_20_n_0 ;
  wire \rgf_c1bus_wb[21]_i_21_n_0 ;
  wire \rgf_c1bus_wb[21]_i_22_n_0 ;
  wire \rgf_c1bus_wb[21]_i_23_n_0 ;
  wire \rgf_c1bus_wb[21]_i_24_n_0 ;
  wire \rgf_c1bus_wb[21]_i_25_n_0 ;
  wire \rgf_c1bus_wb[21]_i_26_n_0 ;
  wire \rgf_c1bus_wb[21]_i_27_n_0 ;
  wire \rgf_c1bus_wb[21]_i_28_n_0 ;
  wire \rgf_c1bus_wb[21]_i_2_n_0 ;
  wire \rgf_c1bus_wb[21]_i_3_n_0 ;
  wire \rgf_c1bus_wb[21]_i_4_n_0 ;
  wire \rgf_c1bus_wb[21]_i_5_n_0 ;
  wire \rgf_c1bus_wb[21]_i_6_n_0 ;
  wire \rgf_c1bus_wb[21]_i_7_n_0 ;
  wire \rgf_c1bus_wb[21]_i_8_n_0 ;
  wire \rgf_c1bus_wb[21]_i_9_n_0 ;
  wire \rgf_c1bus_wb[22]_i_10_n_0 ;
  wire \rgf_c1bus_wb[22]_i_11_n_0 ;
  wire \rgf_c1bus_wb[22]_i_12_n_0 ;
  wire \rgf_c1bus_wb[22]_i_13_n_0 ;
  wire \rgf_c1bus_wb[22]_i_14_n_0 ;
  wire \rgf_c1bus_wb[22]_i_15_n_0 ;
  wire \rgf_c1bus_wb[22]_i_16_n_0 ;
  wire \rgf_c1bus_wb[22]_i_17_n_0 ;
  wire \rgf_c1bus_wb[22]_i_18_n_0 ;
  wire \rgf_c1bus_wb[22]_i_19_n_0 ;
  wire \rgf_c1bus_wb[22]_i_20_n_0 ;
  wire \rgf_c1bus_wb[22]_i_21_n_0 ;
  wire \rgf_c1bus_wb[22]_i_22_n_0 ;
  wire \rgf_c1bus_wb[22]_i_23_n_0 ;
  wire \rgf_c1bus_wb[22]_i_2_n_0 ;
  wire \rgf_c1bus_wb[22]_i_3_n_0 ;
  wire \rgf_c1bus_wb[22]_i_4_n_0 ;
  wire \rgf_c1bus_wb[22]_i_5_n_0 ;
  wire \rgf_c1bus_wb[22]_i_6_n_0 ;
  wire \rgf_c1bus_wb[22]_i_7_n_0 ;
  wire \rgf_c1bus_wb[22]_i_8_n_0 ;
  wire \rgf_c1bus_wb[22]_i_9_n_0 ;
  wire \rgf_c1bus_wb[23]_i_10_n_0 ;
  wire \rgf_c1bus_wb[23]_i_12_n_0 ;
  wire \rgf_c1bus_wb[23]_i_13_n_0 ;
  wire \rgf_c1bus_wb[23]_i_14_n_0 ;
  wire \rgf_c1bus_wb[23]_i_15_n_0 ;
  wire \rgf_c1bus_wb[23]_i_16_n_0 ;
  wire \rgf_c1bus_wb[23]_i_17_n_0 ;
  wire \rgf_c1bus_wb[23]_i_18_n_0 ;
  wire \rgf_c1bus_wb[23]_i_19_n_0 ;
  wire \rgf_c1bus_wb[23]_i_20_n_0 ;
  wire \rgf_c1bus_wb[23]_i_21_n_0 ;
  wire \rgf_c1bus_wb[23]_i_22_n_0 ;
  wire \rgf_c1bus_wb[23]_i_23_n_0 ;
  wire \rgf_c1bus_wb[23]_i_24_n_0 ;
  wire \rgf_c1bus_wb[23]_i_25_n_0 ;
  wire \rgf_c1bus_wb[23]_i_26_n_0 ;
  wire \rgf_c1bus_wb[23]_i_2_n_0 ;
  wire \rgf_c1bus_wb[23]_i_30_n_0 ;
  wire \rgf_c1bus_wb[23]_i_31_n_0 ;
  wire \rgf_c1bus_wb[23]_i_32_n_0 ;
  wire \rgf_c1bus_wb[23]_i_33_n_0 ;
  wire \rgf_c1bus_wb[23]_i_34_n_0 ;
  wire \rgf_c1bus_wb[23]_i_35_n_0 ;
  wire \rgf_c1bus_wb[23]_i_36_n_0 ;
  wire \rgf_c1bus_wb[23]_i_37_n_0 ;
  wire \rgf_c1bus_wb[23]_i_38_n_0 ;
  wire \rgf_c1bus_wb[23]_i_39_n_0 ;
  wire \rgf_c1bus_wb[23]_i_3_n_0 ;
  wire \rgf_c1bus_wb[23]_i_40_n_0 ;
  wire \rgf_c1bus_wb[23]_i_41_n_0 ;
  wire \rgf_c1bus_wb[23]_i_42_n_0 ;
  wire \rgf_c1bus_wb[23]_i_4_n_0 ;
  wire \rgf_c1bus_wb[23]_i_5_n_0 ;
  wire \rgf_c1bus_wb[23]_i_6_n_0 ;
  wire \rgf_c1bus_wb[23]_i_7_n_0 ;
  wire \rgf_c1bus_wb[23]_i_8_n_0 ;
  wire \rgf_c1bus_wb[23]_i_9_n_0 ;
  wire \rgf_c1bus_wb[24]_i_10_n_0 ;
  wire \rgf_c1bus_wb[24]_i_11_n_0 ;
  wire \rgf_c1bus_wb[24]_i_12_n_0 ;
  wire \rgf_c1bus_wb[24]_i_13_n_0 ;
  wire \rgf_c1bus_wb[24]_i_14_n_0 ;
  wire \rgf_c1bus_wb[24]_i_15_n_0 ;
  wire \rgf_c1bus_wb[24]_i_16_n_0 ;
  wire \rgf_c1bus_wb[24]_i_17_n_0 ;
  wire \rgf_c1bus_wb[24]_i_18_n_0 ;
  wire \rgf_c1bus_wb[24]_i_19_n_0 ;
  wire \rgf_c1bus_wb[24]_i_20_n_0 ;
  wire \rgf_c1bus_wb[24]_i_21_n_0 ;
  wire \rgf_c1bus_wb[24]_i_22_n_0 ;
  wire \rgf_c1bus_wb[24]_i_23_n_0 ;
  wire \rgf_c1bus_wb[24]_i_24_n_0 ;
  wire \rgf_c1bus_wb[24]_i_25_n_0 ;
  wire \rgf_c1bus_wb[24]_i_26_n_0 ;
  wire \rgf_c1bus_wb[24]_i_27_n_0 ;
  wire \rgf_c1bus_wb[24]_i_28_n_0 ;
  wire \rgf_c1bus_wb[24]_i_29_n_0 ;
  wire \rgf_c1bus_wb[24]_i_30_n_0 ;
  wire \rgf_c1bus_wb[24]_i_31_n_0 ;
  wire \rgf_c1bus_wb[24]_i_32_n_0 ;
  wire \rgf_c1bus_wb[24]_i_33_n_0 ;
  wire \rgf_c1bus_wb[24]_i_34_n_0 ;
  wire \rgf_c1bus_wb[24]_i_3_n_0 ;
  wire \rgf_c1bus_wb[24]_i_4_n_0 ;
  wire \rgf_c1bus_wb[24]_i_7_n_0 ;
  wire \rgf_c1bus_wb[24]_i_8_n_0 ;
  wire \rgf_c1bus_wb[24]_i_9_n_0 ;
  wire \rgf_c1bus_wb[25]_i_10_n_0 ;
  wire \rgf_c1bus_wb[25]_i_11_n_0 ;
  wire \rgf_c1bus_wb[25]_i_12_n_0 ;
  wire \rgf_c1bus_wb[25]_i_13_n_0 ;
  wire \rgf_c1bus_wb[25]_i_14_n_0 ;
  wire \rgf_c1bus_wb[25]_i_15_n_0 ;
  wire \rgf_c1bus_wb[25]_i_16_n_0 ;
  wire \rgf_c1bus_wb[25]_i_17_n_0 ;
  wire \rgf_c1bus_wb[25]_i_18_n_0 ;
  wire \rgf_c1bus_wb[25]_i_19_n_0 ;
  wire \rgf_c1bus_wb[25]_i_20_n_0 ;
  wire \rgf_c1bus_wb[25]_i_21_n_0 ;
  wire \rgf_c1bus_wb[25]_i_22_n_0 ;
  wire \rgf_c1bus_wb[25]_i_23_n_0 ;
  wire \rgf_c1bus_wb[25]_i_24_n_0 ;
  wire \rgf_c1bus_wb[25]_i_25_n_0 ;
  wire \rgf_c1bus_wb[25]_i_26_n_0 ;
  wire \rgf_c1bus_wb[25]_i_27_n_0 ;
  wire \rgf_c1bus_wb[25]_i_28_n_0 ;
  wire \rgf_c1bus_wb[25]_i_29_n_0 ;
  wire \rgf_c1bus_wb[25]_i_2_n_0 ;
  wire \rgf_c1bus_wb[25]_i_30_n_0 ;
  wire \rgf_c1bus_wb[25]_i_3_n_0 ;
  wire \rgf_c1bus_wb[25]_i_4_n_0 ;
  wire \rgf_c1bus_wb[25]_i_5_n_0 ;
  wire \rgf_c1bus_wb[25]_i_6_n_0 ;
  wire \rgf_c1bus_wb[25]_i_7_n_0 ;
  wire \rgf_c1bus_wb[25]_i_8_n_0 ;
  wire \rgf_c1bus_wb[25]_i_9_n_0 ;
  wire \rgf_c1bus_wb[26]_i_10_n_0 ;
  wire \rgf_c1bus_wb[26]_i_11_n_0 ;
  wire \rgf_c1bus_wb[26]_i_12_n_0 ;
  wire \rgf_c1bus_wb[26]_i_13_n_0 ;
  wire \rgf_c1bus_wb[26]_i_14_n_0 ;
  wire \rgf_c1bus_wb[26]_i_15_n_0 ;
  wire \rgf_c1bus_wb[26]_i_16_n_0 ;
  wire \rgf_c1bus_wb[26]_i_17_n_0 ;
  wire \rgf_c1bus_wb[26]_i_18_n_0 ;
  wire \rgf_c1bus_wb[26]_i_19_n_0 ;
  wire \rgf_c1bus_wb[26]_i_20_n_0 ;
  wire \rgf_c1bus_wb[26]_i_21_n_0 ;
  wire \rgf_c1bus_wb[26]_i_22_n_0 ;
  wire \rgf_c1bus_wb[26]_i_23_n_0 ;
  wire \rgf_c1bus_wb[26]_i_24_n_0 ;
  wire \rgf_c1bus_wb[26]_i_25_n_0 ;
  wire \rgf_c1bus_wb[26]_i_26_n_0 ;
  wire \rgf_c1bus_wb[26]_i_27_n_0 ;
  wire \rgf_c1bus_wb[26]_i_28_n_0 ;
  wire \rgf_c1bus_wb[26]_i_29_n_0 ;
  wire \rgf_c1bus_wb[26]_i_30_n_0 ;
  wire \rgf_c1bus_wb[26]_i_31_n_0 ;
  wire \rgf_c1bus_wb[26]_i_32_n_0 ;
  wire \rgf_c1bus_wb[26]_i_3_n_0 ;
  wire \rgf_c1bus_wb[26]_i_4_n_0 ;
  wire \rgf_c1bus_wb[26]_i_7_n_0 ;
  wire \rgf_c1bus_wb[26]_i_8_n_0 ;
  wire \rgf_c1bus_wb[26]_i_9_n_0 ;
  wire \rgf_c1bus_wb[27]_i_11_n_0 ;
  wire \rgf_c1bus_wb[27]_i_12_n_0 ;
  wire \rgf_c1bus_wb[27]_i_13_n_0 ;
  wire \rgf_c1bus_wb[27]_i_14_n_0 ;
  wire \rgf_c1bus_wb[27]_i_15_n_0 ;
  wire \rgf_c1bus_wb[27]_i_16_n_0 ;
  wire \rgf_c1bus_wb[27]_i_17_n_0 ;
  wire \rgf_c1bus_wb[27]_i_18_n_0 ;
  wire \rgf_c1bus_wb[27]_i_19_n_0 ;
  wire \rgf_c1bus_wb[27]_i_20_n_0 ;
  wire \rgf_c1bus_wb[27]_i_25_n_0 ;
  wire \rgf_c1bus_wb[27]_i_26_n_0 ;
  wire \rgf_c1bus_wb[27]_i_27_n_0 ;
  wire \rgf_c1bus_wb[27]_i_28_n_0 ;
  wire \rgf_c1bus_wb[27]_i_29_n_0 ;
  wire \rgf_c1bus_wb[27]_i_2_n_0 ;
  wire \rgf_c1bus_wb[27]_i_30_n_0 ;
  wire \rgf_c1bus_wb[27]_i_31_n_0 ;
  wire \rgf_c1bus_wb[27]_i_32_n_0 ;
  wire \rgf_c1bus_wb[27]_i_33_n_0 ;
  wire \rgf_c1bus_wb[27]_i_34_n_0 ;
  wire \rgf_c1bus_wb[27]_i_35_n_0 ;
  wire \rgf_c1bus_wb[27]_i_36_n_0 ;
  wire \rgf_c1bus_wb[27]_i_37_n_0 ;
  wire \rgf_c1bus_wb[27]_i_38_n_0 ;
  wire \rgf_c1bus_wb[27]_i_39_n_0 ;
  wire \rgf_c1bus_wb[27]_i_3_n_0 ;
  wire \rgf_c1bus_wb[27]_i_40_n_0 ;
  wire \rgf_c1bus_wb[27]_i_41_n_0 ;
  wire \rgf_c1bus_wb[27]_i_42_n_0 ;
  wire \rgf_c1bus_wb[27]_i_43_n_0 ;
  wire \rgf_c1bus_wb[27]_i_44_n_0 ;
  wire \rgf_c1bus_wb[27]_i_45_n_0 ;
  wire \rgf_c1bus_wb[27]_i_46_n_0 ;
  wire \rgf_c1bus_wb[27]_i_4_n_0 ;
  wire \rgf_c1bus_wb[27]_i_5_n_0 ;
  wire \rgf_c1bus_wb[27]_i_6_n_0 ;
  wire \rgf_c1bus_wb[27]_i_7_n_0 ;
  wire \rgf_c1bus_wb[27]_i_8_n_0 ;
  wire \rgf_c1bus_wb[27]_i_9_n_0 ;
  wire \rgf_c1bus_wb[28]_i_10_n_0 ;
  wire \rgf_c1bus_wb[28]_i_11_n_0 ;
  wire \rgf_c1bus_wb[28]_i_12_n_0 ;
  wire \rgf_c1bus_wb[28]_i_13_n_0 ;
  wire \rgf_c1bus_wb[28]_i_14_n_0 ;
  wire \rgf_c1bus_wb[28]_i_15_n_0 ;
  wire \rgf_c1bus_wb[28]_i_16_n_0 ;
  wire \rgf_c1bus_wb[28]_i_17_n_0 ;
  wire \rgf_c1bus_wb[28]_i_18_n_0 ;
  wire \rgf_c1bus_wb[28]_i_19_n_0 ;
  wire \rgf_c1bus_wb[28]_i_20_n_0 ;
  wire \rgf_c1bus_wb[28]_i_21_n_0 ;
  wire \rgf_c1bus_wb[28]_i_22_n_0 ;
  wire \rgf_c1bus_wb[28]_i_23_n_0 ;
  wire \rgf_c1bus_wb[28]_i_24_n_0 ;
  wire \rgf_c1bus_wb[28]_i_25_n_0 ;
  wire \rgf_c1bus_wb[28]_i_26_n_0 ;
  wire \rgf_c1bus_wb[28]_i_27_n_0 ;
  wire \rgf_c1bus_wb[28]_i_28_n_0 ;
  wire \rgf_c1bus_wb[28]_i_29_n_0 ;
  wire \rgf_c1bus_wb[28]_i_2_n_0 ;
  wire \rgf_c1bus_wb[28]_i_30_n_0 ;
  wire \rgf_c1bus_wb[28]_i_31_n_0 ;
  wire \rgf_c1bus_wb[28]_i_32_n_0 ;
  wire \rgf_c1bus_wb[28]_i_33_n_0 ;
  wire \rgf_c1bus_wb[28]_i_34_n_0 ;
  wire \rgf_c1bus_wb[28]_i_35_n_0 ;
  wire \rgf_c1bus_wb[28]_i_36_n_0 ;
  wire \rgf_c1bus_wb[28]_i_37_n_0 ;
  wire \rgf_c1bus_wb[28]_i_38_n_0 ;
  wire \rgf_c1bus_wb[28]_i_39_n_0 ;
  wire \rgf_c1bus_wb[28]_i_3_n_0 ;
  wire \rgf_c1bus_wb[28]_i_40_n_0 ;
  wire \rgf_c1bus_wb[28]_i_41_n_0 ;
  wire \rgf_c1bus_wb[28]_i_42_n_0 ;
  wire \rgf_c1bus_wb[28]_i_4_n_0 ;
  wire \rgf_c1bus_wb[28]_i_5_n_0 ;
  wire \rgf_c1bus_wb[28]_i_69_n_0 ;
  wire \rgf_c1bus_wb[28]_i_6_n_0 ;
  wire \rgf_c1bus_wb[28]_i_70_n_0 ;
  wire \rgf_c1bus_wb[28]_i_71_n_0 ;
  wire \rgf_c1bus_wb[28]_i_72_n_0 ;
  wire \rgf_c1bus_wb[28]_i_73_n_0 ;
  wire \rgf_c1bus_wb[28]_i_74_n_0 ;
  wire \rgf_c1bus_wb[28]_i_75_n_0 ;
  wire \rgf_c1bus_wb[28]_i_76_n_0 ;
  wire \rgf_c1bus_wb[28]_i_77_n_0 ;
  wire \rgf_c1bus_wb[28]_i_78_n_0 ;
  wire \rgf_c1bus_wb[28]_i_79_n_0 ;
  wire \rgf_c1bus_wb[28]_i_7_n_0 ;
  wire \rgf_c1bus_wb[28]_i_80_n_0 ;
  wire \rgf_c1bus_wb[28]_i_81_n_0 ;
  wire \rgf_c1bus_wb[28]_i_82_n_0 ;
  wire \rgf_c1bus_wb[28]_i_83_n_0 ;
  wire \rgf_c1bus_wb[28]_i_84_n_0 ;
  wire \rgf_c1bus_wb[28]_i_85_n_0 ;
  wire \rgf_c1bus_wb[28]_i_86_n_0 ;
  wire \rgf_c1bus_wb[28]_i_87_n_0 ;
  wire \rgf_c1bus_wb[28]_i_88_n_0 ;
  wire \rgf_c1bus_wb[28]_i_89_n_0 ;
  wire \rgf_c1bus_wb[28]_i_8_n_0 ;
  wire \rgf_c1bus_wb[28]_i_90_n_0 ;
  wire \rgf_c1bus_wb[28]_i_91_n_0 ;
  wire \rgf_c1bus_wb[28]_i_92_n_0 ;
  wire \rgf_c1bus_wb[28]_i_9_n_0 ;
  wire \rgf_c1bus_wb[29]_i_10_n_0 ;
  wire \rgf_c1bus_wb[29]_i_11_n_0 ;
  wire \rgf_c1bus_wb[29]_i_12_n_0 ;
  wire \rgf_c1bus_wb[29]_i_13_n_0 ;
  wire \rgf_c1bus_wb[29]_i_14_n_0 ;
  wire \rgf_c1bus_wb[29]_i_15_n_0 ;
  wire \rgf_c1bus_wb[29]_i_16_n_0 ;
  wire \rgf_c1bus_wb[29]_i_17_n_0 ;
  wire \rgf_c1bus_wb[29]_i_18_n_0 ;
  wire \rgf_c1bus_wb[29]_i_19_n_0 ;
  wire \rgf_c1bus_wb[29]_i_20_n_0 ;
  wire \rgf_c1bus_wb[29]_i_21_n_0 ;
  wire \rgf_c1bus_wb[29]_i_22_n_0 ;
  wire \rgf_c1bus_wb[29]_i_23_n_0 ;
  wire \rgf_c1bus_wb[29]_i_24_n_0 ;
  wire \rgf_c1bus_wb[29]_i_25_n_0 ;
  wire \rgf_c1bus_wb[29]_i_26_n_0 ;
  wire \rgf_c1bus_wb[29]_i_27_n_0 ;
  wire \rgf_c1bus_wb[29]_i_28_n_0 ;
  wire \rgf_c1bus_wb[29]_i_29_n_0 ;
  wire \rgf_c1bus_wb[29]_i_2_n_0 ;
  wire \rgf_c1bus_wb[29]_i_30_n_0 ;
  wire \rgf_c1bus_wb[29]_i_31_n_0 ;
  wire \rgf_c1bus_wb[29]_i_32_n_0 ;
  wire \rgf_c1bus_wb[29]_i_33_n_0 ;
  wire \rgf_c1bus_wb[29]_i_34_n_0 ;
  wire \rgf_c1bus_wb[29]_i_35_n_0 ;
  wire \rgf_c1bus_wb[29]_i_36_n_0 ;
  wire \rgf_c1bus_wb[29]_i_37_n_0 ;
  wire \rgf_c1bus_wb[29]_i_38_n_0 ;
  wire \rgf_c1bus_wb[29]_i_39_n_0 ;
  wire \rgf_c1bus_wb[29]_i_3_n_0 ;
  wire \rgf_c1bus_wb[29]_i_40_n_0 ;
  wire \rgf_c1bus_wb[29]_i_41_n_0 ;
  wire \rgf_c1bus_wb[29]_i_42_n_0 ;
  wire \rgf_c1bus_wb[29]_i_43_n_0 ;
  wire \rgf_c1bus_wb[29]_i_44_n_0 ;
  wire \rgf_c1bus_wb[29]_i_45_n_0 ;
  wire \rgf_c1bus_wb[29]_i_46_n_0 ;
  wire \rgf_c1bus_wb[29]_i_4_n_0 ;
  wire \rgf_c1bus_wb[29]_i_5_n_0 ;
  wire \rgf_c1bus_wb[29]_i_6_n_0 ;
  wire \rgf_c1bus_wb[29]_i_7_n_0 ;
  wire \rgf_c1bus_wb[29]_i_8_n_0 ;
  wire \rgf_c1bus_wb[29]_i_9_n_0 ;
  wire \rgf_c1bus_wb[2]_i_10_n_0 ;
  wire \rgf_c1bus_wb[2]_i_11_n_0 ;
  wire \rgf_c1bus_wb[2]_i_12_n_0 ;
  wire \rgf_c1bus_wb[2]_i_13_n_0 ;
  wire \rgf_c1bus_wb[2]_i_14_n_0 ;
  wire \rgf_c1bus_wb[2]_i_15_n_0 ;
  wire \rgf_c1bus_wb[2]_i_16_n_0 ;
  wire \rgf_c1bus_wb[2]_i_17_n_0 ;
  wire \rgf_c1bus_wb[2]_i_18_n_0 ;
  wire \rgf_c1bus_wb[2]_i_19_n_0 ;
  wire \rgf_c1bus_wb[2]_i_20_n_0 ;
  wire \rgf_c1bus_wb[2]_i_21_n_0 ;
  wire \rgf_c1bus_wb[2]_i_22_n_0 ;
  wire \rgf_c1bus_wb[2]_i_23_n_0 ;
  wire \rgf_c1bus_wb[2]_i_24_n_0 ;
  wire \rgf_c1bus_wb[2]_i_25_n_0 ;
  wire \rgf_c1bus_wb[2]_i_2_n_0 ;
  wire \rgf_c1bus_wb[2]_i_3_n_0 ;
  wire \rgf_c1bus_wb[2]_i_4_n_0 ;
  wire \rgf_c1bus_wb[2]_i_5_n_0 ;
  wire \rgf_c1bus_wb[2]_i_6_n_0 ;
  wire \rgf_c1bus_wb[2]_i_7_n_0 ;
  wire \rgf_c1bus_wb[2]_i_8_n_0 ;
  wire \rgf_c1bus_wb[2]_i_9_n_0 ;
  wire \rgf_c1bus_wb[30]_i_10_n_0 ;
  wire \rgf_c1bus_wb[30]_i_11_n_0 ;
  wire \rgf_c1bus_wb[30]_i_12_n_0 ;
  wire \rgf_c1bus_wb[30]_i_13_n_0 ;
  wire \rgf_c1bus_wb[30]_i_14_n_0 ;
  wire \rgf_c1bus_wb[30]_i_15_n_0 ;
  wire \rgf_c1bus_wb[30]_i_16_n_0 ;
  wire \rgf_c1bus_wb[30]_i_17_n_0 ;
  wire \rgf_c1bus_wb[30]_i_18_n_0 ;
  wire \rgf_c1bus_wb[30]_i_19_n_0 ;
  wire \rgf_c1bus_wb[30]_i_20_n_0 ;
  wire \rgf_c1bus_wb[30]_i_21_n_0 ;
  wire \rgf_c1bus_wb[30]_i_22_n_0 ;
  wire \rgf_c1bus_wb[30]_i_23_n_0 ;
  wire \rgf_c1bus_wb[30]_i_24_n_0 ;
  wire \rgf_c1bus_wb[30]_i_25_n_0 ;
  wire \rgf_c1bus_wb[30]_i_26_n_0 ;
  wire \rgf_c1bus_wb[30]_i_27_n_0 ;
  wire \rgf_c1bus_wb[30]_i_28_n_0 ;
  wire \rgf_c1bus_wb[30]_i_29_n_0 ;
  wire \rgf_c1bus_wb[30]_i_30_n_0 ;
  wire \rgf_c1bus_wb[30]_i_31_n_0 ;
  wire \rgf_c1bus_wb[30]_i_32_n_0 ;
  wire \rgf_c1bus_wb[30]_i_33_n_0 ;
  wire \rgf_c1bus_wb[30]_i_34_n_0 ;
  wire \rgf_c1bus_wb[30]_i_35_n_0 ;
  wire \rgf_c1bus_wb[30]_i_36_n_0 ;
  wire \rgf_c1bus_wb[30]_i_37_n_0 ;
  wire \rgf_c1bus_wb[30]_i_38_n_0 ;
  wire \rgf_c1bus_wb[30]_i_39_n_0 ;
  wire \rgf_c1bus_wb[30]_i_3_n_0 ;
  wire \rgf_c1bus_wb[30]_i_40_n_0 ;
  wire \rgf_c1bus_wb[30]_i_41_n_0 ;
  wire \rgf_c1bus_wb[30]_i_42_n_0 ;
  wire \rgf_c1bus_wb[30]_i_43_n_0 ;
  wire \rgf_c1bus_wb[30]_i_44_n_0 ;
  wire \rgf_c1bus_wb[30]_i_45_n_0 ;
  wire \rgf_c1bus_wb[30]_i_46_n_0 ;
  wire \rgf_c1bus_wb[30]_i_47_n_0 ;
  wire \rgf_c1bus_wb[30]_i_48_n_0 ;
  wire \rgf_c1bus_wb[30]_i_49_n_0 ;
  wire \rgf_c1bus_wb[30]_i_4_n_0 ;
  wire \rgf_c1bus_wb[30]_i_50_n_0 ;
  wire \rgf_c1bus_wb[30]_i_51_n_0 ;
  wire \rgf_c1bus_wb[30]_i_52_n_0 ;
  wire \rgf_c1bus_wb[30]_i_53_n_0 ;
  wire \rgf_c1bus_wb[30]_i_7_n_0 ;
  wire \rgf_c1bus_wb[30]_i_8_n_0 ;
  wire \rgf_c1bus_wb[30]_i_9_n_0 ;
  wire \rgf_c1bus_wb[31]_i_10_n_0 ;
  wire \rgf_c1bus_wb[31]_i_12_n_0 ;
  wire \rgf_c1bus_wb[31]_i_13_n_0 ;
  wire \rgf_c1bus_wb[31]_i_14_n_0 ;
  wire \rgf_c1bus_wb[31]_i_15_n_0 ;
  wire \rgf_c1bus_wb[31]_i_16_n_0 ;
  wire \rgf_c1bus_wb[31]_i_17_n_0 ;
  wire \rgf_c1bus_wb[31]_i_18_n_0 ;
  wire \rgf_c1bus_wb[31]_i_19_n_0 ;
  wire \rgf_c1bus_wb[31]_i_20_n_0 ;
  wire \rgf_c1bus_wb[31]_i_21_n_0 ;
  wire \rgf_c1bus_wb[31]_i_22_n_0 ;
  wire \rgf_c1bus_wb[31]_i_23_n_0 ;
  wire \rgf_c1bus_wb[31]_i_24_n_0 ;
  wire \rgf_c1bus_wb[31]_i_25_n_0 ;
  wire \rgf_c1bus_wb[31]_i_26_n_0 ;
  wire \rgf_c1bus_wb[31]_i_27_n_0 ;
  wire \rgf_c1bus_wb[31]_i_28_n_0 ;
  wire \rgf_c1bus_wb[31]_i_33_n_0 ;
  wire \rgf_c1bus_wb[31]_i_34_n_0 ;
  wire \rgf_c1bus_wb[31]_i_35_n_0 ;
  wire \rgf_c1bus_wb[31]_i_36_n_0 ;
  wire \rgf_c1bus_wb[31]_i_37_n_0 ;
  wire \rgf_c1bus_wb[31]_i_38_n_0 ;
  wire \rgf_c1bus_wb[31]_i_39_n_0 ;
  wire \rgf_c1bus_wb[31]_i_3_n_0 ;
  wire \rgf_c1bus_wb[31]_i_40_n_0 ;
  wire \rgf_c1bus_wb[31]_i_41_n_0 ;
  wire \rgf_c1bus_wb[31]_i_42_n_0 ;
  wire \rgf_c1bus_wb[31]_i_43_n_0 ;
  wire \rgf_c1bus_wb[31]_i_44_n_0 ;
  wire \rgf_c1bus_wb[31]_i_45_n_0 ;
  wire \rgf_c1bus_wb[31]_i_46_n_0 ;
  wire \rgf_c1bus_wb[31]_i_47_n_0 ;
  wire \rgf_c1bus_wb[31]_i_48_n_0 ;
  wire \rgf_c1bus_wb[31]_i_49_n_0 ;
  wire \rgf_c1bus_wb[31]_i_4_n_0 ;
  wire \rgf_c1bus_wb[31]_i_50_n_0 ;
  wire \rgf_c1bus_wb[31]_i_51_n_0 ;
  wire \rgf_c1bus_wb[31]_i_52_n_0 ;
  wire \rgf_c1bus_wb[31]_i_53_n_0 ;
  wire \rgf_c1bus_wb[31]_i_54_n_0 ;
  wire \rgf_c1bus_wb[31]_i_55_n_0 ;
  wire \rgf_c1bus_wb[31]_i_56_n_0 ;
  wire \rgf_c1bus_wb[31]_i_57_n_0 ;
  wire \rgf_c1bus_wb[31]_i_58_n_0 ;
  wire \rgf_c1bus_wb[31]_i_59_n_0 ;
  wire \rgf_c1bus_wb[31]_i_5_n_0 ;
  wire \rgf_c1bus_wb[31]_i_60_n_0 ;
  wire \rgf_c1bus_wb[31]_i_61_n_0 ;
  wire \rgf_c1bus_wb[31]_i_62_n_0 ;
  wire \rgf_c1bus_wb[31]_i_63_n_0 ;
  wire \rgf_c1bus_wb[31]_i_64_n_0 ;
  wire \rgf_c1bus_wb[31]_i_65_n_0 ;
  wire \rgf_c1bus_wb[31]_i_66_n_0 ;
  wire \rgf_c1bus_wb[31]_i_67_n_0 ;
  wire \rgf_c1bus_wb[31]_i_70_n_0 ;
  wire \rgf_c1bus_wb[31]_i_71_n_0 ;
  wire \rgf_c1bus_wb[31]_i_72_n_0 ;
  wire \rgf_c1bus_wb[31]_i_73_n_0 ;
  wire \rgf_c1bus_wb[31]_i_74_n_0 ;
  wire \rgf_c1bus_wb[31]_i_75_n_0 ;
  wire \rgf_c1bus_wb[31]_i_76_n_0 ;
  wire \rgf_c1bus_wb[31]_i_77_n_0 ;
  wire \rgf_c1bus_wb[31]_i_78_n_0 ;
  wire \rgf_c1bus_wb[31]_i_83_n_0 ;
  wire \rgf_c1bus_wb[31]_i_85_n_0 ;
  wire \rgf_c1bus_wb[31]_i_87_n_0 ;
  wire \rgf_c1bus_wb[31]_i_88_n_0 ;
  wire \rgf_c1bus_wb[31]_i_89_n_0 ;
  wire \rgf_c1bus_wb[31]_i_8_n_0 ;
  wire \rgf_c1bus_wb[31]_i_90_n_0 ;
  wire \rgf_c1bus_wb[31]_i_9_n_0 ;
  wire \rgf_c1bus_wb[3]_i_10_n_0 ;
  wire \rgf_c1bus_wb[3]_i_11_n_0 ;
  wire \rgf_c1bus_wb[3]_i_12_n_0 ;
  wire \rgf_c1bus_wb[3]_i_13_n_0 ;
  wire \rgf_c1bus_wb[3]_i_14_n_0 ;
  wire \rgf_c1bus_wb[3]_i_15_n_0 ;
  wire \rgf_c1bus_wb[3]_i_16_n_0 ;
  wire \rgf_c1bus_wb[3]_i_17_n_0 ;
  wire \rgf_c1bus_wb[3]_i_18_n_0 ;
  wire \rgf_c1bus_wb[3]_i_19_n_0 ;
  wire \rgf_c1bus_wb[3]_i_21_n_0 ;
  wire \rgf_c1bus_wb[3]_i_22_n_0 ;
  wire \rgf_c1bus_wb[3]_i_23_n_0 ;
  wire \rgf_c1bus_wb[3]_i_24_n_0 ;
  wire \rgf_c1bus_wb[3]_i_25_n_0 ;
  wire \rgf_c1bus_wb[3]_i_26_n_0 ;
  wire \rgf_c1bus_wb[3]_i_2_n_0 ;
  wire \rgf_c1bus_wb[3]_i_31_n_0 ;
  wire \rgf_c1bus_wb[3]_i_3_n_0 ;
  wire \rgf_c1bus_wb[3]_i_4_n_0 ;
  wire \rgf_c1bus_wb[3]_i_5_n_0 ;
  wire \rgf_c1bus_wb[3]_i_6_n_0 ;
  wire \rgf_c1bus_wb[3]_i_7_n_0 ;
  wire \rgf_c1bus_wb[3]_i_8_n_0 ;
  wire \rgf_c1bus_wb[3]_i_9_n_0 ;
  wire \rgf_c1bus_wb[4]_i_10_n_0 ;
  wire \rgf_c1bus_wb[4]_i_11_n_0 ;
  wire \rgf_c1bus_wb[4]_i_12_n_0 ;
  wire \rgf_c1bus_wb[4]_i_13_n_0 ;
  wire \rgf_c1bus_wb[4]_i_14_n_0 ;
  wire \rgf_c1bus_wb[4]_i_15_n_0 ;
  wire \rgf_c1bus_wb[4]_i_16_n_0 ;
  wire \rgf_c1bus_wb[4]_i_17_n_0 ;
  wire \rgf_c1bus_wb[4]_i_18_n_0 ;
  wire \rgf_c1bus_wb[4]_i_19_n_0 ;
  wire \rgf_c1bus_wb[4]_i_20_n_0 ;
  wire \rgf_c1bus_wb[4]_i_21_n_0 ;
  wire \rgf_c1bus_wb[4]_i_22_n_0 ;
  wire \rgf_c1bus_wb[4]_i_23_n_0 ;
  wire \rgf_c1bus_wb[4]_i_24_n_0 ;
  wire \rgf_c1bus_wb[4]_i_25_n_0 ;
  wire \rgf_c1bus_wb[4]_i_26_n_0 ;
  wire \rgf_c1bus_wb[4]_i_27_n_0 ;
  wire \rgf_c1bus_wb[4]_i_2_n_0 ;
  wire \rgf_c1bus_wb[4]_i_30_n_0 ;
  wire \rgf_c1bus_wb[4]_i_31_n_0 ;
  wire \rgf_c1bus_wb[4]_i_3_n_0 ;
  wire \rgf_c1bus_wb[4]_i_4_n_0 ;
  wire \rgf_c1bus_wb[4]_i_5_n_0 ;
  wire \rgf_c1bus_wb[4]_i_6_n_0 ;
  wire \rgf_c1bus_wb[4]_i_7_n_0 ;
  wire \rgf_c1bus_wb[4]_i_8_n_0 ;
  wire \rgf_c1bus_wb[4]_i_9_n_0 ;
  wire \rgf_c1bus_wb[5]_i_10_n_0 ;
  wire \rgf_c1bus_wb[5]_i_11_n_0 ;
  wire \rgf_c1bus_wb[5]_i_12_n_0 ;
  wire \rgf_c1bus_wb[5]_i_13_n_0 ;
  wire \rgf_c1bus_wb[5]_i_14_n_0 ;
  wire \rgf_c1bus_wb[5]_i_15_n_0 ;
  wire \rgf_c1bus_wb[5]_i_16_n_0 ;
  wire \rgf_c1bus_wb[5]_i_17_n_0 ;
  wire \rgf_c1bus_wb[5]_i_18_n_0 ;
  wire \rgf_c1bus_wb[5]_i_19_n_0 ;
  wire \rgf_c1bus_wb[5]_i_20_n_0 ;
  wire \rgf_c1bus_wb[5]_i_21_n_0 ;
  wire \rgf_c1bus_wb[5]_i_22_n_0 ;
  wire \rgf_c1bus_wb[5]_i_23_n_0 ;
  wire \rgf_c1bus_wb[5]_i_24_n_0 ;
  wire \rgf_c1bus_wb[5]_i_25_n_0 ;
  wire \rgf_c1bus_wb[5]_i_26_n_0 ;
  wire \rgf_c1bus_wb[5]_i_27_n_0 ;
  wire \rgf_c1bus_wb[5]_i_2_n_0 ;
  wire \rgf_c1bus_wb[5]_i_3_n_0 ;
  wire \rgf_c1bus_wb[5]_i_4_n_0 ;
  wire \rgf_c1bus_wb[5]_i_5_n_0 ;
  wire \rgf_c1bus_wb[5]_i_6_n_0 ;
  wire \rgf_c1bus_wb[5]_i_7_n_0 ;
  wire \rgf_c1bus_wb[5]_i_8_n_0 ;
  wire \rgf_c1bus_wb[5]_i_9_n_0 ;
  wire \rgf_c1bus_wb[6]_i_10_n_0 ;
  wire \rgf_c1bus_wb[6]_i_11_n_0 ;
  wire \rgf_c1bus_wb[6]_i_12_n_0 ;
  wire \rgf_c1bus_wb[6]_i_13_n_0 ;
  wire \rgf_c1bus_wb[6]_i_14_n_0 ;
  wire \rgf_c1bus_wb[6]_i_15_n_0 ;
  wire \rgf_c1bus_wb[6]_i_16_n_0 ;
  wire \rgf_c1bus_wb[6]_i_17_n_0 ;
  wire \rgf_c1bus_wb[6]_i_18_n_0 ;
  wire \rgf_c1bus_wb[6]_i_19_n_0 ;
  wire \rgf_c1bus_wb[6]_i_20_n_0 ;
  wire \rgf_c1bus_wb[6]_i_21_n_0 ;
  wire \rgf_c1bus_wb[6]_i_22_n_0 ;
  wire \rgf_c1bus_wb[6]_i_23_n_0 ;
  wire \rgf_c1bus_wb[6]_i_24_n_0 ;
  wire \rgf_c1bus_wb[6]_i_25_n_0 ;
  wire \rgf_c1bus_wb[6]_i_26_n_0 ;
  wire \rgf_c1bus_wb[6]_i_2_n_0 ;
  wire \rgf_c1bus_wb[6]_i_3_n_0 ;
  wire \rgf_c1bus_wb[6]_i_4_n_0 ;
  wire \rgf_c1bus_wb[6]_i_5_n_0 ;
  wire \rgf_c1bus_wb[6]_i_6_n_0 ;
  wire \rgf_c1bus_wb[6]_i_7_n_0 ;
  wire \rgf_c1bus_wb[6]_i_8_n_0 ;
  wire \rgf_c1bus_wb[6]_i_9_n_0 ;
  wire \rgf_c1bus_wb[7]_i_10_n_0 ;
  wire \rgf_c1bus_wb[7]_i_11_n_0 ;
  wire \rgf_c1bus_wb[7]_i_12_n_0 ;
  wire \rgf_c1bus_wb[7]_i_13_n_0 ;
  wire \rgf_c1bus_wb[7]_i_14_n_0 ;
  wire \rgf_c1bus_wb[7]_i_15_n_0 ;
  wire \rgf_c1bus_wb[7]_i_16_n_0 ;
  wire \rgf_c1bus_wb[7]_i_17_n_0 ;
  wire \rgf_c1bus_wb[7]_i_18_n_0 ;
  wire \rgf_c1bus_wb[7]_i_19_n_0 ;
  wire \rgf_c1bus_wb[7]_i_20_n_0 ;
  wire \rgf_c1bus_wb[7]_i_21_n_0 ;
  wire \rgf_c1bus_wb[7]_i_22_n_0 ;
  wire \rgf_c1bus_wb[7]_i_24_n_0 ;
  wire \rgf_c1bus_wb[7]_i_25_n_0 ;
  wire \rgf_c1bus_wb[7]_i_26_n_0 ;
  wire \rgf_c1bus_wb[7]_i_27_n_0 ;
  wire \rgf_c1bus_wb[7]_i_28_n_0 ;
  wire \rgf_c1bus_wb[7]_i_29_n_0 ;
  wire \rgf_c1bus_wb[7]_i_2_n_0 ;
  wire \rgf_c1bus_wb[7]_i_30_n_0 ;
  wire \rgf_c1bus_wb[7]_i_35_n_0 ;
  wire \rgf_c1bus_wb[7]_i_3_n_0 ;
  wire \rgf_c1bus_wb[7]_i_4_n_0 ;
  wire \rgf_c1bus_wb[7]_i_5_n_0 ;
  wire \rgf_c1bus_wb[7]_i_6_n_0 ;
  wire \rgf_c1bus_wb[7]_i_7_n_0 ;
  wire \rgf_c1bus_wb[7]_i_8_n_0 ;
  wire \rgf_c1bus_wb[7]_i_9_n_0 ;
  wire \rgf_c1bus_wb[8]_i_10_n_0 ;
  wire \rgf_c1bus_wb[8]_i_11_n_0 ;
  wire \rgf_c1bus_wb[8]_i_12_n_0 ;
  wire \rgf_c1bus_wb[8]_i_13_n_0 ;
  wire \rgf_c1bus_wb[8]_i_14_n_0 ;
  wire \rgf_c1bus_wb[8]_i_15_n_0 ;
  wire \rgf_c1bus_wb[8]_i_16_n_0 ;
  wire \rgf_c1bus_wb[8]_i_17_n_0 ;
  wire \rgf_c1bus_wb[8]_i_18_n_0 ;
  wire \rgf_c1bus_wb[8]_i_19_n_0 ;
  wire \rgf_c1bus_wb[8]_i_20_n_0 ;
  wire \rgf_c1bus_wb[8]_i_21_n_0 ;
  wire \rgf_c1bus_wb[8]_i_22_n_0 ;
  wire \rgf_c1bus_wb[8]_i_23_n_0 ;
  wire \rgf_c1bus_wb[8]_i_24_n_0 ;
  wire \rgf_c1bus_wb[8]_i_25_n_0 ;
  wire \rgf_c1bus_wb[8]_i_26_n_0 ;
  wire \rgf_c1bus_wb[8]_i_27_n_0 ;
  wire \rgf_c1bus_wb[8]_i_2_n_0 ;
  wire \rgf_c1bus_wb[8]_i_3_n_0 ;
  wire \rgf_c1bus_wb[8]_i_4_n_0 ;
  wire \rgf_c1bus_wb[8]_i_5_n_0 ;
  wire \rgf_c1bus_wb[8]_i_6_n_0 ;
  wire \rgf_c1bus_wb[8]_i_7_n_0 ;
  wire \rgf_c1bus_wb[8]_i_8_n_0 ;
  wire \rgf_c1bus_wb[8]_i_9_n_0 ;
  wire \rgf_c1bus_wb[9]_i_10_n_0 ;
  wire \rgf_c1bus_wb[9]_i_11_n_0 ;
  wire \rgf_c1bus_wb[9]_i_12_n_0 ;
  wire \rgf_c1bus_wb[9]_i_13_n_0 ;
  wire \rgf_c1bus_wb[9]_i_14_n_0 ;
  wire \rgf_c1bus_wb[9]_i_15_n_0 ;
  wire \rgf_c1bus_wb[9]_i_16_n_0 ;
  wire \rgf_c1bus_wb[9]_i_17_n_0 ;
  wire \rgf_c1bus_wb[9]_i_18_n_0 ;
  wire \rgf_c1bus_wb[9]_i_19_n_0 ;
  wire \rgf_c1bus_wb[9]_i_20_n_0 ;
  wire \rgf_c1bus_wb[9]_i_21_n_0 ;
  wire \rgf_c1bus_wb[9]_i_22_n_0 ;
  wire \rgf_c1bus_wb[9]_i_23_n_0 ;
  wire \rgf_c1bus_wb[9]_i_24_n_0 ;
  wire \rgf_c1bus_wb[9]_i_25_n_0 ;
  wire \rgf_c1bus_wb[9]_i_26_n_0 ;
  wire \rgf_c1bus_wb[9]_i_2_n_0 ;
  wire \rgf_c1bus_wb[9]_i_3_n_0 ;
  wire \rgf_c1bus_wb[9]_i_4_n_0 ;
  wire \rgf_c1bus_wb[9]_i_5_n_0 ;
  wire \rgf_c1bus_wb[9]_i_6_n_0 ;
  wire \rgf_c1bus_wb[9]_i_7_n_0 ;
  wire \rgf_c1bus_wb[9]_i_8_n_0 ;
  wire \rgf_c1bus_wb[9]_i_9_n_0 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_0 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_1 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_2 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_3 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_4 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_5 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_6 ;
  wire \rgf_c1bus_wb_reg[11]_i_10_n_7 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_0 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_1 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_2 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_3 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_4 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_5 ;
  wire \rgf_c1bus_wb_reg[19]_i_10_n_7 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_0 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_1 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_2 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_3 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_4 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_5 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_6 ;
  wire \rgf_c1bus_wb_reg[19]_i_18_n_7 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_0 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_1 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_2 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_3 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_4 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_5 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_6 ;
  wire \rgf_c1bus_wb_reg[23]_i_11_n_7 ;
  wire \rgf_c1bus_wb_reg[24]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[24]_i_5_n_0 ;
  wire \rgf_c1bus_wb_reg[24]_i_6_n_0 ;
  wire \rgf_c1bus_wb_reg[26]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[26]_i_5_n_0 ;
  wire \rgf_c1bus_wb_reg[26]_i_6_n_0 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_0 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_1 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_2 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_3 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_4 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_5 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_6 ;
  wire \rgf_c1bus_wb_reg[27]_i_10_n_7 ;
  wire \rgf_c1bus_wb_reg[30]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[30]_i_5_n_0 ;
  wire \rgf_c1bus_wb_reg[30]_i_6_n_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_1 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_2 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_3 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_4 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_5 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_6 ;
  wire \rgf_c1bus_wb_reg[31]_i_11_n_7 ;
  wire \rgf_c1bus_wb_reg[31]_i_2_n_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_6_n_0 ;
  wire \rgf_c1bus_wb_reg[31]_i_7_n_0 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_0 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_1 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_2 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_3 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_4 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_5 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_6 ;
  wire \rgf_c1bus_wb_reg[3]_i_20_n_7 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_0 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_1 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_2 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_3 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_4 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_5 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_6 ;
  wire \rgf_c1bus_wb_reg[7]_i_23_n_7 ;
  wire \rgf_selc0_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_1_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_1_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_24_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_25_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_26_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_27_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc0_rn_wb[2]_i_9_n_0 ;
  wire rgf_selc0_stat_i_1_n_0;
  wire rgf_selc0_stat_i_2_n_0;
  wire \rgf_selc0_wb[0]_i_10_n_0 ;
  wire \rgf_selc0_wb[0]_i_11_n_0 ;
  wire \rgf_selc0_wb[0]_i_12_n_0 ;
  wire \rgf_selc0_wb[0]_i_13_n_0 ;
  wire \rgf_selc0_wb[0]_i_14_n_0 ;
  wire \rgf_selc0_wb[0]_i_15_n_0 ;
  wire \rgf_selc0_wb[0]_i_16_n_0 ;
  wire \rgf_selc0_wb[0]_i_17_n_0 ;
  wire \rgf_selc0_wb[0]_i_2_n_0 ;
  wire \rgf_selc0_wb[0]_i_3_n_0 ;
  wire \rgf_selc0_wb[0]_i_4_n_0 ;
  wire \rgf_selc0_wb[0]_i_5_n_0 ;
  wire \rgf_selc0_wb[0]_i_6_n_0 ;
  wire \rgf_selc0_wb[0]_i_7_n_0 ;
  wire \rgf_selc0_wb[0]_i_8_n_0 ;
  wire \rgf_selc0_wb[0]_i_9_n_0 ;
  wire \rgf_selc0_wb[1]_i_10_n_0 ;
  wire \rgf_selc0_wb[1]_i_11_n_0 ;
  wire \rgf_selc0_wb[1]_i_12_n_0 ;
  wire \rgf_selc0_wb[1]_i_13_n_0 ;
  wire \rgf_selc0_wb[1]_i_14_n_0 ;
  wire \rgf_selc0_wb[1]_i_15_n_0 ;
  wire \rgf_selc0_wb[1]_i_16_n_0 ;
  wire \rgf_selc0_wb[1]_i_17_n_0 ;
  wire \rgf_selc0_wb[1]_i_18_n_0 ;
  wire \rgf_selc0_wb[1]_i_19_n_0 ;
  wire \rgf_selc0_wb[1]_i_20_n_0 ;
  wire \rgf_selc0_wb[1]_i_21_n_0 ;
  wire \rgf_selc0_wb[1]_i_22_n_0 ;
  wire \rgf_selc0_wb[1]_i_23_n_0 ;
  wire \rgf_selc0_wb[1]_i_24_n_0 ;
  wire \rgf_selc0_wb[1]_i_25_n_0 ;
  wire \rgf_selc0_wb[1]_i_26_n_0 ;
  wire \rgf_selc0_wb[1]_i_27_n_0 ;
  wire \rgf_selc0_wb[1]_i_28_n_0 ;
  wire \rgf_selc0_wb[1]_i_29_n_0 ;
  wire \rgf_selc0_wb[1]_i_2_n_0 ;
  wire \rgf_selc0_wb[1]_i_30_n_0 ;
  wire \rgf_selc0_wb[1]_i_31_n_0 ;
  wire \rgf_selc0_wb[1]_i_32_n_0 ;
  wire \rgf_selc0_wb[1]_i_33_n_0 ;
  wire \rgf_selc0_wb[1]_i_34_n_0 ;
  wire \rgf_selc0_wb[1]_i_35_n_0 ;
  wire \rgf_selc0_wb[1]_i_36_n_0 ;
  wire \rgf_selc0_wb[1]_i_37_n_0 ;
  wire \rgf_selc0_wb[1]_i_38_n_0 ;
  wire \rgf_selc0_wb[1]_i_39_n_0 ;
  wire \rgf_selc0_wb[1]_i_3_n_0 ;
  wire \rgf_selc0_wb[1]_i_4_n_0 ;
  wire \rgf_selc0_wb[1]_i_5_n_0 ;
  wire \rgf_selc0_wb[1]_i_6_n_0 ;
  wire \rgf_selc0_wb[1]_i_7_n_0 ;
  wire \rgf_selc0_wb[1]_i_8_n_0 ;
  wire \rgf_selc0_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_29_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_30_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_31_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_32_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_33_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_34_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_35_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_1_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_29_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_30_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_31_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_10_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_11_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_12_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_13_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_14_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_15_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_16_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_17_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_18_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_19_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_1_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_20_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_21_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_22_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_23_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_24_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_25_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_26_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_27_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_28_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_2_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_3_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_4_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_5_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_6_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_7_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_8_n_0 ;
  wire \rgf_selc1_rn_wb[2]_i_9_n_0 ;
  wire rgf_selc1_stat_i_1_n_0;
  wire rgf_selc1_stat_i_2_n_0;
  wire \rgf_selc1_wb[0]_i_10_n_0 ;
  wire \rgf_selc1_wb[0]_i_11_n_0 ;
  wire \rgf_selc1_wb[0]_i_12_n_0 ;
  wire \rgf_selc1_wb[0]_i_13_n_0 ;
  wire \rgf_selc1_wb[0]_i_14_n_0 ;
  wire \rgf_selc1_wb[0]_i_15_n_0 ;
  wire \rgf_selc1_wb[0]_i_16_n_0 ;
  wire \rgf_selc1_wb[0]_i_17_n_0 ;
  wire \rgf_selc1_wb[0]_i_18_n_0 ;
  wire \rgf_selc1_wb[0]_i_19_n_0 ;
  wire \rgf_selc1_wb[0]_i_20_n_0 ;
  wire \rgf_selc1_wb[0]_i_2_n_0 ;
  wire \rgf_selc1_wb[0]_i_3_n_0 ;
  wire \rgf_selc1_wb[0]_i_4_n_0 ;
  wire \rgf_selc1_wb[0]_i_5_n_0 ;
  wire \rgf_selc1_wb[0]_i_6_n_0 ;
  wire \rgf_selc1_wb[0]_i_7_n_0 ;
  wire \rgf_selc1_wb[0]_i_8_n_0 ;
  wire \rgf_selc1_wb[0]_i_9_n_0 ;
  wire \rgf_selc1_wb[1]_i_10_n_0 ;
  wire \rgf_selc1_wb[1]_i_11_n_0 ;
  wire \rgf_selc1_wb[1]_i_12_n_0 ;
  wire \rgf_selc1_wb[1]_i_13_n_0 ;
  wire \rgf_selc1_wb[1]_i_14_n_0 ;
  wire \rgf_selc1_wb[1]_i_15_n_0 ;
  wire \rgf_selc1_wb[1]_i_16_n_0 ;
  wire \rgf_selc1_wb[1]_i_17_n_0 ;
  wire \rgf_selc1_wb[1]_i_18_n_0 ;
  wire \rgf_selc1_wb[1]_i_19_n_0 ;
  wire \rgf_selc1_wb[1]_i_20_n_0 ;
  wire \rgf_selc1_wb[1]_i_21_n_0 ;
  wire \rgf_selc1_wb[1]_i_22_n_0 ;
  wire \rgf_selc1_wb[1]_i_23_n_0 ;
  wire \rgf_selc1_wb[1]_i_24_n_0 ;
  wire \rgf_selc1_wb[1]_i_25_n_0 ;
  wire \rgf_selc1_wb[1]_i_26_n_0 ;
  wire \rgf_selc1_wb[1]_i_27_n_0 ;
  wire \rgf_selc1_wb[1]_i_28_n_0 ;
  wire \rgf_selc1_wb[1]_i_29_n_0 ;
  wire \rgf_selc1_wb[1]_i_2_n_0 ;
  wire \rgf_selc1_wb[1]_i_30_n_0 ;
  wire \rgf_selc1_wb[1]_i_31_n_0 ;
  wire \rgf_selc1_wb[1]_i_32_n_0 ;
  wire \rgf_selc1_wb[1]_i_33_n_0 ;
  wire \rgf_selc1_wb[1]_i_34_n_0 ;
  wire \rgf_selc1_wb[1]_i_35_n_0 ;
  wire \rgf_selc1_wb[1]_i_36_n_0 ;
  wire \rgf_selc1_wb[1]_i_37_n_0 ;
  wire \rgf_selc1_wb[1]_i_38_n_0 ;
  wire \rgf_selc1_wb[1]_i_39_n_0 ;
  wire \rgf_selc1_wb[1]_i_3_n_0 ;
  wire \rgf_selc1_wb[1]_i_40_n_0 ;
  wire \rgf_selc1_wb[1]_i_41_n_0 ;
  wire \rgf_selc1_wb[1]_i_42_n_0 ;
  wire \rgf_selc1_wb[1]_i_5_n_0 ;
  wire \rgf_selc1_wb[1]_i_6_n_0 ;
  wire \rgf_selc1_wb[1]_i_7_n_0 ;
  wire \rgf_selc1_wb[1]_i_8_n_0 ;
  wire \rgf_selc1_wb[1]_i_9_n_0 ;
  wire \rgf_selc1_wb_reg[1]_i_4_n_0 ;
  wire rst_n;
  wire \sp[0]_i_1_n_0 ;
  wire \sp[0]_i_2_n_0 ;
  wire \sp[10]_i_1_n_0 ;
  wire \sp[10]_i_2_n_0 ;
  wire \sp[11]_i_1_n_0 ;
  wire \sp[11]_i_2_n_0 ;
  wire \sp[12]_i_1_n_0 ;
  wire \sp[12]_i_2_n_0 ;
  wire \sp[13]_i_1_n_0 ;
  wire \sp[13]_i_2_n_0 ;
  wire \sp[14]_i_1_n_0 ;
  wire \sp[14]_i_2_n_0 ;
  wire \sp[15]_i_1_n_0 ;
  wire \sp[15]_i_2_n_0 ;
  wire \sp[16]_i_1_n_0 ;
  wire \sp[16]_i_2_n_0 ;
  wire \sp[17]_i_1_n_0 ;
  wire \sp[17]_i_2_n_0 ;
  wire \sp[18]_i_1_n_0 ;
  wire \sp[18]_i_2_n_0 ;
  wire \sp[19]_i_1_n_0 ;
  wire \sp[19]_i_2_n_0 ;
  wire \sp[1]_i_1_n_0 ;
  wire \sp[1]_i_2_n_0 ;
  wire \sp[20]_i_1_n_0 ;
  wire \sp[20]_i_2_n_0 ;
  wire \sp[21]_i_1_n_0 ;
  wire \sp[21]_i_2_n_0 ;
  wire \sp[22]_i_1_n_0 ;
  wire \sp[22]_i_2_n_0 ;
  wire \sp[23]_i_1_n_0 ;
  wire \sp[23]_i_2_n_0 ;
  wire \sp[24]_i_1_n_0 ;
  wire \sp[24]_i_2_n_0 ;
  wire \sp[25]_i_1_n_0 ;
  wire \sp[25]_i_2_n_0 ;
  wire \sp[26]_i_1_n_0 ;
  wire \sp[26]_i_2_n_0 ;
  wire \sp[27]_i_1_n_0 ;
  wire \sp[27]_i_2_n_0 ;
  wire \sp[28]_i_1_n_0 ;
  wire \sp[28]_i_2_n_0 ;
  wire \sp[29]_i_1_n_0 ;
  wire \sp[29]_i_2_n_0 ;
  wire \sp[2]_i_1_n_0 ;
  wire \sp[2]_i_2_n_0 ;
  wire \sp[30]_i_1_n_0 ;
  wire \sp[30]_i_2_n_0 ;
  wire \sp[31]_i_10_n_0 ;
  wire \sp[31]_i_11_n_0 ;
  wire \sp[31]_i_12_n_0 ;
  wire \sp[31]_i_15_n_0 ;
  wire \sp[31]_i_16_n_0 ;
  wire \sp[31]_i_17_n_0 ;
  wire \sp[31]_i_18_n_0 ;
  wire \sp[31]_i_19_n_0 ;
  wire \sp[31]_i_1_n_0 ;
  wire \sp[31]_i_20_n_0 ;
  wire \sp[31]_i_21_n_0 ;
  wire \sp[31]_i_22_n_0 ;
  wire \sp[31]_i_24_n_0 ;
  wire \sp[31]_i_25_n_0 ;
  wire \sp[31]_i_26_n_0 ;
  wire \sp[31]_i_27_n_0 ;
  wire \sp[31]_i_28_n_0 ;
  wire \sp[31]_i_29_n_0 ;
  wire \sp[31]_i_2_n_0 ;
  wire \sp[31]_i_30_n_0 ;
  wire \sp[31]_i_31_n_0 ;
  wire \sp[31]_i_32_n_0 ;
  wire \sp[31]_i_7_n_0 ;
  wire \sp[31]_i_8_n_0 ;
  wire \sp[3]_i_1_n_0 ;
  wire \sp[3]_i_2_n_0 ;
  wire \sp[3]_i_4_n_0 ;
  wire \sp[3]_i_5_n_0 ;
  wire \sp[4]_i_1_n_0 ;
  wire \sp[4]_i_2_n_0 ;
  wire \sp[5]_i_1_n_0 ;
  wire \sp[5]_i_2_n_0 ;
  wire \sp[6]_i_1_n_0 ;
  wire \sp[6]_i_2_n_0 ;
  wire \sp[7]_i_1_n_0 ;
  wire \sp[7]_i_2_n_0 ;
  wire \sp[8]_i_1_n_0 ;
  wire \sp[8]_i_2_n_0 ;
  wire \sp[9]_i_1_n_0 ;
  wire \sp[9]_i_2_n_0 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[15]_i_3_n_0 ;
  wire \sp_reg[15]_i_3_n_1 ;
  wire \sp_reg[15]_i_3_n_2 ;
  wire \sp_reg[15]_i_3_n_3 ;
  wire \sp_reg[19]_i_5_n_0 ;
  wire \sp_reg[19]_i_5_n_1 ;
  wire \sp_reg[19]_i_5_n_2 ;
  wire \sp_reg[19]_i_5_n_3 ;
  wire \sp_reg[23]_i_5_n_0 ;
  wire \sp_reg[23]_i_5_n_1 ;
  wire \sp_reg[23]_i_5_n_2 ;
  wire \sp_reg[23]_i_5_n_3 ;
  wire \sp_reg[27]_i_5_n_0 ;
  wire \sp_reg[27]_i_5_n_1 ;
  wire \sp_reg[27]_i_5_n_2 ;
  wire \sp_reg[27]_i_5_n_3 ;
  wire \sp_reg[31]_i_23_n_0 ;
  wire \sp_reg[31]_i_9_n_1 ;
  wire \sp_reg[31]_i_9_n_2 ;
  wire \sp_reg[31]_i_9_n_3 ;
  wire \sp_reg[3]_i_3_n_0 ;
  wire \sp_reg[3]_i_3_n_1 ;
  wire \sp_reg[3]_i_3_n_2 ;
  wire \sp_reg[3]_i_3_n_3 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sr[0]_i_2_n_0 ;
  wire \sr[10]_i_2_n_0 ;
  wire \sr[11]_i_12_n_0 ;
  wire \sr[11]_i_13_n_0 ;
  wire \sr[11]_i_14_n_0 ;
  wire \sr[11]_i_15_n_0 ;
  wire \sr[11]_i_16_n_0 ;
  wire \sr[11]_i_2_n_0 ;
  wire \sr[11]_i_3_n_0 ;
  wire \sr[11]_i_4_n_0 ;
  wire \sr[13]_i_2_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire \sr[15]_i_10_n_0 ;
  wire \sr[15]_i_2_n_0 ;
  wire \sr[15]_i_6_n_0 ;
  wire \sr[15]_i_7_n_0 ;
  wire \sr[15]_i_8_n_0 ;
  wire \sr[15]_i_9_n_0 ;
  wire \sr[1]_i_2_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[2]_i_3_n_0 ;
  wire \sr[2]_i_4_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[3]_i_3_n_0 ;
  wire \sr[3]_i_4_n_0 ;
  wire \sr[3]_i_5_n_0 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_14_n_0 ;
  wire \sr[4]_i_15_n_0 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_17_n_0 ;
  wire \sr[4]_i_18_n_0 ;
  wire \sr[4]_i_19_n_0 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_25_n_0 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_29_n_0 ;
  wire \sr[4]_i_2_n_0 ;
  wire \sr[4]_i_30_n_0 ;
  wire \sr[4]_i_31_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_35_n_0 ;
  wire \sr[4]_i_36_n_0 ;
  wire \sr[4]_i_37_n_0 ;
  wire \sr[4]_i_38_n_0 ;
  wire \sr[4]_i_39_n_0 ;
  wire \sr[4]_i_40_n_0 ;
  wire \sr[4]_i_41_n_0 ;
  wire \sr[4]_i_42_n_0 ;
  wire \sr[4]_i_43_n_0 ;
  wire \sr[4]_i_44_n_0 ;
  wire \sr[4]_i_45_n_0 ;
  wire \sr[4]_i_46_n_0 ;
  wire \sr[4]_i_47_n_0 ;
  wire \sr[4]_i_48_n_0 ;
  wire \sr[4]_i_49_n_0 ;
  wire \sr[4]_i_4_n_0 ;
  wire \sr[4]_i_50_n_0 ;
  wire \sr[4]_i_51_n_0 ;
  wire \sr[4]_i_52_n_0 ;
  wire \sr[4]_i_53_n_0 ;
  wire \sr[4]_i_54_n_0 ;
  wire \sr[4]_i_55_n_0 ;
  wire \sr[4]_i_56_n_0 ;
  wire \sr[4]_i_57_n_0 ;
  wire \sr[4]_i_58_n_0 ;
  wire \sr[4]_i_59_n_0 ;
  wire \sr[4]_i_5_n_0 ;
  wire \sr[4]_i_60_n_0 ;
  wire \sr[4]_i_61_n_0 ;
  wire \sr[4]_i_62_n_0 ;
  wire \sr[4]_i_63_n_0 ;
  wire \sr[4]_i_64_n_0 ;
  wire \sr[4]_i_65_n_0 ;
  wire \sr[4]_i_66_n_0 ;
  wire \sr[4]_i_67_n_0 ;
  wire \sr[4]_i_68_n_0 ;
  wire \sr[4]_i_69_n_0 ;
  wire \sr[4]_i_6_n_0 ;
  wire \sr[4]_i_70_n_0 ;
  wire \sr[4]_i_71_n_0 ;
  wire \sr[4]_i_72_n_0 ;
  wire \sr[4]_i_73_n_0 ;
  wire \sr[4]_i_74_n_0 ;
  wire \sr[4]_i_75_n_0 ;
  wire \sr[4]_i_76_n_0 ;
  wire \sr[4]_i_77_n_0 ;
  wire \sr[4]_i_78_n_0 ;
  wire \sr[4]_i_79_n_0 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[4]_i_80_n_0 ;
  wire \sr[4]_i_81_n_0 ;
  wire \sr[4]_i_82_n_0 ;
  wire \sr[4]_i_83_n_0 ;
  wire \sr[4]_i_84_n_0 ;
  wire \sr[4]_i_85_n_0 ;
  wire \sr[4]_i_86_n_0 ;
  wire \sr[4]_i_87_n_0 ;
  wire \sr[4]_i_88_n_0 ;
  wire \sr[4]_i_89_n_0 ;
  wire \sr[4]_i_8_n_0 ;
  wire \sr[4]_i_90_n_0 ;
  wire \sr[4]_i_91_n_0 ;
  wire \sr[4]_i_92_n_0 ;
  wire \sr[4]_i_93_n_0 ;
  wire \sr[4]_i_94_n_0 ;
  wire \sr[4]_i_95_n_0 ;
  wire \sr[4]_i_96_n_0 ;
  wire \sr[4]_i_97_n_0 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_10_n_0 ;
  wire \sr[5]_i_11_n_0 ;
  wire \sr[5]_i_12_n_0 ;
  wire \sr[5]_i_13_n_0 ;
  wire \sr[5]_i_14_n_0 ;
  wire \sr[5]_i_15_n_0 ;
  wire \sr[5]_i_17_n_0 ;
  wire \sr[5]_i_18_n_0 ;
  wire \sr[5]_i_20_n_0 ;
  wire \sr[5]_i_21_n_0 ;
  wire \sr[5]_i_22_n_0 ;
  wire \sr[5]_i_23_n_0 ;
  wire \sr[5]_i_2_n_0 ;
  wire \sr[5]_i_3_n_0 ;
  wire \sr[5]_i_6_n_0 ;
  wire \sr[5]_i_7_n_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[5]_i_9_n_0 ;
  wire \sr[6]_i_10_n_0 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_12_n_0 ;
  wire \sr[6]_i_13_n_0 ;
  wire \sr[6]_i_16_n_0 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr[6]_i_18_n_0 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_21_n_0 ;
  wire \sr[6]_i_22_n_0 ;
  wire \sr[6]_i_23_n_0 ;
  wire \sr[6]_i_24_n_0 ;
  wire \sr[6]_i_25_n_0 ;
  wire \sr[6]_i_26_n_0 ;
  wire \sr[6]_i_27_n_0 ;
  wire \sr[6]_i_28_n_0 ;
  wire \sr[6]_i_30_n_0 ;
  wire \sr[6]_i_31_n_0 ;
  wire \sr[6]_i_32_n_0 ;
  wire \sr[6]_i_33_n_0 ;
  wire \sr[6]_i_34_n_0 ;
  wire \sr[6]_i_35_n_0 ;
  wire \sr[6]_i_36_n_0 ;
  wire \sr[6]_i_37_n_0 ;
  wire \sr[6]_i_38_n_0 ;
  wire \sr[6]_i_39_n_0 ;
  wire \sr[6]_i_40_n_0 ;
  wire \sr[6]_i_41_n_0 ;
  wire \sr[6]_i_42_n_0 ;
  wire \sr[6]_i_43_n_0 ;
  wire \sr[6]_i_44_n_0 ;
  wire \sr[6]_i_45_n_0 ;
  wire \sr[6]_i_46_n_0 ;
  wire \sr[6]_i_4_n_0 ;
  wire \sr[6]_i_5_n_0 ;
  wire \sr[6]_i_6_n_0 ;
  wire \sr[6]_i_7_n_0 ;
  wire \sr[6]_i_8_n_0 ;
  wire \sr[6]_i_9_n_0 ;
  wire \sr[7]_i_11_n_0 ;
  wire \sr[7]_i_12_n_0 ;
  wire \sr[7]_i_2_n_0 ;
  wire \sr[7]_i_3_n_0 ;
  wire \sr[7]_i_4_n_0 ;
  wire \sr[7]_i_5_n_0 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_8_n_0 ;
  wire \sr[7]_i_9_n_0 ;
  wire \sr[8]_i_2_n_0 ;
  wire \sr[9]_i_2_n_0 ;
  wire [2:0]stat;
  wire \stat[0]_i_10__0_n_0 ;
  wire \stat[0]_i_10__1_n_0 ;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_11__0_n_0 ;
  wire \stat[0]_i_11__1_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12__0_n_0 ;
  wire \stat[0]_i_12__1_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13__0_n_0 ;
  wire \stat[0]_i_13__1_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14__0_n_0 ;
  wire \stat[0]_i_14__1_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15__0_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16__0_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_17__0_n_0 ;
  wire \stat[0]_i_17_n_0 ;
  wire \stat[0]_i_18__0_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_19__0_n_0 ;
  wire \stat[0]_i_19_n_0 ;
  wire \stat[0]_i_1__2_n_0 ;
  wire \stat[0]_i_20__0_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21__0_n_0 ;
  wire \stat[0]_i_21_n_0 ;
  wire \stat[0]_i_22__0_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23__0_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24__0_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25__0_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26__0_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_27__0_n_0 ;
  wire \stat[0]_i_27_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2__0_n_0 ;
  wire \stat[0]_i_2__1_n_0 ;
  wire \stat[0]_i_2__2_n_0 ;
  wire \stat[0]_i_2_n_0 ;
  wire \stat[0]_i_3__0_n_0 ;
  wire \stat[0]_i_3__1_n_0 ;
  wire \stat[0]_i_3__2_n_0 ;
  wire \stat[0]_i_3_n_0 ;
  wire \stat[0]_i_4__0_n_0 ;
  wire \stat[0]_i_4__1_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5__0_n_0 ;
  wire \stat[0]_i_5__1_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6__0_n_0 ;
  wire \stat[0]_i_6__1_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7__0_n_0 ;
  wire \stat[0]_i_7__1_n_0 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8__0_n_0 ;
  wire \stat[0]_i_8__1_n_0 ;
  wire \stat[0]_i_8_n_0 ;
  wire \stat[0]_i_9__0_n_0 ;
  wire \stat[0]_i_9__1_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_10__0_n_0 ;
  wire \stat[1]_i_10_n_0 ;
  wire \stat[1]_i_11__0_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_12__0_n_0 ;
  wire \stat[1]_i_12_n_0 ;
  wire \stat[1]_i_13__0_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_14__0_n_0 ;
  wire \stat[1]_i_14_n_0 ;
  wire \stat[1]_i_15__0_n_0 ;
  wire \stat[1]_i_15_n_0 ;
  wire \stat[1]_i_16__0_n_0 ;
  wire \stat[1]_i_16_n_0 ;
  wire \stat[1]_i_17__0_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18__0_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_19__0_n_0 ;
  wire \stat[1]_i_19_n_0 ;
  wire \stat[1]_i_20__0_n_0 ;
  wire \stat[1]_i_20_n_0 ;
  wire \stat[1]_i_21__0_n_0 ;
  wire \stat[1]_i_21_n_0 ;
  wire \stat[1]_i_22__0_n_0 ;
  wire \stat[1]_i_22_n_0 ;
  wire \stat[1]_i_23__0_n_0 ;
  wire \stat[1]_i_23_n_0 ;
  wire \stat[1]_i_24__0_n_0 ;
  wire \stat[1]_i_24_n_0 ;
  wire \stat[1]_i_25_n_0 ;
  wire \stat[1]_i_26_n_0 ;
  wire \stat[1]_i_27_n_0 ;
  wire \stat[1]_i_2__0_n_0 ;
  wire \stat[1]_i_2__1_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3__0_n_0 ;
  wire \stat[1]_i_3__1_n_0 ;
  wire \stat[1]_i_3_n_0 ;
  wire \stat[1]_i_4__0_n_0 ;
  wire \stat[1]_i_4_n_0 ;
  wire \stat[1]_i_5__0_n_0 ;
  wire \stat[1]_i_5_n_0 ;
  wire \stat[1]_i_6__0_n_0 ;
  wire \stat[1]_i_6_n_0 ;
  wire \stat[1]_i_7__0_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8__0_n_0 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[1]_i_9__0_n_0 ;
  wire \stat[1]_i_9_n_0 ;
  wire \stat[2]_i_10__0_n_0 ;
  wire \stat[2]_i_10_n_0 ;
  wire \stat[2]_i_11__0_n_0 ;
  wire \stat[2]_i_11_n_0 ;
  wire \stat[2]_i_12__0_n_0 ;
  wire \stat[2]_i_12_n_0 ;
  wire \stat[2]_i_13__0_n_0 ;
  wire \stat[2]_i_13_n_0 ;
  wire \stat[2]_i_14__0_n_0 ;
  wire \stat[2]_i_14_n_0 ;
  wire \stat[2]_i_15_n_0 ;
  wire \stat[2]_i_16_n_0 ;
  wire \stat[2]_i_1__1_n_0 ;
  wire \stat[2]_i_1_n_0 ;
  wire \stat[2]_i_2__0_n_0 ;
  wire \stat[2]_i_2__1_n_0 ;
  wire \stat[2]_i_3__0_n_0 ;
  wire \stat[2]_i_3__1_n_0 ;
  wire \stat[2]_i_3_n_0 ;
  wire \stat[2]_i_4__0_n_0 ;
  wire \stat[2]_i_4_n_0 ;
  wire \stat[2]_i_5__0_n_0 ;
  wire \stat[2]_i_5_n_0 ;
  wire \stat[2]_i_6__0_n_0 ;
  wire \stat[2]_i_6_n_0 ;
  wire \stat[2]_i_7__0_n_0 ;
  wire \stat[2]_i_7_n_0 ;
  wire \stat[2]_i_8__0_n_0 ;
  wire \stat[2]_i_8_n_0 ;
  wire \stat[2]_i_9__0_n_0 ;
  wire \stat[2]_i_9_n_0 ;
  wire \tr[31]_i_4_n_0 ;
  wire [3:0]\NLW_pc0_reg[3]_i_3_O_UNCONNECTED ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(a0bus_0[0]),
        .I1(ccmd[4]),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(a0bus_0[10]),
        .I1(ccmd[4]),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(a0bus_0[11]),
        .I1(ccmd[4]),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(a0bus_0[12]),
        .I1(ccmd[4]),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(a0bus_0[13]),
        .I1(ccmd[4]),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(a0bus_0[14]),
        .I1(ccmd[4]),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(a0bus_0[15]),
        .I1(ccmd[4]),
        .O(abus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[16]_INST_0 
       (.I0(a0bus_0[16]),
        .I1(ccmd[4]),
        .O(abus_o[16]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[17]_INST_0 
       (.I0(a0bus_0[17]),
        .I1(ccmd[4]),
        .O(abus_o[17]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[18]_INST_0 
       (.I0(a0bus_0[18]),
        .I1(ccmd[4]),
        .O(abus_o[18]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[19]_INST_0 
       (.I0(a0bus_0[19]),
        .I1(ccmd[4]),
        .O(abus_o[19]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(a0bus_0[1]),
        .I1(ccmd[4]),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[20]_INST_0 
       (.I0(a0bus_0[20]),
        .I1(ccmd[4]),
        .O(abus_o[20]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[21]_INST_0 
       (.I0(a0bus_0[21]),
        .I1(ccmd[4]),
        .O(abus_o[21]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[22]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[22]),
        .O(abus_o[22]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[23]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[23]),
        .O(abus_o[23]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[24]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[24]),
        .O(abus_o[24]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[25]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[25]),
        .O(abus_o[25]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[26]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[26]),
        .O(abus_o[26]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[27]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[27]),
        .O(abus_o[27]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[28]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[28]),
        .O(abus_o[28]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[29]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[29]),
        .O(abus_o[29]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(a0bus_0[2]),
        .I1(ccmd[4]),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[30]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[30]),
        .O(abus_o[30]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[31]_INST_0 
       (.I0(ccmd[4]),
        .I1(a0bus_0[31]),
        .O(abus_o[31]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(a0bus_0[3]),
        .I1(ccmd[4]),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(a0bus_0[4]),
        .I1(ccmd[4]),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(a0bus_0[5]),
        .I1(ccmd[4]),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(a0bus_0[6]),
        .I1(ccmd[4]),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(a0bus_0[7]),
        .I1(ccmd[4]),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(a0bus_0[8]),
        .I1(ccmd[4]),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(a0bus_0[9]),
        .I1(ccmd[4]),
        .O(abus_o[9]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [7]),
        .O(add_out0_carry__0_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_14_n_0),
        .I3(\alu0/div/rem [6]),
        .I4(\alu0/div/dso_0 [6]),
        .O(\alu0/div/p_0_out [6]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_14__0_n_0),
        .I3(\alu1/div/rem [6]),
        .I4(\alu1/div/dso_0 [6]),
        .O(\alu1/div/p_0_out [6]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_15_n_0),
        .I3(\alu0/div/rem [5]),
        .I4(\alu0/div/dso_0 [5]),
        .O(\alu0/div/p_0_out [5]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_15__0_n_0),
        .I3(\alu1/div/rem [5]),
        .I4(\alu1/div/dso_0 [5]),
        .O(\alu1/div/p_0_out [5]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_16_n_0),
        .I3(\alu0/div/rem [4]),
        .I4(\alu0/div/dso_0 [4]),
        .O(\alu0/div/p_0_out [4]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_16__0_n_0),
        .I3(\alu1/div/rem [4]),
        .I4(\alu1/div/dso_0 [4]),
        .O(\alu1/div/p_0_out [4]));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__0_i_13
       (.I0(\alu0/div/quo [7]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [7]),
        .I4(\alu0/div/den [7]),
        .O(add_out0_carry__0_i_13_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__0_i_13__0
       (.I0(\alu1/div/quo [7]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [7]),
        .I4(\alu1/div/den [7]),
        .O(add_out0_carry__0_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_14
       (.I0(\alu0/div/den [6]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [6]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [6]),
        .O(add_out0_carry__0_i_14_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_14__0
       (.I0(\alu1/div/den [6]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [6]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [6]),
        .O(add_out0_carry__0_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__0_i_15
       (.I0(\alu0/div/quo [5]),
        .I1(\alu0/div/dso_0 [5]),
        .I2(\alu0/div/den [5]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__0_i_15_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__0_i_15__0
       (.I0(\alu1/div/quo [5]),
        .I1(\alu1/div/dso_0 [5]),
        .I2(\alu1/div/den [5]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__0_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_16
       (.I0(\alu0/div/den [4]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [4]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [4]),
        .O(add_out0_carry__0_i_16_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__0_i_16__0
       (.I0(\alu1/div/den [4]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [4]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [4]),
        .O(add_out0_carry__0_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [7]),
        .O(add_out0_carry__0_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [6]),
        .O(add_out0_carry__0_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [6]),
        .O(add_out0_carry__0_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [5]),
        .O(add_out0_carry__0_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [5]),
        .O(add_out0_carry__0_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [4]),
        .O(add_out0_carry__0_i_4_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__0_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [4]),
        .O(add_out0_carry__0_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [7]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [7]),
        .O(add_out0_carry__0_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [7]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [7]),
        .O(add_out0_carry__0_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [6]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [6]),
        .O(add_out0_carry__0_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [6]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [6]),
        .O(add_out0_carry__0_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [5]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [5]),
        .O(add_out0_carry__0_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [5]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [5]),
        .O(add_out0_carry__0_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [4]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [4]),
        .O(add_out0_carry__0_i_8_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__0_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [4]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [4]),
        .O(add_out0_carry__0_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__0_i_13_n_0),
        .I3(\alu0/div/rem [7]),
        .I4(\alu0/div/dso_0 [7]),
        .O(\alu0/div/p_0_out [7]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__0_i_13__0_n_0),
        .I3(\alu1/div/rem [7]),
        .I4(\alu1/div/dso_0 [7]),
        .O(\alu1/div/p_0_out [7]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [11]),
        .O(add_out0_carry__1_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_14_n_0),
        .I3(\alu0/div/rem [10]),
        .I4(\alu0/div/dso_0 [10]),
        .O(\alu0/div/p_0_out [10]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_14__0_n_0),
        .I3(\alu1/div/rem [10]),
        .I4(\alu1/div/dso_0 [10]),
        .O(\alu1/div/p_0_out [10]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_15_n_0),
        .I3(\alu0/div/rem [9]),
        .I4(\alu0/div/dso_0 [9]),
        .O(\alu0/div/p_0_out [9]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_15__0_n_0),
        .I3(\alu1/div/rem [9]),
        .I4(\alu1/div/dso_0 [9]),
        .O(\alu1/div/p_0_out [9]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_16_n_0),
        .I3(\alu0/div/rem [8]),
        .I4(\alu0/div/dso_0 [8]),
        .O(\alu0/div/p_0_out [8]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_16__0_n_0),
        .I3(\alu1/div/rem [8]),
        .I4(\alu1/div/dso_0 [8]),
        .O(\alu1/div/p_0_out [8]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_13
       (.I0(\alu0/div/den [11]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [11]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [11]),
        .O(add_out0_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_13__0
       (.I0(\alu1/div/den [11]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [11]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [11]),
        .O(add_out0_carry__1_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_14
       (.I0(\alu0/div/quo [10]),
        .I1(\alu0/div/dso_0 [10]),
        .I2(\alu0/div/den [10]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__1_i_14_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_14__0
       (.I0(\alu1/div/quo [10]),
        .I1(\alu1/div/dso_0 [10]),
        .I2(\alu1/div/den [10]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__1_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_15
       (.I0(\alu0/div/den [9]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [9]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [9]),
        .O(add_out0_carry__1_i_15_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__1_i_15__0
       (.I0(\alu1/div/den [9]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [9]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [9]),
        .O(add_out0_carry__1_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_16
       (.I0(\alu0/div/quo [8]),
        .I1(\alu0/div/dso_0 [8]),
        .I2(\alu0/div/den [8]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__1_i_16_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__1_i_16__0
       (.I0(\alu1/div/quo [8]),
        .I1(\alu1/div/dso_0 [8]),
        .I2(\alu1/div/den [8]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__1_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [11]),
        .O(add_out0_carry__1_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [10]),
        .O(add_out0_carry__1_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [10]),
        .O(add_out0_carry__1_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [9]),
        .O(add_out0_carry__1_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [9]),
        .O(add_out0_carry__1_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [8]),
        .O(add_out0_carry__1_i_4_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__1_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [8]),
        .O(add_out0_carry__1_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [11]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [11]),
        .O(add_out0_carry__1_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [11]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [11]),
        .O(add_out0_carry__1_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [10]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [10]),
        .O(add_out0_carry__1_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [10]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [10]),
        .O(add_out0_carry__1_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [9]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [9]),
        .O(add_out0_carry__1_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [9]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [9]),
        .O(add_out0_carry__1_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [8]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [8]),
        .O(add_out0_carry__1_i_8_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__1_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [8]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [8]),
        .O(add_out0_carry__1_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__1_i_13_n_0),
        .I3(\alu0/div/rem [11]),
        .I4(\alu0/div/dso_0 [11]),
        .O(\alu0/div/p_0_out [11]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__1_i_13__0_n_0),
        .I3(\alu1/div/rem [11]),
        .I4(\alu1/div/dso_0 [11]),
        .O(\alu1/div/p_0_out [11]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [15]),
        .O(add_out0_carry__2_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_14_n_0),
        .I3(\alu0/div/rem [14]),
        .I4(\alu0/div/dso_0 [14]),
        .O(\alu0/div/p_0_out [14]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_14__0_n_0),
        .I3(\alu1/div/rem [14]),
        .I4(\alu1/div/dso_0 [14]),
        .O(\alu1/div/p_0_out [14]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_15_n_0),
        .I3(\alu0/div/rem [13]),
        .I4(\alu0/div/dso_0 [13]),
        .O(\alu0/div/p_0_out [13]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_15__0_n_0),
        .I3(\alu1/div/rem [13]),
        .I4(\alu1/div/dso_0 [13]),
        .O(\alu1/div/p_0_out [13]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_16_n_0),
        .I3(\alu0/div/rem [12]),
        .I4(\alu0/div/dso_0 [12]),
        .O(\alu0/div/p_0_out [12]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_16__0_n_0),
        .I3(\alu1/div/rem [12]),
        .I4(\alu1/div/dso_0 [12]),
        .O(\alu1/div/p_0_out [12]));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__2_i_13
       (.I0(\alu0/div/den [15]),
        .I1(\alu0/div/quo [15]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [15]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__2_i_13_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__2_i_13__0
       (.I0(\alu1/div/den [15]),
        .I1(\alu1/div/quo [15]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [15]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__2_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__2_i_14
       (.I0(\alu0/div/quo [14]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [14]),
        .I4(\alu0/div/den [14]),
        .O(add_out0_carry__2_i_14_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__2_i_14__0
       (.I0(\alu1/div/quo [14]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [14]),
        .I4(\alu1/div/den [14]),
        .O(add_out0_carry__2_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__2_i_15
       (.I0(\alu0/div/den [13]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [13]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [13]),
        .O(add_out0_carry__2_i_15_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__2_i_15__0
       (.I0(\alu1/div/den [13]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [13]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [13]),
        .O(add_out0_carry__2_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__2_i_16
       (.I0(\alu0/div/quo [12]),
        .I1(\alu0/div/dso_0 [12]),
        .I2(\alu0/div/den [12]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__2_i_16_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__2_i_16__0
       (.I0(\alu1/div/quo [12]),
        .I1(\alu1/div/dso_0 [12]),
        .I2(\alu1/div/den [12]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__2_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [15]),
        .O(add_out0_carry__2_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [14]),
        .O(add_out0_carry__2_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [14]),
        .O(add_out0_carry__2_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [13]),
        .O(add_out0_carry__2_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [13]),
        .O(add_out0_carry__2_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [12]),
        .O(add_out0_carry__2_i_4_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__2_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [12]),
        .O(add_out0_carry__2_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [15]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [15]),
        .O(add_out0_carry__2_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [15]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [15]),
        .O(add_out0_carry__2_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [14]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [14]),
        .O(add_out0_carry__2_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [14]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [14]),
        .O(add_out0_carry__2_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [13]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [13]),
        .O(add_out0_carry__2_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [13]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [13]),
        .O(add_out0_carry__2_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [12]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [12]),
        .O(add_out0_carry__2_i_8_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__2_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [12]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [12]),
        .O(add_out0_carry__2_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__2_i_13_n_0),
        .I3(\alu0/div/rem [15]),
        .I4(\alu0/div/dso_0 [15]),
        .O(\alu0/div/p_0_out [15]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__2_i_13__0_n_0),
        .I3(\alu1/div/rem [15]),
        .I4(\alu1/div/dso_0 [15]),
        .O(\alu1/div/p_0_out [15]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [19]),
        .O(add_out0_carry__3_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_14_n_0),
        .I3(\alu0/div/rem [18]),
        .I4(\alu0/div/dso_0 [18]),
        .O(\alu0/div/p_0_out [18]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_14__0_n_0),
        .I3(\alu1/div/rem [18]),
        .I4(\alu1/div/dso_0 [18]),
        .O(\alu1/div/p_0_out [18]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_15_n_0),
        .I3(\alu0/div/rem [17]),
        .I4(\alu0/div/dso_0 [17]),
        .O(\alu0/div/p_0_out [17]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_15__0_n_0),
        .I3(\alu1/div/rem [17]),
        .I4(\alu1/div/dso_0 [17]),
        .O(\alu1/div/p_0_out [17]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_16_n_0),
        .I3(\alu0/div/rem [16]),
        .I4(\alu0/div/dso_0 [16]),
        .O(\alu0/div/p_0_out [16]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_16__0_n_0),
        .I3(\alu1/div/rem [16]),
        .I4(\alu1/div/dso_0 [16]),
        .O(\alu1/div/p_0_out [16]));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_13
       (.I0(\alu0/div/den [19]),
        .I1(\alu0/div/quo [19]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [19]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__3_i_13_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_13__0
       (.I0(\alu1/div/den [19]),
        .I1(\alu1/div/quo [19]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [19]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__3_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_14
       (.I0(\alu0/div/den [18]),
        .I1(\alu0/div/quo [18]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [18]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__3_i_14_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__3_i_14__0
       (.I0(\alu1/div/den [18]),
        .I1(\alu1/div/quo [18]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [18]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__3_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__3_i_15
       (.I0(\alu0/div/quo [17]),
        .I1(\alu0/div/dso_0 [17]),
        .I2(\alu0/div/den [17]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry__3_i_15_n_0));
  LUT5 #(
    .INIT(32'h0F550033)) 
    add_out0_carry__3_i_15__0
       (.I0(\alu1/div/quo [17]),
        .I1(\alu1/div/dso_0 [17]),
        .I2(\alu1/div/den [17]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry__3_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__3_i_16
       (.I0(\alu0/div/quo [16]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [16]),
        .I4(\alu0/div/den [16]),
        .O(add_out0_carry__3_i_16_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__3_i_16__0
       (.I0(\alu1/div/quo [16]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [16]),
        .I4(\alu1/div/den [16]),
        .O(add_out0_carry__3_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [19]),
        .O(add_out0_carry__3_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [18]),
        .O(add_out0_carry__3_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [18]),
        .O(add_out0_carry__3_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [17]),
        .O(add_out0_carry__3_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [17]),
        .O(add_out0_carry__3_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [16]),
        .O(add_out0_carry__3_i_4_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__3_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [16]),
        .O(add_out0_carry__3_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [19]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [19]),
        .O(add_out0_carry__3_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [19]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [19]),
        .O(add_out0_carry__3_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [18]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [18]),
        .O(add_out0_carry__3_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [18]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [18]),
        .O(add_out0_carry__3_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [17]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [17]),
        .O(add_out0_carry__3_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [17]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [17]),
        .O(add_out0_carry__3_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [16]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [16]),
        .O(add_out0_carry__3_i_8_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__3_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [16]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [16]),
        .O(add_out0_carry__3_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__3_i_13_n_0),
        .I3(\alu0/div/rem [19]),
        .I4(\alu0/div/dso_0 [19]),
        .O(\alu0/div/p_0_out [19]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__3_i_13__0_n_0),
        .I3(\alu1/div/rem [19]),
        .I4(\alu1/div/dso_0 [19]),
        .O(\alu1/div/p_0_out [19]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [23]),
        .O(add_out0_carry__4_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_14_n_0),
        .I3(\alu0/div/rem [22]),
        .I4(\alu0/div/dso_0 [22]),
        .O(\alu0/div/p_0_out [22]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_14__0_n_0),
        .I3(\alu1/div/rem [22]),
        .I4(\alu1/div/dso_0 [22]),
        .O(\alu1/div/p_0_out [22]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_15_n_0),
        .I3(\alu0/div/rem [21]),
        .I4(\alu0/div/dso_0 [21]),
        .O(\alu0/div/p_0_out [21]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_15__0_n_0),
        .I3(\alu1/div/rem [21]),
        .I4(\alu1/div/dso_0 [21]),
        .O(\alu1/div/p_0_out [21]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_16_n_0),
        .I3(\alu0/div/rem [20]),
        .I4(\alu0/div/dso_0 [20]),
        .O(\alu0/div/p_0_out [20]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_16__0_n_0),
        .I3(\alu1/div/rem [20]),
        .I4(\alu1/div/dso_0 [20]),
        .O(\alu1/div/p_0_out [20]));
  LUT5 #(
    .INIT(32'h0131C1F1)) 
    add_out0_carry__4_i_13
       (.I0(\alu0/div/dso_0 [23]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/quo [23]),
        .I4(\alu0/div/den [23]),
        .O(add_out0_carry__4_i_13_n_0));
  LUT5 #(
    .INIT(32'h0131C1F1)) 
    add_out0_carry__4_i_13__0
       (.I0(\alu1/div/dso_0 [23]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/quo [23]),
        .I4(\alu1/div/den [23]),
        .O(add_out0_carry__4_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_14
       (.I0(\alu0/div/quo [22]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [22]),
        .I4(\alu0/div/den [22]),
        .O(add_out0_carry__4_i_14_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_14__0
       (.I0(\alu1/div/quo [22]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [22]),
        .I4(\alu1/div/den [22]),
        .O(add_out0_carry__4_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_15
       (.I0(\alu0/div/quo [21]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [21]),
        .I4(\alu0/div/den [21]),
        .O(add_out0_carry__4_i_15_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__4_i_15__0
       (.I0(\alu1/div/quo [21]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [21]),
        .I4(\alu1/div/den [21]),
        .O(add_out0_carry__4_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__4_i_16
       (.I0(\alu0/div/den [20]),
        .I1(\alu0/div/quo [20]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [20]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry__4_i_16_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry__4_i_16__0
       (.I0(\alu1/div/den [20]),
        .I1(\alu1/div/quo [20]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [20]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry__4_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [23]),
        .O(add_out0_carry__4_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [22]),
        .O(add_out0_carry__4_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [22]),
        .O(add_out0_carry__4_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [21]),
        .O(add_out0_carry__4_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [21]),
        .O(add_out0_carry__4_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [20]),
        .O(add_out0_carry__4_i_4_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__4_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [20]),
        .O(add_out0_carry__4_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [23]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [23]),
        .O(add_out0_carry__4_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [23]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [23]),
        .O(add_out0_carry__4_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [22]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [22]),
        .O(add_out0_carry__4_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [22]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [22]),
        .O(add_out0_carry__4_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [21]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [21]),
        .O(add_out0_carry__4_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [21]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [21]),
        .O(add_out0_carry__4_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [20]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [20]),
        .O(add_out0_carry__4_i_8_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__4_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [20]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [20]),
        .O(add_out0_carry__4_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__4_i_13_n_0),
        .I3(\alu0/div/rem [23]),
        .I4(\alu0/div/dso_0 [23]),
        .O(\alu0/div/p_0_out [23]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__4_i_13__0_n_0),
        .I3(\alu1/div/rem [23]),
        .I4(\alu1/div/dso_0 [23]),
        .O(\alu1/div/p_0_out [23]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [27]),
        .O(add_out0_carry__5_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_14_n_0),
        .I3(\alu0/div/rem [26]),
        .I4(\alu0/div/dso_0 [26]),
        .O(\alu0/div/p_0_out [26]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_14__0_n_0),
        .I3(\alu1/div/rem [26]),
        .I4(\alu1/div/dso_0 [26]),
        .O(\alu1/div/p_0_out [26]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_15_n_0),
        .I3(\alu0/div/rem [25]),
        .I4(\alu0/div/dso_0 [25]),
        .O(\alu0/div/p_0_out [25]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_15__0_n_0),
        .I3(\alu1/div/rem [25]),
        .I4(\alu1/div/dso_0 [25]),
        .O(\alu1/div/p_0_out [25]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_16_n_0),
        .I3(\alu0/div/rem [24]),
        .I4(\alu0/div/dso_0 [24]),
        .O(\alu0/div/p_0_out [24]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_16__0_n_0),
        .I3(\alu1/div/rem [24]),
        .I4(\alu1/div/dso_0 [24]),
        .O(\alu1/div/p_0_out [24]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_13
       (.I0(\alu0/div/den [27]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [27]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [27]),
        .O(add_out0_carry__5_i_13_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_13__0
       (.I0(\alu1/div/den [27]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [27]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [27]),
        .O(add_out0_carry__5_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_14
       (.I0(\alu0/div/den [26]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [26]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [26]),
        .O(add_out0_carry__5_i_14_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_14__0
       (.I0(\alu1/div/den [26]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [26]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [26]),
        .O(add_out0_carry__5_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_15
       (.I0(\alu0/div/den [25]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [25]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [25]),
        .O(add_out0_carry__5_i_15_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__5_i_15__0
       (.I0(\alu1/div/den [25]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [25]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [25]),
        .O(add_out0_carry__5_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__5_i_16
       (.I0(\alu0/div/quo [24]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [24]),
        .I4(\alu0/div/den [24]),
        .O(add_out0_carry__5_i_16_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__5_i_16__0
       (.I0(\alu1/div/quo [24]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [24]),
        .I4(\alu1/div/den [24]),
        .O(add_out0_carry__5_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [27]),
        .O(add_out0_carry__5_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [26]),
        .O(add_out0_carry__5_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [26]),
        .O(add_out0_carry__5_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [25]),
        .O(add_out0_carry__5_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [25]),
        .O(add_out0_carry__5_i_3__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_4
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [24]),
        .O(add_out0_carry__5_i_4_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__5_i_4__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [24]),
        .O(add_out0_carry__5_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [27]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [27]),
        .O(add_out0_carry__5_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [27]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [27]),
        .O(add_out0_carry__5_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [26]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [26]),
        .O(add_out0_carry__5_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [26]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [26]),
        .O(add_out0_carry__5_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [25]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [25]),
        .O(add_out0_carry__5_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [25]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [25]),
        .O(add_out0_carry__5_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [24]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [24]),
        .O(add_out0_carry__5_i_8_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__5_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [24]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [24]),
        .O(add_out0_carry__5_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__5_i_13_n_0),
        .I3(\alu0/div/rem [27]),
        .I4(\alu0/div/dso_0 [27]),
        .O(\alu0/div/p_0_out [27]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__5_i_13__0_n_0),
        .I3(\alu1/div/rem [27]),
        .I4(\alu1/div/dso_0 [27]),
        .O(\alu1/div/p_0_out [27]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [30]),
        .O(add_out0_carry__6_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__6_i_13_n_0),
        .I3(\alu0/div/rem [28]),
        .I4(\alu0/div/dso_0 [28]),
        .O(\alu0/div/p_0_out [28]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__6_i_13__0_n_0),
        .I3(\alu1/div/rem [28]),
        .I4(\alu1/div/dso_0 [28]),
        .O(\alu1/div/p_0_out [28]));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_11
       (.I0(\alu0/div/den [30]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo__0 [30]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [30]),
        .O(add_out0_carry__6_i_11_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_11__0
       (.I0(\alu1/div/den [30]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo__0 [30]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [30]),
        .O(add_out0_carry__6_i_11__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__6_i_12
       (.I0(\alu0/div/quo__0 [29]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [29]),
        .I4(\alu0/div/den [29]),
        .O(add_out0_carry__6_i_12_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry__6_i_12__0
       (.I0(\alu1/div/quo__0 [29]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [29]),
        .I4(\alu1/div/den [29]),
        .O(add_out0_carry__6_i_12__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_13
       (.I0(\alu0/div/den [28]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo__0 [28]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [28]),
        .O(add_out0_carry__6_i_13_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry__6_i_13__0
       (.I0(\alu1/div/den [28]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo__0 [28]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [28]),
        .O(add_out0_carry__6_i_13__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [30]),
        .O(add_out0_carry__6_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [29]),
        .O(add_out0_carry__6_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [29]),
        .O(add_out0_carry__6_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [28]),
        .O(add_out0_carry__6_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry__6_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [28]),
        .O(add_out0_carry__6_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h003300555ABB0F5F)) 
    add_out0_carry__6_i_4
       (.I0(\alu0/div/dso_0 [31]),
        .I1(\alu0/div/quo__0 [31]),
        .I2(\alu0/div/rem [31]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\dso[31]_i_3_n_0 ),
        .I5(\rem[31]_i_3_n_0 ),
        .O(add_out0_carry__6_i_4_n_0));
  LUT6 #(
    .INIT(64'h003300555ABB0F5F)) 
    add_out0_carry__6_i_4__0
       (.I0(\alu1/div/dso_0 [31]),
        .I1(\alu1/div/quo__0 [31]),
        .I2(\alu1/div/rem [31]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\dso[31]_i_3__0_n_0 ),
        .I5(\rem[31]_i_3__0_n_0 ),
        .O(add_out0_carry__6_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [30]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [30]),
        .O(add_out0_carry__6_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [30]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [30]),
        .O(add_out0_carry__6_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [29]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [29]),
        .O(add_out0_carry__6_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [29]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [29]),
        .O(add_out0_carry__6_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [28]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [28]),
        .O(add_out0_carry__6_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry__6_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [28]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [28]),
        .O(add_out0_carry__6_i_7__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_8
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__6_i_11_n_0),
        .I3(\alu0/div/rem [30]),
        .I4(\alu0/div/dso_0 [30]),
        .O(\alu0/div/p_0_out [30]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_8__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__6_i_11__0_n_0),
        .I3(\alu1/div/rem [30]),
        .I4(\alu1/div/dso_0 [30]),
        .O(\alu1/div/p_0_out [30]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry__6_i_12_n_0),
        .I3(\alu0/div/rem [29]),
        .I4(\alu0/div/dso_0 [29]),
        .O(\alu0/div/p_0_out [29]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry__6_i_12__0_n_0),
        .I3(\alu1/div/rem [29]),
        .I4(\alu1/div/dso_0 [29]),
        .O(\alu1/div/p_0_out [29]));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_1
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [3]),
        .O(add_out0_carry_i_1_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_14_n_0),
        .I3(\alu0/div/rem [2]),
        .I4(\alu0/div/dso_0 [2]),
        .O(\alu0/div/p_0_out [2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_10__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_14__0_n_0),
        .I3(\alu1/div/rem [2]),
        .I4(\alu1/div/dso_0 [2]),
        .O(\alu1/div/p_0_out [2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_15_n_0),
        .I3(\alu0/div/rem [1]),
        .I4(\alu0/div/dso_0 [1]),
        .O(\alu0/div/p_0_out [1]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_11__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_15__0_n_0),
        .I3(\alu1/div/rem [1]),
        .I4(\alu1/div/dso_0 [1]),
        .O(\alu1/div/p_0_out [1]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_16_n_0),
        .I3(\alu0/div/rem [0]),
        .I4(\alu0/div/dso_0 [0]),
        .O(\alu0/div/p_0_out [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_12__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_16__0_n_0),
        .I3(\alu1/div/rem [0]),
        .I4(\alu1/div/dso_0 [0]),
        .O(\alu1/div/p_0_out [0]));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_13
       (.I0(\alu0/div/quo [3]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [3]),
        .I4(\alu0/div/den [3]),
        .O(add_out0_carry_i_13_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_13__0
       (.I0(\alu1/div/quo [3]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [3]),
        .I4(\alu1/div/den [3]),
        .O(add_out0_carry_i_13__0_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry_i_14
       (.I0(\alu0/div/den [2]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/quo [2]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [2]),
        .O(add_out0_carry_i_14_n_0));
  LUT5 #(
    .INIT(32'h47004733)) 
    add_out0_carry_i_14__0
       (.I0(\alu1/div/den [2]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/quo [2]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [2]),
        .O(add_out0_carry_i_14__0_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_15
       (.I0(\alu0/div/quo [1]),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [1]),
        .I4(\alu0/div/den [1]),
        .O(add_out0_carry_i_15_n_0));
  LUT5 #(
    .INIT(32'h1013D0D3)) 
    add_out0_carry_i_15__0
       (.I0(\alu1/div/quo [1]),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [1]),
        .I4(\alu1/div/den [1]),
        .O(add_out0_carry_i_15__0_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry_i_16
       (.I0(\alu0/div/den [0]),
        .I1(\alu0/div/quo [0]),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(\alu0/div/dso_0 [0]),
        .I4(\dso[31]_i_4_n_0 ),
        .O(add_out0_carry_i_16_n_0));
  LUT5 #(
    .INIT(32'h5050303F)) 
    add_out0_carry_i_16__0
       (.I0(\alu1/div/den [0]),
        .I1(\alu1/div/quo [0]),
        .I2(\dso[31]_i_3__0_n_0 ),
        .I3(\alu1/div/dso_0 [0]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .O(add_out0_carry_i_16__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_1__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [3]),
        .O(add_out0_carry_i_1__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_2
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [2]),
        .O(add_out0_carry_i_2_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_2__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [2]),
        .O(add_out0_carry_i_2__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_3
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [1]),
        .O(add_out0_carry_i_3_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    add_out0_carry_i_3__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [1]),
        .O(add_out0_carry_i_3__0_n_0));
  LUT4 #(
    .INIT(16'hFC77)) 
    add_out0_carry_i_4
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [0]),
        .I3(\dso[31]_i_3_n_0 ),
        .O(add_out0_carry_i_4_n_0));
  LUT4 #(
    .INIT(16'hFC77)) 
    add_out0_carry_i_4__0
       (.I0(\dso[31]_i_4__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [0]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .O(add_out0_carry_i_4__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_5
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [3]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [3]),
        .O(add_out0_carry_i_5_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_5__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [3]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [3]),
        .O(add_out0_carry_i_5__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_6
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [2]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [2]),
        .O(add_out0_carry_i_6_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_6__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [2]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [2]),
        .O(add_out0_carry_i_6__0_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_7
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [1]),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [1]),
        .O(add_out0_carry_i_7_n_0));
  LUT5 #(
    .INIT(32'hDFFF2000)) 
    add_out0_carry_i_7__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [1]),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [1]),
        .O(add_out0_carry_i_7__0_n_0));
  LUT5 #(
    .INIT(32'h5202ADFD)) 
    add_out0_carry_i_8
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\alu0/div/rem [0]),
        .I2(\rem[31]_i_3_n_0 ),
        .I3(\dso[31]_i_4_n_0 ),
        .I4(\alu0/div/p_0_out [0]),
        .O(add_out0_carry_i_8_n_0));
  LUT5 #(
    .INIT(32'h5202ADFD)) 
    add_out0_carry_i_8__0
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\alu1/div/rem [0]),
        .I2(\rem[31]_i_3__0_n_0 ),
        .I3(\dso[31]_i_4__0_n_0 ),
        .I4(\alu1/div/p_0_out [0]),
        .O(add_out0_carry_i_8__0_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_13_n_0),
        .I3(\alu0/div/rem [3]),
        .I4(\alu0/div/dso_0 [3]),
        .O(\alu0/div/p_0_out [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_9__0
       (.I0(\rem[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(add_out0_carry_i_13__0_n_0),
        .I3(\alu1/div/rem [3]),
        .I4(\alu1/div/dso_0 [3]),
        .O(\alu1/div/p_0_out [3]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry 
       (.CI(\<const0> ),
        .CO({\alu0/div/dadd/add_out0_carry_n_0 ,\alu0/div/dadd/add_out0_carry_n_1 ,\alu0/div/dadd/add_out0_carry_n_2 ,\alu0/div/dadd/add_out0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry_i_1_n_0,add_out0_carry_i_2_n_0,add_out0_carry_i_3_n_0,add_out0_carry_i_4_n_0}),
        .O(\alu0/div/add_out [3:0]),
        .S({add_out0_carry_i_5_n_0,add_out0_carry_i_6_n_0,add_out0_carry_i_7_n_0,add_out0_carry_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry__0 
       (.CI(\alu0/div/dadd/add_out0_carry_n_0 ),
        .CO({\alu0/div/dadd/add_out0_carry__0_n_0 ,\alu0/div/dadd/add_out0_carry__0_n_1 ,\alu0/div/dadd/add_out0_carry__0_n_2 ,\alu0/div/dadd/add_out0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__0_i_1_n_0,add_out0_carry__0_i_2_n_0,add_out0_carry__0_i_3_n_0,add_out0_carry__0_i_4_n_0}),
        .O(\alu0/div/add_out [7:4]),
        .S({add_out0_carry__0_i_5_n_0,add_out0_carry__0_i_6_n_0,add_out0_carry__0_i_7_n_0,add_out0_carry__0_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry__1 
       (.CI(\alu0/div/dadd/add_out0_carry__0_n_0 ),
        .CO({\alu0/div/dadd/add_out0_carry__1_n_0 ,\alu0/div/dadd/add_out0_carry__1_n_1 ,\alu0/div/dadd/add_out0_carry__1_n_2 ,\alu0/div/dadd/add_out0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__1_i_1_n_0,add_out0_carry__1_i_2_n_0,add_out0_carry__1_i_3_n_0,add_out0_carry__1_i_4_n_0}),
        .O(\alu0/div/add_out [11:8]),
        .S({add_out0_carry__1_i_5_n_0,add_out0_carry__1_i_6_n_0,add_out0_carry__1_i_7_n_0,add_out0_carry__1_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry__2 
       (.CI(\alu0/div/dadd/add_out0_carry__1_n_0 ),
        .CO({\alu0/div/dadd/add_out0_carry__2_n_0 ,\alu0/div/dadd/add_out0_carry__2_n_1 ,\alu0/div/dadd/add_out0_carry__2_n_2 ,\alu0/div/dadd/add_out0_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__2_i_1_n_0,add_out0_carry__2_i_2_n_0,add_out0_carry__2_i_3_n_0,add_out0_carry__2_i_4_n_0}),
        .O(\alu0/div/add_out [15:12]),
        .S({add_out0_carry__2_i_5_n_0,add_out0_carry__2_i_6_n_0,add_out0_carry__2_i_7_n_0,add_out0_carry__2_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry__3 
       (.CI(\alu0/div/dadd/add_out0_carry__2_n_0 ),
        .CO({\alu0/div/dadd/add_out0_carry__3_n_0 ,\alu0/div/dadd/add_out0_carry__3_n_1 ,\alu0/div/dadd/add_out0_carry__3_n_2 ,\alu0/div/dadd/add_out0_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__3_i_1_n_0,add_out0_carry__3_i_2_n_0,add_out0_carry__3_i_3_n_0,add_out0_carry__3_i_4_n_0}),
        .O(\alu0/div/add_out [19:16]),
        .S({add_out0_carry__3_i_5_n_0,add_out0_carry__3_i_6_n_0,add_out0_carry__3_i_7_n_0,add_out0_carry__3_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry__4 
       (.CI(\alu0/div/dadd/add_out0_carry__3_n_0 ),
        .CO({\alu0/div/dadd/add_out0_carry__4_n_0 ,\alu0/div/dadd/add_out0_carry__4_n_1 ,\alu0/div/dadd/add_out0_carry__4_n_2 ,\alu0/div/dadd/add_out0_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__4_i_1_n_0,add_out0_carry__4_i_2_n_0,add_out0_carry__4_i_3_n_0,add_out0_carry__4_i_4_n_0}),
        .O(\alu0/div/add_out [23:20]),
        .S({add_out0_carry__4_i_5_n_0,add_out0_carry__4_i_6_n_0,add_out0_carry__4_i_7_n_0,add_out0_carry__4_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry__5 
       (.CI(\alu0/div/dadd/add_out0_carry__4_n_0 ),
        .CO({\alu0/div/dadd/add_out0_carry__5_n_0 ,\alu0/div/dadd/add_out0_carry__5_n_1 ,\alu0/div/dadd/add_out0_carry__5_n_2 ,\alu0/div/dadd/add_out0_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__5_i_1_n_0,add_out0_carry__5_i_2_n_0,add_out0_carry__5_i_3_n_0,add_out0_carry__5_i_4_n_0}),
        .O(\alu0/div/add_out [27:24]),
        .S({add_out0_carry__5_i_5_n_0,add_out0_carry__5_i_6_n_0,add_out0_carry__5_i_7_n_0,add_out0_carry__5_i_8_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/dadd/add_out0_carry__6 
       (.CI(\alu0/div/dadd/add_out0_carry__5_n_0 ),
        .CO({\alu0/div/dadd/add_out0_carry__6_n_1 ,\alu0/div/dadd/add_out0_carry__6_n_2 ,\alu0/div/dadd/add_out0_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,add_out0_carry__6_i_1_n_0,add_out0_carry__6_i_2_n_0,add_out0_carry__6_i_3_n_0}),
        .O(\alu0/div/add_out [31:28]),
        .S({add_out0_carry__6_i_4_n_0,add_out0_carry__6_i_5_n_0,add_out0_carry__6_i_6_n_0,add_out0_carry__6_i_7_n_0}));
  FDRE \alu0/div/dctl/dctl_long_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/div/dctl_long ),
        .Q(\alu0/div/dctl/dctl_long_f ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/dctl_sign_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/div/dctl/dctl_sign ),
        .Q(\alu0/div/dctl/dctl_sign_f ),
        .R(\alu1/div/p_0_in__0 ));
  FDSE \alu0/div/dctl/div_crdy_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(div_crdy_i_1_n_0),
        .Q(div_crdy0),
        .S(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/fsm/chg_quo_sgn_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_quo_sgn_i_1_n_0),
        .Q(\alu0/div/chg_quo_sgn ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/fsm/chg_rem_sgn_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_rem_sgn_i_1_n_0),
        .Q(\alu0/div/chg_rem_sgn ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/fsm/dctl_stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/div/dctl/fsm/dctl_next [0]),
        .Q(\alu0/div/dctl_stat [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/fsm/dctl_stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/div/dctl/fsm/dctl_next [1]),
        .Q(\alu0/div/dctl_stat [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/fsm/dctl_stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/div/dctl/fsm/dctl_next [2]),
        .Q(\alu0/div/dctl_stat [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/fsm/dctl_stat_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/div/dctl/fsm/dctl_next [3]),
        .Q(\alu0/div/dctl_stat [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/dctl/fsm/fdiv_rem_msb_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/div/p_0_in0 ),
        .Q(\alu0/div/fdiv_rem_msb_f ),
        .R(\alu1/div/p_0_in__0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry 
       (.CI(\<const0> ),
        .CO({\alu0/div/fdiv/rem0_carry_n_0 ,\alu0/div/fdiv/rem0_carry_n_1 ,\alu0/div/fdiv/rem0_carry_n_2 ,\alu0/div/fdiv/rem0_carry_n_3 }),
        .CYINIT(rem0_carry_i_1_n_0),
        .DI({\alu0/div/rem1__0 [3:1],\alu0/div/den [28]}),
        .O(\alu0/div/fdiv_rem [3:0]),
        .S({rem0_carry_i_2_n_0,rem0_carry_i_3_n_0,rem0_carry_i_4_n_0,rem0_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__0 
       (.CI(\alu0/div/fdiv/rem0_carry_n_0 ),
        .CO({\alu0/div/fdiv/rem0_carry__0_n_0 ,\alu0/div/fdiv/rem0_carry__0_n_1 ,\alu0/div/fdiv/rem0_carry__0_n_2 ,\alu0/div/fdiv/rem0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem1__0 [7:4]),
        .O(\alu0/div/fdiv_rem [7:4]),
        .S({rem0_carry__0_i_1_n_0,rem0_carry__0_i_2_n_0,rem0_carry__0_i_3_n_0,rem0_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__1 
       (.CI(\alu0/div/fdiv/rem0_carry__0_n_0 ),
        .CO({\alu0/div/fdiv/rem0_carry__1_n_0 ,\alu0/div/fdiv/rem0_carry__1_n_1 ,\alu0/div/fdiv/rem0_carry__1_n_2 ,\alu0/div/fdiv/rem0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem1__0 [11:8]),
        .O(\alu0/div/fdiv_rem [11:8]),
        .S({rem0_carry__1_i_1_n_0,rem0_carry__1_i_2_n_0,rem0_carry__1_i_3_n_0,rem0_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__2 
       (.CI(\alu0/div/fdiv/rem0_carry__1_n_0 ),
        .CO({\alu0/div/fdiv/rem0_carry__2_n_0 ,\alu0/div/fdiv/rem0_carry__2_n_1 ,\alu0/div/fdiv/rem0_carry__2_n_2 ,\alu0/div/fdiv/rem0_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem1__0 [15:12]),
        .O(\alu0/div/fdiv_rem [15:12]),
        .S({rem0_carry__2_i_1_n_0,rem0_carry__2_i_2_n_0,rem0_carry__2_i_3_n_0,rem0_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__3 
       (.CI(\alu0/div/fdiv/rem0_carry__2_n_0 ),
        .CO({\alu0/div/fdiv/rem0_carry__3_n_0 ,\alu0/div/fdiv/rem0_carry__3_n_1 ,\alu0/div/fdiv/rem0_carry__3_n_2 ,\alu0/div/fdiv/rem0_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem1__0 [19:16]),
        .O(\alu0/div/fdiv_rem [19:16]),
        .S({rem0_carry__3_i_1_n_0,rem0_carry__3_i_2_n_0,rem0_carry__3_i_3_n_0,rem0_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__4 
       (.CI(\alu0/div/fdiv/rem0_carry__3_n_0 ),
        .CO({\alu0/div/fdiv/rem0_carry__4_n_0 ,\alu0/div/fdiv/rem0_carry__4_n_1 ,\alu0/div/fdiv/rem0_carry__4_n_2 ,\alu0/div/fdiv/rem0_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem1__0 [23:20]),
        .O(\alu0/div/fdiv_rem [23:20]),
        .S({rem0_carry__4_i_1_n_0,rem0_carry__4_i_2_n_0,rem0_carry__4_i_3_n_0,rem0_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__5 
       (.CI(\alu0/div/fdiv/rem0_carry__4_n_0 ),
        .CO({\alu0/div/fdiv/rem0_carry__5_n_0 ,\alu0/div/fdiv/rem0_carry__5_n_1 ,\alu0/div/fdiv/rem0_carry__5_n_2 ,\alu0/div/fdiv/rem0_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem1__0 [27:24]),
        .O(\alu0/div/fdiv_rem [27:24]),
        .S({rem0_carry__5_i_1_n_0,rem0_carry__5_i_2_n_0,rem0_carry__5_i_3_n_0,rem0_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__6 
       (.CI(\alu0/div/fdiv/rem0_carry__5_n_0 ),
        .CO({\alu0/div/fdiv/rem0_carry__6_n_0 ,\alu0/div/fdiv/rem0_carry__6_n_1 ,\alu0/div/fdiv/rem0_carry__6_n_2 ,\alu0/div/fdiv/rem0_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem1__0 [31:28]),
        .O(\alu0/div/fdiv_rem [31:28]),
        .S({rem0_carry__6_i_1_n_0,rem0_carry__6_i_2_n_0,rem0_carry__6_i_3_n_0,rem0_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem0_carry__7 
       (.CI(\alu0/div/fdiv/rem0_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu0/div/p_0_in0 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem0_carry__7_i_1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry 
       (.CI(\<const0> ),
        .CO({\alu0/div/fdiv/rem1_carry_n_0 ,\alu0/div/fdiv/rem1_carry_n_1 ,\alu0/div/fdiv/rem1_carry_n_2 ,\alu0/div/fdiv/rem1_carry_n_3 }),
        .CYINIT(rem1_carry_i_1_n_0),
        .DI({\alu0/div/rem2__0 [3:1],\alu0/div/den [29]}),
        .O(\alu0/div/rem1__0 [4:1]),
        .S({rem1_carry_i_2_n_0,rem1_carry_i_3_n_0,rem1_carry_i_4_n_0,rem1_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__0 
       (.CI(\alu0/div/fdiv/rem1_carry_n_0 ),
        .CO({\alu0/div/fdiv/rem1_carry__0_n_0 ,\alu0/div/fdiv/rem1_carry__0_n_1 ,\alu0/div/fdiv/rem1_carry__0_n_2 ,\alu0/div/fdiv/rem1_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem2__0 [7:4]),
        .O(\alu0/div/rem1__0 [8:5]),
        .S({rem1_carry__0_i_1_n_0,rem1_carry__0_i_2_n_0,rem1_carry__0_i_3_n_0,rem1_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__1 
       (.CI(\alu0/div/fdiv/rem1_carry__0_n_0 ),
        .CO({\alu0/div/fdiv/rem1_carry__1_n_0 ,\alu0/div/fdiv/rem1_carry__1_n_1 ,\alu0/div/fdiv/rem1_carry__1_n_2 ,\alu0/div/fdiv/rem1_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem2__0 [11:8]),
        .O(\alu0/div/rem1__0 [12:9]),
        .S({rem1_carry__1_i_1_n_0,rem1_carry__1_i_2_n_0,rem1_carry__1_i_3_n_0,rem1_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__2 
       (.CI(\alu0/div/fdiv/rem1_carry__1_n_0 ),
        .CO({\alu0/div/fdiv/rem1_carry__2_n_0 ,\alu0/div/fdiv/rem1_carry__2_n_1 ,\alu0/div/fdiv/rem1_carry__2_n_2 ,\alu0/div/fdiv/rem1_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem2__0 [15:12]),
        .O(\alu0/div/rem1__0 [16:13]),
        .S({rem1_carry__2_i_1_n_0,rem1_carry__2_i_2_n_0,rem1_carry__2_i_3_n_0,rem1_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__3 
       (.CI(\alu0/div/fdiv/rem1_carry__2_n_0 ),
        .CO({\alu0/div/fdiv/rem1_carry__3_n_0 ,\alu0/div/fdiv/rem1_carry__3_n_1 ,\alu0/div/fdiv/rem1_carry__3_n_2 ,\alu0/div/fdiv/rem1_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem2__0 [19:16]),
        .O(\alu0/div/rem1__0 [20:17]),
        .S({rem1_carry__3_i_1_n_0,rem1_carry__3_i_2_n_0,rem1_carry__3_i_3_n_0,rem1_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__4 
       (.CI(\alu0/div/fdiv/rem1_carry__3_n_0 ),
        .CO({\alu0/div/fdiv/rem1_carry__4_n_0 ,\alu0/div/fdiv/rem1_carry__4_n_1 ,\alu0/div/fdiv/rem1_carry__4_n_2 ,\alu0/div/fdiv/rem1_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem2__0 [23:20]),
        .O(\alu0/div/rem1__0 [24:21]),
        .S({rem1_carry__4_i_1_n_0,rem1_carry__4_i_2_n_0,rem1_carry__4_i_3_n_0,rem1_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__5 
       (.CI(\alu0/div/fdiv/rem1_carry__4_n_0 ),
        .CO({\alu0/div/fdiv/rem1_carry__5_n_0 ,\alu0/div/fdiv/rem1_carry__5_n_1 ,\alu0/div/fdiv/rem1_carry__5_n_2 ,\alu0/div/fdiv/rem1_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem2__0 [27:24]),
        .O(\alu0/div/rem1__0 [28:25]),
        .S({rem1_carry__5_i_1_n_0,rem1_carry__5_i_2_n_0,rem1_carry__5_i_3_n_0,rem1_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__6 
       (.CI(\alu0/div/fdiv/rem1_carry__5_n_0 ),
        .CO({\alu0/div/fdiv/rem1_carry__6_n_0 ,\alu0/div/fdiv/rem1_carry__6_n_1 ,\alu0/div/fdiv/rem1_carry__6_n_2 ,\alu0/div/fdiv/rem1_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem2__0 [31:28]),
        .O(\alu0/div/rem1__0 [32:29]),
        .S({rem1_carry__6_i_1_n_0,rem1_carry__6_i_2_n_0,rem1_carry__6_i_3_n_0,rem1_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem1_carry__7 
       (.CI(\alu0/div/fdiv/rem1_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu0/div/rem1 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem1_carry__7_i_1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry 
       (.CI(\<const0> ),
        .CO({\alu0/div/fdiv/rem2_carry_n_0 ,\alu0/div/fdiv/rem2_carry_n_1 ,\alu0/div/fdiv/rem2_carry_n_2 ,\alu0/div/fdiv/rem2_carry_n_3 }),
        .CYINIT(\alu0/div/fdiv/p_1_in3_in ),
        .DI({\alu0/div/rem3__0 [3:1],\alu0/div/den [30]}),
        .O(\alu0/div/rem2__0 [4:1]),
        .S({rem2_carry_i_2_n_0,rem2_carry_i_3_n_0,rem2_carry_i_4_n_0,rem2_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__0 
       (.CI(\alu0/div/fdiv/rem2_carry_n_0 ),
        .CO({\alu0/div/fdiv/rem2_carry__0_n_0 ,\alu0/div/fdiv/rem2_carry__0_n_1 ,\alu0/div/fdiv/rem2_carry__0_n_2 ,\alu0/div/fdiv/rem2_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem3__0 [7:4]),
        .O(\alu0/div/rem2__0 [8:5]),
        .S({rem2_carry__0_i_1_n_0,rem2_carry__0_i_2_n_0,rem2_carry__0_i_3_n_0,rem2_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__1 
       (.CI(\alu0/div/fdiv/rem2_carry__0_n_0 ),
        .CO({\alu0/div/fdiv/rem2_carry__1_n_0 ,\alu0/div/fdiv/rem2_carry__1_n_1 ,\alu0/div/fdiv/rem2_carry__1_n_2 ,\alu0/div/fdiv/rem2_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem3__0 [11:8]),
        .O(\alu0/div/rem2__0 [12:9]),
        .S({rem2_carry__1_i_1_n_0,rem2_carry__1_i_2_n_0,rem2_carry__1_i_3_n_0,rem2_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__2 
       (.CI(\alu0/div/fdiv/rem2_carry__1_n_0 ),
        .CO({\alu0/div/fdiv/rem2_carry__2_n_0 ,\alu0/div/fdiv/rem2_carry__2_n_1 ,\alu0/div/fdiv/rem2_carry__2_n_2 ,\alu0/div/fdiv/rem2_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem3__0 [15:12]),
        .O(\alu0/div/rem2__0 [16:13]),
        .S({rem2_carry__2_i_1_n_0,rem2_carry__2_i_2_n_0,rem2_carry__2_i_3_n_0,rem2_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__3 
       (.CI(\alu0/div/fdiv/rem2_carry__2_n_0 ),
        .CO({\alu0/div/fdiv/rem2_carry__3_n_0 ,\alu0/div/fdiv/rem2_carry__3_n_1 ,\alu0/div/fdiv/rem2_carry__3_n_2 ,\alu0/div/fdiv/rem2_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem3__0 [19:16]),
        .O(\alu0/div/rem2__0 [20:17]),
        .S({rem2_carry__3_i_1_n_0,rem2_carry__3_i_2_n_0,rem2_carry__3_i_3_n_0,rem2_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__4 
       (.CI(\alu0/div/fdiv/rem2_carry__3_n_0 ),
        .CO({\alu0/div/fdiv/rem2_carry__4_n_0 ,\alu0/div/fdiv/rem2_carry__4_n_1 ,\alu0/div/fdiv/rem2_carry__4_n_2 ,\alu0/div/fdiv/rem2_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem3__0 [23:20]),
        .O(\alu0/div/rem2__0 [24:21]),
        .S({rem2_carry__4_i_1_n_0,rem2_carry__4_i_2_n_0,rem2_carry__4_i_3_n_0,rem2_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__5 
       (.CI(\alu0/div/fdiv/rem2_carry__4_n_0 ),
        .CO({\alu0/div/fdiv/rem2_carry__5_n_0 ,\alu0/div/fdiv/rem2_carry__5_n_1 ,\alu0/div/fdiv/rem2_carry__5_n_2 ,\alu0/div/fdiv/rem2_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem3__0 [27:24]),
        .O(\alu0/div/rem2__0 [28:25]),
        .S({rem2_carry__5_i_1_n_0,rem2_carry__5_i_2_n_0,rem2_carry__5_i_3_n_0,rem2_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__6 
       (.CI(\alu0/div/fdiv/rem2_carry__5_n_0 ),
        .CO({\alu0/div/fdiv/rem2_carry__6_n_0 ,\alu0/div/fdiv/rem2_carry__6_n_1 ,\alu0/div/fdiv/rem2_carry__6_n_2 ,\alu0/div/fdiv/rem2_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/rem3__0 [31:28]),
        .O(\alu0/div/rem2__0 [32:29]),
        .S({rem2_carry__6_i_1_n_0,rem2_carry__6_i_2_n_0,rem2_carry__6_i_3_n_0,rem2_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem2_carry__7 
       (.CI(\alu0/div/fdiv/rem2_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu0/div/rem2 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem2_carry__7_i_1_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry 
       (.CI(\<const0> ),
        .CO({\alu0/div/fdiv/rem3_carry_n_0 ,\alu0/div/fdiv/rem3_carry_n_1 ,\alu0/div/fdiv/rem3_carry_n_2 ,\alu0/div/fdiv/rem3_carry_n_3 }),
        .CYINIT(\alu0/div/fdiv/p_1_in5_in ),
        .DI({\alu0/div/den [34:32],\alu0/div/den2 }),
        .O(\alu0/div/rem3__0 [4:1]),
        .S({rem3_carry_i_2_n_0,rem3_carry_i_3_n_0,rem3_carry_i_4_n_0,rem3_carry_i_5_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__0 
       (.CI(\alu0/div/fdiv/rem3_carry_n_0 ),
        .CO({\alu0/div/fdiv/rem3_carry__0_n_0 ,\alu0/div/fdiv/rem3_carry__0_n_1 ,\alu0/div/fdiv/rem3_carry__0_n_2 ,\alu0/div/fdiv/rem3_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/den [38:35]),
        .O(\alu0/div/rem3__0 [8:5]),
        .S({rem3_carry__0_i_1_n_0,rem3_carry__0_i_2_n_0,rem3_carry__0_i_3_n_0,rem3_carry__0_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__1 
       (.CI(\alu0/div/fdiv/rem3_carry__0_n_0 ),
        .CO({\alu0/div/fdiv/rem3_carry__1_n_0 ,\alu0/div/fdiv/rem3_carry__1_n_1 ,\alu0/div/fdiv/rem3_carry__1_n_2 ,\alu0/div/fdiv/rem3_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/den [42:39]),
        .O(\alu0/div/rem3__0 [12:9]),
        .S({rem3_carry__1_i_1_n_0,rem3_carry__1_i_2_n_0,rem3_carry__1_i_3_n_0,rem3_carry__1_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__2 
       (.CI(\alu0/div/fdiv/rem3_carry__1_n_0 ),
        .CO({\alu0/div/fdiv/rem3_carry__2_n_0 ,\alu0/div/fdiv/rem3_carry__2_n_1 ,\alu0/div/fdiv/rem3_carry__2_n_2 ,\alu0/div/fdiv/rem3_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/den [46:43]),
        .O(\alu0/div/rem3__0 [16:13]),
        .S({rem3_carry__2_i_1_n_0,rem3_carry__2_i_2_n_0,rem3_carry__2_i_3_n_0,rem3_carry__2_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__3 
       (.CI(\alu0/div/fdiv/rem3_carry__2_n_0 ),
        .CO({\alu0/div/fdiv/rem3_carry__3_n_0 ,\alu0/div/fdiv/rem3_carry__3_n_1 ,\alu0/div/fdiv/rem3_carry__3_n_2 ,\alu0/div/fdiv/rem3_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/den [50:47]),
        .O(\alu0/div/rem3__0 [20:17]),
        .S({rem3_carry__3_i_1_n_0,rem3_carry__3_i_2_n_0,rem3_carry__3_i_3_n_0,rem3_carry__3_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__4 
       (.CI(\alu0/div/fdiv/rem3_carry__3_n_0 ),
        .CO({\alu0/div/fdiv/rem3_carry__4_n_0 ,\alu0/div/fdiv/rem3_carry__4_n_1 ,\alu0/div/fdiv/rem3_carry__4_n_2 ,\alu0/div/fdiv/rem3_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/den [54:51]),
        .O(\alu0/div/rem3__0 [24:21]),
        .S({rem3_carry__4_i_1_n_0,rem3_carry__4_i_2_n_0,rem3_carry__4_i_3_n_0,rem3_carry__4_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__5 
       (.CI(\alu0/div/fdiv/rem3_carry__4_n_0 ),
        .CO({\alu0/div/fdiv/rem3_carry__5_n_0 ,\alu0/div/fdiv/rem3_carry__5_n_1 ,\alu0/div/fdiv/rem3_carry__5_n_2 ,\alu0/div/fdiv/rem3_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/den [58:55]),
        .O(\alu0/div/rem3__0 [28:25]),
        .S({rem3_carry__5_i_1_n_0,rem3_carry__5_i_2_n_0,rem3_carry__5_i_3_n_0,rem3_carry__5_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__6 
       (.CI(\alu0/div/fdiv/rem3_carry__5_n_0 ),
        .CO({\alu0/div/fdiv/rem3_carry__6_n_0 ,\alu0/div/fdiv/rem3_carry__6_n_1 ,\alu0/div/fdiv/rem3_carry__6_n_2 ,\alu0/div/fdiv/rem3_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu0/div/den [62:59]),
        .O(\alu0/div/rem3__0 [32:29]),
        .S({rem3_carry__6_i_1_n_0,rem3_carry__6_i_2_n_0,rem3_carry__6_i_3_n_0,rem3_carry__6_i_4_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu0/div/fdiv/rem3_carry__7 
       (.CI(\alu0/div/fdiv/rem3_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu0/div/rem3 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem3_carry__7_i_1_n_0}));
  FDRE \alu0/div/rden/remden_reg[0] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[0]_i_1_n_0 ),
        .Q(\alu0/div/den [0]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[10] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[10]_i_1_n_0 ),
        .Q(\alu0/div/den [10]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[11] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[11]_i_1_n_0 ),
        .Q(\alu0/div/den [11]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[12] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[12]_i_1_n_0 ),
        .Q(\alu0/div/den [12]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[13] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[13]_i_1_n_0 ),
        .Q(\alu0/div/den [13]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[14] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[14]_i_1_n_0 ),
        .Q(\alu0/div/den [14]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[15] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[15]_i_1_n_0 ),
        .Q(\alu0/div/den [15]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[16] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[16]_i_1_n_0 ),
        .Q(\alu0/div/den [16]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[17] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[17]_i_1_n_0 ),
        .Q(\alu0/div/den [17]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[18] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[18]_i_1_n_0 ),
        .Q(\alu0/div/den [18]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[19] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[19]_i_1_n_0 ),
        .Q(\alu0/div/den [19]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[1] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[1]_i_1_n_0 ),
        .Q(\alu0/div/den [1]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[20] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[20]_i_1_n_0 ),
        .Q(\alu0/div/den [20]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[21] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[21]_i_1_n_0 ),
        .Q(\alu0/div/den [21]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[22] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[22]_i_1_n_0 ),
        .Q(\alu0/div/den [22]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[23] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[23]_i_1_n_0 ),
        .Q(\alu0/div/den [23]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[24] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[24]_i_1_n_0 ),
        .Q(\alu0/div/den [24]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[25] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[25]_i_1_n_0 ),
        .Q(\alu0/div/den [25]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[26] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[26]_i_1_n_0 ),
        .Q(\alu0/div/den [26]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[27] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[27]_i_1_n_0 ),
        .Q(\alu0/div/den [27]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[28] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[28]_i_1_n_0 ),
        .Q(\alu0/div/den [28]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[29] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[29]_i_1_n_0 ),
        .Q(\alu0/div/den [29]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[2] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[2]_i_1_n_0 ),
        .Q(\alu0/div/den [2]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[30] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[30]_i_1_n_0 ),
        .Q(\alu0/div/den [30]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[31] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[31]_i_2_n_0 ),
        .Q(\alu0/div/den2 ),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[32] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[32]_i_1_n_0 ),
        .Q(\alu0/div/den [32]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[33] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[33]_i_1_n_0 ),
        .Q(\alu0/div/den [33]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[34] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[34]_i_1_n_0 ),
        .Q(\alu0/div/den [34]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[35] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[35]_i_1_n_0 ),
        .Q(\alu0/div/den [35]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[36] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[36]_i_1_n_0 ),
        .Q(\alu0/div/den [36]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[37] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[37]_i_1_n_0 ),
        .Q(\alu0/div/den [37]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[38] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[38]_i_1_n_0 ),
        .Q(\alu0/div/den [38]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[39] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[39]_i_1_n_0 ),
        .Q(\alu0/div/den [39]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[3] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[3]_i_1_n_0 ),
        .Q(\alu0/div/den [3]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[40] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[40]_i_1_n_0 ),
        .Q(\alu0/div/den [40]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[41] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[41]_i_1_n_0 ),
        .Q(\alu0/div/den [41]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[42] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[42]_i_1_n_0 ),
        .Q(\alu0/div/den [42]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[43] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[43]_i_1_n_0 ),
        .Q(\alu0/div/den [43]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[44] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[44]_i_1_n_0 ),
        .Q(\alu0/div/den [44]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[45] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[45]_i_1_n_0 ),
        .Q(\alu0/div/den [45]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[46] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[46]_i_1_n_0 ),
        .Q(\alu0/div/den [46]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[47] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[47]_i_1_n_0 ),
        .Q(\alu0/div/den [47]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[48] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[48]_i_1_n_0 ),
        .Q(\alu0/div/den [48]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[49] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[49]_i_1_n_0 ),
        .Q(\alu0/div/den [49]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[4] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[4]_i_1_n_0 ),
        .Q(\alu0/div/den [4]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[50] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[50]_i_1_n_0 ),
        .Q(\alu0/div/den [50]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[51] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[51]_i_1_n_0 ),
        .Q(\alu0/div/den [51]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[52] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[52]_i_1_n_0 ),
        .Q(\alu0/div/den [52]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[53] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[53]_i_1_n_0 ),
        .Q(\alu0/div/den [53]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[54] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[54]_i_1_n_0 ),
        .Q(\alu0/div/den [54]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[55] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[55]_i_1_n_0 ),
        .Q(\alu0/div/den [55]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[56] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[56]_i_1_n_0 ),
        .Q(\alu0/div/den [56]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[57] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[57]_i_1_n_0 ),
        .Q(\alu0/div/den [57]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[58] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[58]_i_1_n_0 ),
        .Q(\alu0/div/den [58]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[59] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[59]_i_1_n_0 ),
        .Q(\alu0/div/den [59]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[5] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[5]_i_1_n_0 ),
        .Q(\alu0/div/den [5]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[60] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[60]_i_1_n_0 ),
        .Q(\alu0/div/den [60]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[61] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[61]_i_1_n_0 ),
        .Q(\alu0/div/den [61]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[62] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[62]_i_1_n_0 ),
        .Q(\alu0/div/den [62]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[63] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[63]_i_1_n_0 ),
        .Q(\alu0/div/den [63]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[64] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[64]_i_3_n_0 ),
        .Q(\alu0/div/den [64]),
        .R(\remden[64]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[6] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[6]_i_1_n_0 ),
        .Q(\alu0/div/den [6]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[7] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[7]_i_1_n_0 ),
        .Q(\alu0/div/den [7]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[8] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[8]_i_1_n_0 ),
        .Q(\alu0/div/den [8]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rden/remden_reg[9] 
       (.C(clk),
        .CE(\remden[64]_i_2_n_0 ),
        .D(\remden[9]_i_1_n_0 ),
        .Q(\alu0/div/den [9]),
        .R(\remden[31]_i_1_n_0 ));
  FDRE \alu0/div/rdso/dso_reg[0] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_7 ),
        .Q(\alu0/div/dso_0 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[10] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_5 ),
        .Q(\alu0/div/dso_0 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[11] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_4 ),
        .Q(\alu0/div/dso_0 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[12] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_7 ),
        .Q(\alu0/div/dso_0 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[13] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_6 ),
        .Q(\alu0/div/dso_0 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[14] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_5 ),
        .Q(\alu0/div/dso_0 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[15] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[15]_i_1_n_4 ),
        .Q(\alu0/div/dso_0 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[16] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_7 ),
        .Q(\alu0/div/dso_0 [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[17] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_6 ),
        .Q(\alu0/div/dso_0 [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[18] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_5 ),
        .Q(\alu0/div/dso_0 [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[19] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[19]_i_1_n_4 ),
        .Q(\alu0/div/dso_0 [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[1] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_6 ),
        .Q(\alu0/div/dso_0 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[20] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_7 ),
        .Q(\alu0/div/dso_0 [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[21] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_6 ),
        .Q(\alu0/div/dso_0 [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[22] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_5 ),
        .Q(\alu0/div/dso_0 [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[23] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[23]_i_1_n_4 ),
        .Q(\alu0/div/dso_0 [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[24] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_7 ),
        .Q(\alu0/div/dso_0 [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[25] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_6 ),
        .Q(\alu0/div/dso_0 [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[26] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_5 ),
        .Q(\alu0/div/dso_0 [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[27] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[27]_i_1_n_4 ),
        .Q(\alu0/div/dso_0 [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[28] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_7 ),
        .Q(\alu0/div/dso_0 [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[29] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_6 ),
        .Q(\alu0/div/dso_0 [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[2] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_5 ),
        .Q(\alu0/div/dso_0 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[30] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_5 ),
        .Q(\alu0/div/dso_0 [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[31] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[31]_i_2_n_4 ),
        .Q(\alu0/div/dso_0 [31]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[3] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[3]_i_1_n_4 ),
        .Q(\alu0/div/dso_0 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[4] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_7 ),
        .Q(\alu0/div/dso_0 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[5] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_6 ),
        .Q(\alu0/div/dso_0 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[6] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_5 ),
        .Q(\alu0/div/dso_0 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[7] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[7]_i_1_n_4 ),
        .Q(\alu0/div/dso_0 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[8] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_7 ),
        .Q(\alu0/div/dso_0 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rdso/dso_reg[9] 
       (.C(clk),
        .CE(\dso[31]_i_1_n_0 ),
        .D(\dso_reg[11]_i_1_n_6 ),
        .Q(\alu0/div/dso_0 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[0] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [0]),
        .Q(\alu0/div/quo [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[10] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [10]),
        .Q(\alu0/div/quo [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[11] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [11]),
        .Q(\alu0/div/quo [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[12] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [12]),
        .Q(\alu0/div/quo [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[13] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [13]),
        .Q(\alu0/div/quo [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[14] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [14]),
        .Q(\alu0/div/quo [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[15] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [15]),
        .Q(\alu0/div/quo [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[16] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [16]),
        .Q(\alu0/div/quo [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[17] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [17]),
        .Q(\alu0/div/quo [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[18] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [18]),
        .Q(\alu0/div/quo [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[19] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [19]),
        .Q(\alu0/div/quo [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[1] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [1]),
        .Q(\alu0/div/quo [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[20] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [20]),
        .Q(\alu0/div/quo [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[21] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [21]),
        .Q(\alu0/div/quo [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[22] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [22]),
        .Q(\alu0/div/quo [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[23] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [23]),
        .Q(\alu0/div/quo [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[24] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [24]),
        .Q(\alu0/div/quo [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[25] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [25]),
        .Q(\alu0/div/quo [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[26] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [26]),
        .Q(\alu0/div/quo [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[27] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [27]),
        .Q(\alu0/div/quo [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[28] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [28]),
        .Q(\alu0/div/quo__0 [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[29] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [29]),
        .Q(\alu0/div/quo__0 [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[2] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [2]),
        .Q(\alu0/div/quo [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[30] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [30]),
        .Q(\alu0/div/quo__0 [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[31] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [31]),
        .Q(\alu0/div/quo__0 [31]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[3] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [3]),
        .Q(\alu0/div/quo [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[4] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [4]),
        .Q(\alu0/div/quo [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[5] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [5]),
        .Q(\alu0/div/quo [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[6] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [6]),
        .Q(\alu0/div/quo [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[7] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [7]),
        .Q(\alu0/div/quo [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[8] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [8]),
        .Q(\alu0/div/quo [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rquo/quo_reg[9] 
       (.C(clk),
        .CE(\quo[31]_i_1_n_0 ),
        .D(\alu0/div/p_2_in [9]),
        .Q(\alu0/div/quo [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[0] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_7 ),
        .Q(\alu0/div/rem [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[10] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_5 ),
        .Q(\alu0/div/rem [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[11] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_4 ),
        .Q(\alu0/div/rem [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[12] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_7 ),
        .Q(\alu0/div/rem [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[13] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_6 ),
        .Q(\alu0/div/rem [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[14] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_5 ),
        .Q(\alu0/div/rem [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[15] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[15]_i_1_n_4 ),
        .Q(\alu0/div/rem [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[16] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_7 ),
        .Q(\alu0/div/rem [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[17] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_6 ),
        .Q(\alu0/div/rem [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[18] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_5 ),
        .Q(\alu0/div/rem [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[19] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[19]_i_1_n_4 ),
        .Q(\alu0/div/rem [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[1] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_6 ),
        .Q(\alu0/div/rem [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[20] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_7 ),
        .Q(\alu0/div/rem [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[21] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_6 ),
        .Q(\alu0/div/rem [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[22] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_5 ),
        .Q(\alu0/div/rem [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[23] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[23]_i_1_n_4 ),
        .Q(\alu0/div/rem [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[24] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_7 ),
        .Q(\alu0/div/rem [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[25] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_6 ),
        .Q(\alu0/div/rem [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[26] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_5 ),
        .Q(\alu0/div/rem [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[27] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[27]_i_1_n_4 ),
        .Q(\alu0/div/rem [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[28] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_7 ),
        .Q(\alu0/div/rem [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[29] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_6 ),
        .Q(\alu0/div/rem [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[2] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_5 ),
        .Q(\alu0/div/rem [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[30] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_5 ),
        .Q(\alu0/div/rem [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[31] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[31]_i_2_n_4 ),
        .Q(\alu0/div/rem [31]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[3] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[3]_i_1_n_4 ),
        .Q(\alu0/div/rem [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[4] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_7 ),
        .Q(\alu0/div/rem [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[5] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_6 ),
        .Q(\alu0/div/rem [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[6] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_5 ),
        .Q(\alu0/div/rem [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[7] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[7]_i_1_n_4 ),
        .Q(\alu0/div/rem [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[8] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_7 ),
        .Q(\alu0/div/rem [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/div/rrem/rem_reg[9] 
       (.C(clk),
        .CE(\rem[31]_i_1_n_0 ),
        .D(\rem_reg[11]_i_1_n_6 ),
        .Q(\alu0/div/rem [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[0] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[0]),
        .Q(\alu0/mul/mul_a [0]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[10] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[10]),
        .Q(\alu0/mul/mul_a [10]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[11] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[11]),
        .Q(\alu0/mul/mul_a [11]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[12] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[12]),
        .Q(\alu0/mul/mul_a [12]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[13] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[13]),
        .Q(\alu0/mul/mul_a [13]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[14] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[14]),
        .Q(\alu0/mul/mul_a [14]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[15] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[15]),
        .Q(\alu0/mul/mul_a [15]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[16] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\mul_a[16]_i_1_n_0 ),
        .Q(\alu0/mul/mul_a [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[17] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [17]),
        .Q(\alu0/mul/mul_a [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[18] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [18]),
        .Q(\alu0/mul/mul_a [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[19] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [19]),
        .Q(\alu0/mul/mul_a [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[1] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[1]),
        .Q(\alu0/mul/mul_a [1]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[20] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [20]),
        .Q(\alu0/mul/mul_a [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[21] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [21]),
        .Q(\alu0/mul/mul_a [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[22] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [22]),
        .Q(\alu0/mul/mul_a [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[23] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [23]),
        .Q(\alu0/mul/mul_a [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[24] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [24]),
        .Q(\alu0/mul/mul_a [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[25] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [25]),
        .Q(\alu0/mul/mul_a [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[26] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [26]),
        .Q(\alu0/mul/mul_a [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[27] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [27]),
        .Q(\alu0/mul/mul_a [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[28] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [28]),
        .Q(\alu0/mul/mul_a [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[29] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [29]),
        .Q(\alu0/mul/mul_a [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[2] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[2]),
        .Q(\alu0/mul/mul_a [2]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[30] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\alu0/mul_a_i [30]),
        .Q(\alu0/mul/mul_a [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mul_a_reg[31] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\mul_a[31]_i_1__0_n_0 ),
        .Q(\alu0/mul/mul_a [31]),
        .R(\<const0> ));
  FDRE \alu0/mul/mul_a_reg[32] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\mul_a[32]_i_1__0_n_0 ),
        .Q(\alu0/mul/mul_a [32]),
        .R(\<const0> ));
  FDRE \alu0/mul/mul_a_reg[3] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[3]),
        .Q(\alu0/mul/mul_a [3]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[4] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[4]),
        .Q(\alu0/mul/mul_a [4]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[5] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[5]),
        .Q(\alu0/mul/mul_a [5]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[6] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[6]),
        .Q(\alu0/mul/mul_a [6]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[7] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[7]),
        .Q(\alu0/mul/mul_a [7]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[8] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[8]),
        .Q(\alu0/mul/mul_a [8]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_a_reg[9] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(a0bus_0[9]),
        .Q(\alu0/mul/mul_a [9]),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[0] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[0]),
        .Q(\alu0/mul/mul_b_reg_n_0_[0] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[10] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[10]),
        .Q(\alu0/mul/mul_b_reg_n_0_[10] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[11] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[11]),
        .Q(\alu0/mul/mul_b_reg_n_0_[11] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[12] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[12]),
        .Q(\alu0/mul/mul_b_reg_n_0_[12] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[13] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[13]),
        .Q(\alu0/mul/mul_b_reg_n_0_[13] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[14] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[14]),
        .Q(\alu0/mul/mul_b_reg_n_0_[14] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[15] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[15]),
        .Q(\alu0/mul/mul_b_reg_n_0_[15] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[16] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[16]),
        .Q(\alu0/mul/mul_b_reg_n_0_[16] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[17] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[17]),
        .Q(\alu0/mul/mul_b_reg_n_0_[17] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[18] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[18]),
        .Q(\alu0/mul/mul_b_reg_n_0_[18] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[19] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[19]),
        .Q(\alu0/mul/mul_b_reg_n_0_[19] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[1] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[1]),
        .Q(\alu0/mul/mul_b_reg_n_0_[1] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[20] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[20]),
        .Q(\alu0/mul/mul_b_reg_n_0_[20] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[21] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[21]),
        .Q(\alu0/mul/mul_b_reg_n_0_[21] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[22] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[22]),
        .Q(\alu0/mul/mul_b_reg_n_0_[22] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[23] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[23]),
        .Q(\alu0/mul/mul_b_reg_n_0_[23] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[24] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[24]),
        .Q(\alu0/mul/mul_b_reg_n_0_[24] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[25] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[25]),
        .Q(\alu0/mul/mul_b_reg_n_0_[25] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[26] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[26]),
        .Q(\alu0/mul/mul_b_reg_n_0_[26] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[27] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[27]),
        .Q(\alu0/mul/mul_b_reg_n_0_[27] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[28] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[28]),
        .Q(\alu0/mul/mul_b_reg_n_0_[28] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[29] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[29]),
        .Q(\alu0/mul/mul_b_reg_n_0_[29] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[2] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[2]),
        .Q(\alu0/mul/mul_b_reg_n_0_[2] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[30] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[30]),
        .Q(\alu0/mul/mul_b_reg_n_0_[30] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[31] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\mul_b[31]_i_1_n_0 ),
        .Q(\alu0/mul/mul_b_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE \alu0/mul/mul_b_reg[32] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(\mul_b[32]_i_1_n_0 ),
        .Q(\alu0/mul/mul_b_reg_n_0_[32] ),
        .R(\<const0> ));
  FDRE \alu0/mul/mul_b_reg[3] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[3]),
        .Q(\alu0/mul/mul_b_reg_n_0_[3] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[4] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[4]),
        .Q(\alu0/mul/mul_b_reg_n_0_[4] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[5] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[5]),
        .Q(\alu0/mul/mul_b_reg_n_0_[5] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[6] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[6]),
        .Q(\alu0/mul/mul_b_reg_n_0_[6] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[7] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[7]),
        .Q(\alu0/mul/mul_b_reg_n_0_[7] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[8] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[8]),
        .Q(\alu0/mul/mul_b_reg_n_0_[8] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_b_reg[9] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(b0bus_0[9]),
        .Q(\alu0/mul/mul_b_reg_n_0_[9] ),
        .R(\mul_a[15]_i_1_n_0 ));
  FDRE \alu0/mul/mul_rslt_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu0/mul/mul_rslt0 ),
        .Q(\alu0/mul/mul_rslt ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu0/mul/mulh_reg[0] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[16]),
        .Q(\alu0/mul/mulh [0]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[10] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[26]),
        .Q(\alu0/mul/mulh [10]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[11] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[27]),
        .Q(\alu0/mul/mulh [11]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[12] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[28]),
        .Q(\alu0/mul/mulh [12]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[13] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[29]),
        .Q(\alu0/mul/mulh [13]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[14] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[30]),
        .Q(\alu0/mul/mulh [14]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[15] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[31]),
        .Q(\alu0/mul/mulh [15]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[1] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[17]),
        .Q(\alu0/mul/mulh [1]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[2] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[18]),
        .Q(\alu0/mul/mulh [2]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[3] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[19]),
        .Q(\alu0/mul/mulh [3]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[4] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[20]),
        .Q(\alu0/mul/mulh [4]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[5] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[21]),
        .Q(\alu0/mul/mulh [5]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[6] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[22]),
        .Q(\alu0/mul/mulh [6]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[7] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[23]),
        .Q(\alu0/mul/mulh [7]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[8] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[24]),
        .Q(\alu0/mul/mulh [8]),
        .R(\mulh[15]_i_1_n_0 ));
  FDRE \alu0/mul/mulh_reg[9] 
       (.C(clk),
        .CE(\alu0/mul/mul_b ),
        .D(niss_dsp_c0[25]),
        .Q(\alu0/mul/mulh [9]),
        .R(\mulh[15]_i_1_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry 
       (.CI(\<const0> ),
        .CO({\alu1/div/dadd/add_out0_carry_n_0 ,\alu1/div/dadd/add_out0_carry_n_1 ,\alu1/div/dadd/add_out0_carry_n_2 ,\alu1/div/dadd/add_out0_carry_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry_i_1__0_n_0,add_out0_carry_i_2__0_n_0,add_out0_carry_i_3__0_n_0,add_out0_carry_i_4__0_n_0}),
        .O(\alu1/div/add_out [3:0]),
        .S({add_out0_carry_i_5__0_n_0,add_out0_carry_i_6__0_n_0,add_out0_carry_i_7__0_n_0,add_out0_carry_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry__0 
       (.CI(\alu1/div/dadd/add_out0_carry_n_0 ),
        .CO({\alu1/div/dadd/add_out0_carry__0_n_0 ,\alu1/div/dadd/add_out0_carry__0_n_1 ,\alu1/div/dadd/add_out0_carry__0_n_2 ,\alu1/div/dadd/add_out0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__0_i_1__0_n_0,add_out0_carry__0_i_2__0_n_0,add_out0_carry__0_i_3__0_n_0,add_out0_carry__0_i_4__0_n_0}),
        .O(\alu1/div/add_out [7:4]),
        .S({add_out0_carry__0_i_5__0_n_0,add_out0_carry__0_i_6__0_n_0,add_out0_carry__0_i_7__0_n_0,add_out0_carry__0_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry__1 
       (.CI(\alu1/div/dadd/add_out0_carry__0_n_0 ),
        .CO({\alu1/div/dadd/add_out0_carry__1_n_0 ,\alu1/div/dadd/add_out0_carry__1_n_1 ,\alu1/div/dadd/add_out0_carry__1_n_2 ,\alu1/div/dadd/add_out0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__1_i_1__0_n_0,add_out0_carry__1_i_2__0_n_0,add_out0_carry__1_i_3__0_n_0,add_out0_carry__1_i_4__0_n_0}),
        .O(\alu1/div/add_out [11:8]),
        .S({add_out0_carry__1_i_5__0_n_0,add_out0_carry__1_i_6__0_n_0,add_out0_carry__1_i_7__0_n_0,add_out0_carry__1_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry__2 
       (.CI(\alu1/div/dadd/add_out0_carry__1_n_0 ),
        .CO({\alu1/div/dadd/add_out0_carry__2_n_0 ,\alu1/div/dadd/add_out0_carry__2_n_1 ,\alu1/div/dadd/add_out0_carry__2_n_2 ,\alu1/div/dadd/add_out0_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__2_i_1__0_n_0,add_out0_carry__2_i_2__0_n_0,add_out0_carry__2_i_3__0_n_0,add_out0_carry__2_i_4__0_n_0}),
        .O(\alu1/div/add_out [15:12]),
        .S({add_out0_carry__2_i_5__0_n_0,add_out0_carry__2_i_6__0_n_0,add_out0_carry__2_i_7__0_n_0,add_out0_carry__2_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry__3 
       (.CI(\alu1/div/dadd/add_out0_carry__2_n_0 ),
        .CO({\alu1/div/dadd/add_out0_carry__3_n_0 ,\alu1/div/dadd/add_out0_carry__3_n_1 ,\alu1/div/dadd/add_out0_carry__3_n_2 ,\alu1/div/dadd/add_out0_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__3_i_1__0_n_0,add_out0_carry__3_i_2__0_n_0,add_out0_carry__3_i_3__0_n_0,add_out0_carry__3_i_4__0_n_0}),
        .O(\alu1/div/add_out [19:16]),
        .S({add_out0_carry__3_i_5__0_n_0,add_out0_carry__3_i_6__0_n_0,add_out0_carry__3_i_7__0_n_0,add_out0_carry__3_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry__4 
       (.CI(\alu1/div/dadd/add_out0_carry__3_n_0 ),
        .CO({\alu1/div/dadd/add_out0_carry__4_n_0 ,\alu1/div/dadd/add_out0_carry__4_n_1 ,\alu1/div/dadd/add_out0_carry__4_n_2 ,\alu1/div/dadd/add_out0_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__4_i_1__0_n_0,add_out0_carry__4_i_2__0_n_0,add_out0_carry__4_i_3__0_n_0,add_out0_carry__4_i_4__0_n_0}),
        .O(\alu1/div/add_out [23:20]),
        .S({add_out0_carry__4_i_5__0_n_0,add_out0_carry__4_i_6__0_n_0,add_out0_carry__4_i_7__0_n_0,add_out0_carry__4_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry__5 
       (.CI(\alu1/div/dadd/add_out0_carry__4_n_0 ),
        .CO({\alu1/div/dadd/add_out0_carry__5_n_0 ,\alu1/div/dadd/add_out0_carry__5_n_1 ,\alu1/div/dadd/add_out0_carry__5_n_2 ,\alu1/div/dadd/add_out0_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({add_out0_carry__5_i_1__0_n_0,add_out0_carry__5_i_2__0_n_0,add_out0_carry__5_i_3__0_n_0,add_out0_carry__5_i_4__0_n_0}),
        .O(\alu1/div/add_out [27:24]),
        .S({add_out0_carry__5_i_5__0_n_0,add_out0_carry__5_i_6__0_n_0,add_out0_carry__5_i_7__0_n_0,add_out0_carry__5_i_8__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/dadd/add_out0_carry__6 
       (.CI(\alu1/div/dadd/add_out0_carry__5_n_0 ),
        .CO({\alu1/div/dadd/add_out0_carry__6_n_1 ,\alu1/div/dadd/add_out0_carry__6_n_2 ,\alu1/div/dadd/add_out0_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,add_out0_carry__6_i_1__0_n_0,add_out0_carry__6_i_2__0_n_0,add_out0_carry__6_i_3__0_n_0}),
        .O(\alu1/div/add_out [31:28]),
        .S({add_out0_carry__6_i_4__0_n_0,add_out0_carry__6_i_5__0_n_0,add_out0_carry__6_i_6__0_n_0,add_out0_carry__6_i_7__0_n_0}));
  FDRE \alu1/div/dctl/dctl_long_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/div/dctl_long ),
        .Q(\alu1/div/dctl/dctl_long_f ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/dctl_sign_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/div/dctl/dctl_sign ),
        .Q(\alu1/div/dctl/dctl_sign_f ),
        .R(\alu1/div/p_0_in__0 ));
  FDSE \alu1/div/dctl/div_crdy_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(div_crdy_i_1__0_n_0),
        .Q(div_crdy1),
        .S(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/fsm/chg_quo_sgn_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_quo_sgn_i_1__0_n_0),
        .Q(\alu1/div/chg_quo_sgn ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/fsm/chg_rem_sgn_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_rem_sgn_i_1__0_n_0),
        .Q(\alu1/div/chg_rem_sgn ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/fsm/dctl_stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/div/dctl/fsm/dctl_next [0]),
        .Q(\alu1/div/dctl_stat [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/fsm/dctl_stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/div/dctl/fsm/dctl_next [1]),
        .Q(\alu1/div/dctl_stat [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/fsm/dctl_stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/div/dctl/fsm/dctl_next [2]),
        .Q(\alu1/div/dctl_stat [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/fsm/dctl_stat_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/div/dctl/fsm/dctl_next [3]),
        .Q(\alu1/div/dctl_stat [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/dctl/fsm/fdiv_rem_msb_f_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/div/p_0_in0 ),
        .Q(\alu1/div/fdiv_rem_msb_f ),
        .R(\alu1/div/p_0_in__0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry 
       (.CI(\<const0> ),
        .CO({\alu1/div/fdiv/rem0_carry_n_0 ,\alu1/div/fdiv/rem0_carry_n_1 ,\alu1/div/fdiv/rem0_carry_n_2 ,\alu1/div/fdiv/rem0_carry_n_3 }),
        .CYINIT(rem0_carry_i_1__0_n_0),
        .DI({\alu1/div/rem1__0 [3:1],\alu1/div/den [28]}),
        .O(\alu1/div/fdiv_rem [3:0]),
        .S({rem0_carry_i_2__0_n_0,rem0_carry_i_3__0_n_0,rem0_carry_i_4__0_n_0,rem0_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__0 
       (.CI(\alu1/div/fdiv/rem0_carry_n_0 ),
        .CO({\alu1/div/fdiv/rem0_carry__0_n_0 ,\alu1/div/fdiv/rem0_carry__0_n_1 ,\alu1/div/fdiv/rem0_carry__0_n_2 ,\alu1/div/fdiv/rem0_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem1__0 [7:4]),
        .O(\alu1/div/fdiv_rem [7:4]),
        .S({rem0_carry__0_i_1__0_n_0,rem0_carry__0_i_2__0_n_0,rem0_carry__0_i_3__0_n_0,rem0_carry__0_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__1 
       (.CI(\alu1/div/fdiv/rem0_carry__0_n_0 ),
        .CO({\alu1/div/fdiv/rem0_carry__1_n_0 ,\alu1/div/fdiv/rem0_carry__1_n_1 ,\alu1/div/fdiv/rem0_carry__1_n_2 ,\alu1/div/fdiv/rem0_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem1__0 [11:8]),
        .O(\alu1/div/fdiv_rem [11:8]),
        .S({rem0_carry__1_i_1__0_n_0,rem0_carry__1_i_2__0_n_0,rem0_carry__1_i_3__0_n_0,rem0_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__2 
       (.CI(\alu1/div/fdiv/rem0_carry__1_n_0 ),
        .CO({\alu1/div/fdiv/rem0_carry__2_n_0 ,\alu1/div/fdiv/rem0_carry__2_n_1 ,\alu1/div/fdiv/rem0_carry__2_n_2 ,\alu1/div/fdiv/rem0_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem1__0 [15:12]),
        .O(\alu1/div/fdiv_rem [15:12]),
        .S({rem0_carry__2_i_1__0_n_0,rem0_carry__2_i_2__0_n_0,rem0_carry__2_i_3__0_n_0,rem0_carry__2_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__3 
       (.CI(\alu1/div/fdiv/rem0_carry__2_n_0 ),
        .CO({\alu1/div/fdiv/rem0_carry__3_n_0 ,\alu1/div/fdiv/rem0_carry__3_n_1 ,\alu1/div/fdiv/rem0_carry__3_n_2 ,\alu1/div/fdiv/rem0_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem1__0 [19:16]),
        .O(\alu1/div/fdiv_rem [19:16]),
        .S({rem0_carry__3_i_1__0_n_0,rem0_carry__3_i_2__0_n_0,rem0_carry__3_i_3__0_n_0,rem0_carry__3_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__4 
       (.CI(\alu1/div/fdiv/rem0_carry__3_n_0 ),
        .CO({\alu1/div/fdiv/rem0_carry__4_n_0 ,\alu1/div/fdiv/rem0_carry__4_n_1 ,\alu1/div/fdiv/rem0_carry__4_n_2 ,\alu1/div/fdiv/rem0_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem1__0 [23:20]),
        .O(\alu1/div/fdiv_rem [23:20]),
        .S({rem0_carry__4_i_1__0_n_0,rem0_carry__4_i_2__0_n_0,rem0_carry__4_i_3__0_n_0,rem0_carry__4_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__5 
       (.CI(\alu1/div/fdiv/rem0_carry__4_n_0 ),
        .CO({\alu1/div/fdiv/rem0_carry__5_n_0 ,\alu1/div/fdiv/rem0_carry__5_n_1 ,\alu1/div/fdiv/rem0_carry__5_n_2 ,\alu1/div/fdiv/rem0_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem1__0 [27:24]),
        .O(\alu1/div/fdiv_rem [27:24]),
        .S({rem0_carry__5_i_1__0_n_0,rem0_carry__5_i_2__0_n_0,rem0_carry__5_i_3__0_n_0,rem0_carry__5_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__6 
       (.CI(\alu1/div/fdiv/rem0_carry__5_n_0 ),
        .CO({\alu1/div/fdiv/rem0_carry__6_n_0 ,\alu1/div/fdiv/rem0_carry__6_n_1 ,\alu1/div/fdiv/rem0_carry__6_n_2 ,\alu1/div/fdiv/rem0_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem1__0 [31:28]),
        .O(\alu1/div/fdiv_rem [31:28]),
        .S({rem0_carry__6_i_1__0_n_0,rem0_carry__6_i_2__0_n_0,rem0_carry__6_i_3__0_n_0,rem0_carry__6_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem0_carry__7 
       (.CI(\alu1/div/fdiv/rem0_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu1/div/p_0_in0 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem0_carry__7_i_1__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry 
       (.CI(\<const0> ),
        .CO({\alu1/div/fdiv/rem1_carry_n_0 ,\alu1/div/fdiv/rem1_carry_n_1 ,\alu1/div/fdiv/rem1_carry_n_2 ,\alu1/div/fdiv/rem1_carry_n_3 }),
        .CYINIT(rem1_carry_i_1__0_n_0),
        .DI({\alu1/div/rem2__0 [3:1],\alu1/div/den [29]}),
        .O(\alu1/div/rem1__0 [4:1]),
        .S({rem1_carry_i_2__0_n_0,rem1_carry_i_3__0_n_0,rem1_carry_i_4__0_n_0,rem1_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__0 
       (.CI(\alu1/div/fdiv/rem1_carry_n_0 ),
        .CO({\alu1/div/fdiv/rem1_carry__0_n_0 ,\alu1/div/fdiv/rem1_carry__0_n_1 ,\alu1/div/fdiv/rem1_carry__0_n_2 ,\alu1/div/fdiv/rem1_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem2__0 [7:4]),
        .O(\alu1/div/rem1__0 [8:5]),
        .S({rem1_carry__0_i_1__0_n_0,rem1_carry__0_i_2__0_n_0,rem1_carry__0_i_3__0_n_0,rem1_carry__0_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__1 
       (.CI(\alu1/div/fdiv/rem1_carry__0_n_0 ),
        .CO({\alu1/div/fdiv/rem1_carry__1_n_0 ,\alu1/div/fdiv/rem1_carry__1_n_1 ,\alu1/div/fdiv/rem1_carry__1_n_2 ,\alu1/div/fdiv/rem1_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem2__0 [11:8]),
        .O(\alu1/div/rem1__0 [12:9]),
        .S({rem1_carry__1_i_1__0_n_0,rem1_carry__1_i_2__0_n_0,rem1_carry__1_i_3__0_n_0,rem1_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__2 
       (.CI(\alu1/div/fdiv/rem1_carry__1_n_0 ),
        .CO({\alu1/div/fdiv/rem1_carry__2_n_0 ,\alu1/div/fdiv/rem1_carry__2_n_1 ,\alu1/div/fdiv/rem1_carry__2_n_2 ,\alu1/div/fdiv/rem1_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem2__0 [15:12]),
        .O(\alu1/div/rem1__0 [16:13]),
        .S({rem1_carry__2_i_1__0_n_0,rem1_carry__2_i_2__0_n_0,rem1_carry__2_i_3__0_n_0,rem1_carry__2_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__3 
       (.CI(\alu1/div/fdiv/rem1_carry__2_n_0 ),
        .CO({\alu1/div/fdiv/rem1_carry__3_n_0 ,\alu1/div/fdiv/rem1_carry__3_n_1 ,\alu1/div/fdiv/rem1_carry__3_n_2 ,\alu1/div/fdiv/rem1_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem2__0 [19:16]),
        .O(\alu1/div/rem1__0 [20:17]),
        .S({rem1_carry__3_i_1__0_n_0,rem1_carry__3_i_2__0_n_0,rem1_carry__3_i_3__0_n_0,rem1_carry__3_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__4 
       (.CI(\alu1/div/fdiv/rem1_carry__3_n_0 ),
        .CO({\alu1/div/fdiv/rem1_carry__4_n_0 ,\alu1/div/fdiv/rem1_carry__4_n_1 ,\alu1/div/fdiv/rem1_carry__4_n_2 ,\alu1/div/fdiv/rem1_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem2__0 [23:20]),
        .O(\alu1/div/rem1__0 [24:21]),
        .S({rem1_carry__4_i_1__0_n_0,rem1_carry__4_i_2__0_n_0,rem1_carry__4_i_3__0_n_0,rem1_carry__4_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__5 
       (.CI(\alu1/div/fdiv/rem1_carry__4_n_0 ),
        .CO({\alu1/div/fdiv/rem1_carry__5_n_0 ,\alu1/div/fdiv/rem1_carry__5_n_1 ,\alu1/div/fdiv/rem1_carry__5_n_2 ,\alu1/div/fdiv/rem1_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem2__0 [27:24]),
        .O(\alu1/div/rem1__0 [28:25]),
        .S({rem1_carry__5_i_1__0_n_0,rem1_carry__5_i_2__0_n_0,rem1_carry__5_i_3__0_n_0,rem1_carry__5_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__6 
       (.CI(\alu1/div/fdiv/rem1_carry__5_n_0 ),
        .CO({\alu1/div/fdiv/rem1_carry__6_n_0 ,\alu1/div/fdiv/rem1_carry__6_n_1 ,\alu1/div/fdiv/rem1_carry__6_n_2 ,\alu1/div/fdiv/rem1_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem2__0 [31:28]),
        .O(\alu1/div/rem1__0 [32:29]),
        .S({rem1_carry__6_i_1__0_n_0,rem1_carry__6_i_2__0_n_0,rem1_carry__6_i_3__0_n_0,rem1_carry__6_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem1_carry__7 
       (.CI(\alu1/div/fdiv/rem1_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu1/div/rem1 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem1_carry__7_i_1__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry 
       (.CI(\<const0> ),
        .CO({\alu1/div/fdiv/rem2_carry_n_0 ,\alu1/div/fdiv/rem2_carry_n_1 ,\alu1/div/fdiv/rem2_carry_n_2 ,\alu1/div/fdiv/rem2_carry_n_3 }),
        .CYINIT(\alu1/div/fdiv/p_1_in3_in ),
        .DI({\alu1/div/rem3__0 [3:1],\alu1/div/den [30]}),
        .O(\alu1/div/rem2__0 [4:1]),
        .S({rem2_carry_i_2__0_n_0,rem2_carry_i_3__0_n_0,rem2_carry_i_4__0_n_0,rem2_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__0 
       (.CI(\alu1/div/fdiv/rem2_carry_n_0 ),
        .CO({\alu1/div/fdiv/rem2_carry__0_n_0 ,\alu1/div/fdiv/rem2_carry__0_n_1 ,\alu1/div/fdiv/rem2_carry__0_n_2 ,\alu1/div/fdiv/rem2_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem3__0 [7:4]),
        .O(\alu1/div/rem2__0 [8:5]),
        .S({rem2_carry__0_i_1__0_n_0,rem2_carry__0_i_2__0_n_0,rem2_carry__0_i_3__0_n_0,rem2_carry__0_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__1 
       (.CI(\alu1/div/fdiv/rem2_carry__0_n_0 ),
        .CO({\alu1/div/fdiv/rem2_carry__1_n_0 ,\alu1/div/fdiv/rem2_carry__1_n_1 ,\alu1/div/fdiv/rem2_carry__1_n_2 ,\alu1/div/fdiv/rem2_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem3__0 [11:8]),
        .O(\alu1/div/rem2__0 [12:9]),
        .S({rem2_carry__1_i_1__0_n_0,rem2_carry__1_i_2__0_n_0,rem2_carry__1_i_3__0_n_0,rem2_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__2 
       (.CI(\alu1/div/fdiv/rem2_carry__1_n_0 ),
        .CO({\alu1/div/fdiv/rem2_carry__2_n_0 ,\alu1/div/fdiv/rem2_carry__2_n_1 ,\alu1/div/fdiv/rem2_carry__2_n_2 ,\alu1/div/fdiv/rem2_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem3__0 [15:12]),
        .O(\alu1/div/rem2__0 [16:13]),
        .S({rem2_carry__2_i_1__0_n_0,rem2_carry__2_i_2__0_n_0,rem2_carry__2_i_3__0_n_0,rem2_carry__2_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__3 
       (.CI(\alu1/div/fdiv/rem2_carry__2_n_0 ),
        .CO({\alu1/div/fdiv/rem2_carry__3_n_0 ,\alu1/div/fdiv/rem2_carry__3_n_1 ,\alu1/div/fdiv/rem2_carry__3_n_2 ,\alu1/div/fdiv/rem2_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem3__0 [19:16]),
        .O(\alu1/div/rem2__0 [20:17]),
        .S({rem2_carry__3_i_1__0_n_0,rem2_carry__3_i_2__0_n_0,rem2_carry__3_i_3__0_n_0,rem2_carry__3_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__4 
       (.CI(\alu1/div/fdiv/rem2_carry__3_n_0 ),
        .CO({\alu1/div/fdiv/rem2_carry__4_n_0 ,\alu1/div/fdiv/rem2_carry__4_n_1 ,\alu1/div/fdiv/rem2_carry__4_n_2 ,\alu1/div/fdiv/rem2_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem3__0 [23:20]),
        .O(\alu1/div/rem2__0 [24:21]),
        .S({rem2_carry__4_i_1__0_n_0,rem2_carry__4_i_2__0_n_0,rem2_carry__4_i_3__0_n_0,rem2_carry__4_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__5 
       (.CI(\alu1/div/fdiv/rem2_carry__4_n_0 ),
        .CO({\alu1/div/fdiv/rem2_carry__5_n_0 ,\alu1/div/fdiv/rem2_carry__5_n_1 ,\alu1/div/fdiv/rem2_carry__5_n_2 ,\alu1/div/fdiv/rem2_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem3__0 [27:24]),
        .O(\alu1/div/rem2__0 [28:25]),
        .S({rem2_carry__5_i_1__0_n_0,rem2_carry__5_i_2__0_n_0,rem2_carry__5_i_3__0_n_0,rem2_carry__5_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__6 
       (.CI(\alu1/div/fdiv/rem2_carry__5_n_0 ),
        .CO({\alu1/div/fdiv/rem2_carry__6_n_0 ,\alu1/div/fdiv/rem2_carry__6_n_1 ,\alu1/div/fdiv/rem2_carry__6_n_2 ,\alu1/div/fdiv/rem2_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/rem3__0 [31:28]),
        .O(\alu1/div/rem2__0 [32:29]),
        .S({rem2_carry__6_i_1__0_n_0,rem2_carry__6_i_2__0_n_0,rem2_carry__6_i_3__0_n_0,rem2_carry__6_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem2_carry__7 
       (.CI(\alu1/div/fdiv/rem2_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu1/div/rem2 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem2_carry__7_i_1__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry 
       (.CI(\<const0> ),
        .CO({\alu1/div/fdiv/rem3_carry_n_0 ,\alu1/div/fdiv/rem3_carry_n_1 ,\alu1/div/fdiv/rem3_carry_n_2 ,\alu1/div/fdiv/rem3_carry_n_3 }),
        .CYINIT(\alu1/div/fdiv/p_1_in5_in ),
        .DI({\alu1/div/den [34:32],\alu1/div/den2 }),
        .O(\alu1/div/rem3__0 [4:1]),
        .S({rem3_carry_i_2__0_n_0,rem3_carry_i_3__0_n_0,rem3_carry_i_4__0_n_0,rem3_carry_i_5__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__0 
       (.CI(\alu1/div/fdiv/rem3_carry_n_0 ),
        .CO({\alu1/div/fdiv/rem3_carry__0_n_0 ,\alu1/div/fdiv/rem3_carry__0_n_1 ,\alu1/div/fdiv/rem3_carry__0_n_2 ,\alu1/div/fdiv/rem3_carry__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/den [38:35]),
        .O(\alu1/div/rem3__0 [8:5]),
        .S({rem3_carry__0_i_1__0_n_0,rem3_carry__0_i_2__0_n_0,rem3_carry__0_i_3__0_n_0,rem3_carry__0_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__1 
       (.CI(\alu1/div/fdiv/rem3_carry__0_n_0 ),
        .CO({\alu1/div/fdiv/rem3_carry__1_n_0 ,\alu1/div/fdiv/rem3_carry__1_n_1 ,\alu1/div/fdiv/rem3_carry__1_n_2 ,\alu1/div/fdiv/rem3_carry__1_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/den [42:39]),
        .O(\alu1/div/rem3__0 [12:9]),
        .S({rem3_carry__1_i_1__0_n_0,rem3_carry__1_i_2__0_n_0,rem3_carry__1_i_3__0_n_0,rem3_carry__1_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__2 
       (.CI(\alu1/div/fdiv/rem3_carry__1_n_0 ),
        .CO({\alu1/div/fdiv/rem3_carry__2_n_0 ,\alu1/div/fdiv/rem3_carry__2_n_1 ,\alu1/div/fdiv/rem3_carry__2_n_2 ,\alu1/div/fdiv/rem3_carry__2_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/den [46:43]),
        .O(\alu1/div/rem3__0 [16:13]),
        .S({rem3_carry__2_i_1__0_n_0,rem3_carry__2_i_2__0_n_0,rem3_carry__2_i_3__0_n_0,rem3_carry__2_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__3 
       (.CI(\alu1/div/fdiv/rem3_carry__2_n_0 ),
        .CO({\alu1/div/fdiv/rem3_carry__3_n_0 ,\alu1/div/fdiv/rem3_carry__3_n_1 ,\alu1/div/fdiv/rem3_carry__3_n_2 ,\alu1/div/fdiv/rem3_carry__3_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/den [50:47]),
        .O(\alu1/div/rem3__0 [20:17]),
        .S({rem3_carry__3_i_1__0_n_0,rem3_carry__3_i_2__0_n_0,rem3_carry__3_i_3__0_n_0,rem3_carry__3_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__4 
       (.CI(\alu1/div/fdiv/rem3_carry__3_n_0 ),
        .CO({\alu1/div/fdiv/rem3_carry__4_n_0 ,\alu1/div/fdiv/rem3_carry__4_n_1 ,\alu1/div/fdiv/rem3_carry__4_n_2 ,\alu1/div/fdiv/rem3_carry__4_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/den [54:51]),
        .O(\alu1/div/rem3__0 [24:21]),
        .S({rem3_carry__4_i_1__0_n_0,rem3_carry__4_i_2__0_n_0,rem3_carry__4_i_3__0_n_0,rem3_carry__4_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__5 
       (.CI(\alu1/div/fdiv/rem3_carry__4_n_0 ),
        .CO({\alu1/div/fdiv/rem3_carry__5_n_0 ,\alu1/div/fdiv/rem3_carry__5_n_1 ,\alu1/div/fdiv/rem3_carry__5_n_2 ,\alu1/div/fdiv/rem3_carry__5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/den [58:55]),
        .O(\alu1/div/rem3__0 [28:25]),
        .S({rem3_carry__5_i_1__0_n_0,rem3_carry__5_i_2__0_n_0,rem3_carry__5_i_3__0_n_0,rem3_carry__5_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__6 
       (.CI(\alu1/div/fdiv/rem3_carry__5_n_0 ),
        .CO({\alu1/div/fdiv/rem3_carry__6_n_0 ,\alu1/div/fdiv/rem3_carry__6_n_1 ,\alu1/div/fdiv/rem3_carry__6_n_2 ,\alu1/div/fdiv/rem3_carry__6_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\alu1/div/den [62:59]),
        .O(\alu1/div/rem3__0 [32:29]),
        .S({rem3_carry__6_i_1__0_n_0,rem3_carry__6_i_2__0_n_0,rem3_carry__6_i_3__0_n_0,rem3_carry__6_i_4__0_n_0}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \alu1/div/fdiv/rem3_carry__7 
       (.CI(\alu1/div/fdiv/rem3_carry__6_n_0 ),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\alu1/div/rem3 ),
        .S({\<const0> ,\<const0> ,\<const0> ,rem3_carry__7_i_1__0_n_0}));
  FDRE \alu1/div/rden/remden_reg[0] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[0]_i_1__0_n_0 ),
        .Q(\alu1/div/den [0]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[10] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[10]_i_1__0_n_0 ),
        .Q(\alu1/div/den [10]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[11] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[11]_i_1__0_n_0 ),
        .Q(\alu1/div/den [11]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[12] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[12]_i_1__0_n_0 ),
        .Q(\alu1/div/den [12]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[13] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[13]_i_1__0_n_0 ),
        .Q(\alu1/div/den [13]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[14] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[14]_i_1__0_n_0 ),
        .Q(\alu1/div/den [14]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[15] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[15]_i_1__0_n_0 ),
        .Q(\alu1/div/den [15]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[16] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[16]_i_1__0_n_0 ),
        .Q(\alu1/div/den [16]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[17] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[17]_i_1__0_n_0 ),
        .Q(\alu1/div/den [17]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[18] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[18]_i_1__0_n_0 ),
        .Q(\alu1/div/den [18]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[19] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[19]_i_1__0_n_0 ),
        .Q(\alu1/div/den [19]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[1] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[1]_i_1__0_n_0 ),
        .Q(\alu1/div/den [1]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[20] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[20]_i_1__0_n_0 ),
        .Q(\alu1/div/den [20]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[21] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[21]_i_1__0_n_0 ),
        .Q(\alu1/div/den [21]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[22] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[22]_i_1__0_n_0 ),
        .Q(\alu1/div/den [22]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[23] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[23]_i_1__0_n_0 ),
        .Q(\alu1/div/den [23]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[24] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[24]_i_1__0_n_0 ),
        .Q(\alu1/div/den [24]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[25] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[25]_i_1__0_n_0 ),
        .Q(\alu1/div/den [25]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[26] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[26]_i_1__0_n_0 ),
        .Q(\alu1/div/den [26]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[27] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[27]_i_1__0_n_0 ),
        .Q(\alu1/div/den [27]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[28] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[28]_i_1__0_n_0 ),
        .Q(\alu1/div/den [28]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[29] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[29]_i_1__0_n_0 ),
        .Q(\alu1/div/den [29]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[2] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[2]_i_1__0_n_0 ),
        .Q(\alu1/div/den [2]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[30] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[30]_i_1__0_n_0 ),
        .Q(\alu1/div/den [30]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[31] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[31]_i_2__0_n_0 ),
        .Q(\alu1/div/den2 ),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[32] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[32]_i_1__0_n_0 ),
        .Q(\alu1/div/den [32]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[33] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[33]_i_1__0_n_0 ),
        .Q(\alu1/div/den [33]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[34] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[34]_i_1__0_n_0 ),
        .Q(\alu1/div/den [34]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[35] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[35]_i_1__0_n_0 ),
        .Q(\alu1/div/den [35]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[36] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[36]_i_1__0_n_0 ),
        .Q(\alu1/div/den [36]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[37] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[37]_i_1__0_n_0 ),
        .Q(\alu1/div/den [37]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[38] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[38]_i_1__0_n_0 ),
        .Q(\alu1/div/den [38]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[39] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[39]_i_1__0_n_0 ),
        .Q(\alu1/div/den [39]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[3] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[3]_i_1__0_n_0 ),
        .Q(\alu1/div/den [3]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[40] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[40]_i_1__0_n_0 ),
        .Q(\alu1/div/den [40]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[41] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[41]_i_1__0_n_0 ),
        .Q(\alu1/div/den [41]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[42] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[42]_i_1__0_n_0 ),
        .Q(\alu1/div/den [42]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[43] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[43]_i_1__0_n_0 ),
        .Q(\alu1/div/den [43]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[44] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[44]_i_1__0_n_0 ),
        .Q(\alu1/div/den [44]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[45] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[45]_i_1__0_n_0 ),
        .Q(\alu1/div/den [45]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[46] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[46]_i_1__0_n_0 ),
        .Q(\alu1/div/den [46]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[47] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[47]_i_1__0_n_0 ),
        .Q(\alu1/div/den [47]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[48] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[48]_i_1__0_n_0 ),
        .Q(\alu1/div/den [48]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[49] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[49]_i_1__0_n_0 ),
        .Q(\alu1/div/den [49]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[4] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[4]_i_1__0_n_0 ),
        .Q(\alu1/div/den [4]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[50] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[50]_i_1__0_n_0 ),
        .Q(\alu1/div/den [50]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[51] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[51]_i_1__0_n_0 ),
        .Q(\alu1/div/den [51]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[52] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[52]_i_1__0_n_0 ),
        .Q(\alu1/div/den [52]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[53] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[53]_i_1__0_n_0 ),
        .Q(\alu1/div/den [53]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[54] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[54]_i_1__0_n_0 ),
        .Q(\alu1/div/den [54]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[55] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[55]_i_1__0_n_0 ),
        .Q(\alu1/div/den [55]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[56] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[56]_i_1__0_n_0 ),
        .Q(\alu1/div/den [56]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[57] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[57]_i_1__0_n_0 ),
        .Q(\alu1/div/den [57]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[58] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[58]_i_1__0_n_0 ),
        .Q(\alu1/div/den [58]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[59] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[59]_i_1__0_n_0 ),
        .Q(\alu1/div/den [59]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[5] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[5]_i_1__0_n_0 ),
        .Q(\alu1/div/den [5]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[60] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[60]_i_1__0_n_0 ),
        .Q(\alu1/div/den [60]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[61] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[61]_i_1__0_n_0 ),
        .Q(\alu1/div/den [61]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[62] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[62]_i_1__0_n_0 ),
        .Q(\alu1/div/den [62]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[63] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[63]_i_1__0_n_0 ),
        .Q(\alu1/div/den [63]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[64] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[64]_i_3__0_n_0 ),
        .Q(\alu1/div/den [64]),
        .R(\remden[64]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[6] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[6]_i_1__0_n_0 ),
        .Q(\alu1/div/den [6]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[7] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[7]_i_1__0_n_0 ),
        .Q(\alu1/div/den [7]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[8] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[8]_i_1__0_n_0 ),
        .Q(\alu1/div/den [8]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rden/remden_reg[9] 
       (.C(clk),
        .CE(\remden[64]_i_2__0_n_0 ),
        .D(\remden[9]_i_1__0_n_0 ),
        .Q(\alu1/div/den [9]),
        .R(\remden[31]_i_1__0_n_0 ));
  FDRE \alu1/div/rdso/dso_reg[0] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[3]_i_1__0_n_7 ),
        .Q(\alu1/div/dso_0 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[10] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[11]_i_1__0_n_5 ),
        .Q(\alu1/div/dso_0 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[11] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[11]_i_1__0_n_4 ),
        .Q(\alu1/div/dso_0 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[12] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[15]_i_1__0_n_7 ),
        .Q(\alu1/div/dso_0 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[13] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[15]_i_1__0_n_6 ),
        .Q(\alu1/div/dso_0 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[14] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[15]_i_1__0_n_5 ),
        .Q(\alu1/div/dso_0 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[15] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[15]_i_1__0_n_4 ),
        .Q(\alu1/div/dso_0 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[16] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[19]_i_1__0_n_7 ),
        .Q(\alu1/div/dso_0 [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[17] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[19]_i_1__0_n_6 ),
        .Q(\alu1/div/dso_0 [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[18] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[19]_i_1__0_n_5 ),
        .Q(\alu1/div/dso_0 [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[19] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[19]_i_1__0_n_4 ),
        .Q(\alu1/div/dso_0 [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[1] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[3]_i_1__0_n_6 ),
        .Q(\alu1/div/dso_0 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[20] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[23]_i_1__0_n_7 ),
        .Q(\alu1/div/dso_0 [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[21] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[23]_i_1__0_n_6 ),
        .Q(\alu1/div/dso_0 [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[22] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[23]_i_1__0_n_5 ),
        .Q(\alu1/div/dso_0 [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[23] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[23]_i_1__0_n_4 ),
        .Q(\alu1/div/dso_0 [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[24] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[27]_i_1__0_n_7 ),
        .Q(\alu1/div/dso_0 [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[25] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[27]_i_1__0_n_6 ),
        .Q(\alu1/div/dso_0 [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[26] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[27]_i_1__0_n_5 ),
        .Q(\alu1/div/dso_0 [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[27] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[27]_i_1__0_n_4 ),
        .Q(\alu1/div/dso_0 [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[28] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[31]_i_2__0_n_7 ),
        .Q(\alu1/div/dso_0 [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[29] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[31]_i_2__0_n_6 ),
        .Q(\alu1/div/dso_0 [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[2] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[3]_i_1__0_n_5 ),
        .Q(\alu1/div/dso_0 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[30] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[31]_i_2__0_n_5 ),
        .Q(\alu1/div/dso_0 [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[31] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[31]_i_2__0_n_4 ),
        .Q(\alu1/div/dso_0 [31]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[3] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[3]_i_1__0_n_4 ),
        .Q(\alu1/div/dso_0 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[4] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[7]_i_1__0_n_7 ),
        .Q(\alu1/div/dso_0 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[5] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[7]_i_1__0_n_6 ),
        .Q(\alu1/div/dso_0 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[6] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[7]_i_1__0_n_5 ),
        .Q(\alu1/div/dso_0 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[7] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[7]_i_1__0_n_4 ),
        .Q(\alu1/div/dso_0 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[8] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[11]_i_1__0_n_7 ),
        .Q(\alu1/div/dso_0 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rdso/dso_reg[9] 
       (.C(clk),
        .CE(\dso[31]_i_1__0_n_0 ),
        .D(\dso_reg[11]_i_1__0_n_6 ),
        .Q(\alu1/div/dso_0 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[0] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [0]),
        .Q(\alu1/div/quo [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[10] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [10]),
        .Q(\alu1/div/quo [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[11] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [11]),
        .Q(\alu1/div/quo [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[12] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [12]),
        .Q(\alu1/div/quo [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[13] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [13]),
        .Q(\alu1/div/quo [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[14] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [14]),
        .Q(\alu1/div/quo [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[15] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [15]),
        .Q(\alu1/div/quo [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[16] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [16]),
        .Q(\alu1/div/quo [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[17] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [17]),
        .Q(\alu1/div/quo [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[18] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [18]),
        .Q(\alu1/div/quo [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[19] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [19]),
        .Q(\alu1/div/quo [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[1] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [1]),
        .Q(\alu1/div/quo [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[20] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [20]),
        .Q(\alu1/div/quo [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[21] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [21]),
        .Q(\alu1/div/quo [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[22] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [22]),
        .Q(\alu1/div/quo [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[23] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [23]),
        .Q(\alu1/div/quo [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[24] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [24]),
        .Q(\alu1/div/quo [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[25] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [25]),
        .Q(\alu1/div/quo [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[26] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [26]),
        .Q(\alu1/div/quo [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[27] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [27]),
        .Q(\alu1/div/quo [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[28] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [28]),
        .Q(\alu1/div/quo__0 [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[29] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [29]),
        .Q(\alu1/div/quo__0 [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[2] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [2]),
        .Q(\alu1/div/quo [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[30] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [30]),
        .Q(\alu1/div/quo__0 [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[31] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [31]),
        .Q(\alu1/div/quo__0 [31]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[3] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [3]),
        .Q(\alu1/div/quo [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[4] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [4]),
        .Q(\alu1/div/quo [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[5] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [5]),
        .Q(\alu1/div/quo [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[6] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [6]),
        .Q(\alu1/div/quo [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[7] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [7]),
        .Q(\alu1/div/quo [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[8] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [8]),
        .Q(\alu1/div/quo [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rquo/quo_reg[9] 
       (.C(clk),
        .CE(\quo[31]_i_1__0_n_0 ),
        .D(\alu1/div/p_2_in [9]),
        .Q(\alu1/div/quo [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[0] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[3]_i_1__0_n_7 ),
        .Q(\alu1/div/rem [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[10] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[11]_i_1__0_n_5 ),
        .Q(\alu1/div/rem [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[11] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[11]_i_1__0_n_4 ),
        .Q(\alu1/div/rem [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[12] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[15]_i_1__0_n_7 ),
        .Q(\alu1/div/rem [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[13] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[15]_i_1__0_n_6 ),
        .Q(\alu1/div/rem [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[14] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[15]_i_1__0_n_5 ),
        .Q(\alu1/div/rem [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[15] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[15]_i_1__0_n_4 ),
        .Q(\alu1/div/rem [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[16] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[19]_i_1__0_n_7 ),
        .Q(\alu1/div/rem [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[17] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[19]_i_1__0_n_6 ),
        .Q(\alu1/div/rem [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[18] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[19]_i_1__0_n_5 ),
        .Q(\alu1/div/rem [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[19] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[19]_i_1__0_n_4 ),
        .Q(\alu1/div/rem [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[1] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[3]_i_1__0_n_6 ),
        .Q(\alu1/div/rem [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[20] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[23]_i_1__0_n_7 ),
        .Q(\alu1/div/rem [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[21] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[23]_i_1__0_n_6 ),
        .Q(\alu1/div/rem [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[22] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[23]_i_1__0_n_5 ),
        .Q(\alu1/div/rem [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[23] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[23]_i_1__0_n_4 ),
        .Q(\alu1/div/rem [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[24] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[27]_i_1__0_n_7 ),
        .Q(\alu1/div/rem [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[25] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[27]_i_1__0_n_6 ),
        .Q(\alu1/div/rem [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[26] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[27]_i_1__0_n_5 ),
        .Q(\alu1/div/rem [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[27] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[27]_i_1__0_n_4 ),
        .Q(\alu1/div/rem [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[28] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[31]_i_2__0_n_7 ),
        .Q(\alu1/div/rem [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[29] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[31]_i_2__0_n_6 ),
        .Q(\alu1/div/rem [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[2] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[3]_i_1__0_n_5 ),
        .Q(\alu1/div/rem [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[30] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[31]_i_2__0_n_5 ),
        .Q(\alu1/div/rem [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[31] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[31]_i_2__0_n_4 ),
        .Q(\alu1/div/rem [31]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[3] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[3]_i_1__0_n_4 ),
        .Q(\alu1/div/rem [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[4] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[7]_i_1__0_n_7 ),
        .Q(\alu1/div/rem [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[5] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[7]_i_1__0_n_6 ),
        .Q(\alu1/div/rem [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[6] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[7]_i_1__0_n_5 ),
        .Q(\alu1/div/rem [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[7] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[7]_i_1__0_n_4 ),
        .Q(\alu1/div/rem [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[8] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[11]_i_1__0_n_7 ),
        .Q(\alu1/div/rem [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/div/rrem/rem_reg[9] 
       (.C(clk),
        .CE(\rem[31]_i_1__0_n_0 ),
        .D(\rem_reg[11]_i_1__0_n_6 ),
        .Q(\alu1/div/rem [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[0] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[0]),
        .Q(\alu1/mul/mul_a [0]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[10] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[10]),
        .Q(\alu1/mul/mul_a [10]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[11] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[11]),
        .Q(\alu1/mul/mul_a [11]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[12] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[12]),
        .Q(\alu1/mul/mul_a [12]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[13] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[13]),
        .Q(\alu1/mul/mul_a [13]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[14] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[14]),
        .Q(\alu1/mul/mul_a [14]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[15] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[15]),
        .Q(\alu1/mul/mul_a [15]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[16] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\mul_a[16]_i_1__0_n_0 ),
        .Q(\alu1/mul/mul_a [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[17] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [17]),
        .Q(\alu1/mul/mul_a [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[18] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [18]),
        .Q(\alu1/mul/mul_a [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[19] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [19]),
        .Q(\alu1/mul/mul_a [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[1] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[1]),
        .Q(\alu1/mul/mul_a [1]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[20] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [20]),
        .Q(\alu1/mul/mul_a [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[21] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [21]),
        .Q(\alu1/mul/mul_a [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[22] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [22]),
        .Q(\alu1/mul/mul_a [22]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[23] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [23]),
        .Q(\alu1/mul/mul_a [23]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[24] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [24]),
        .Q(\alu1/mul/mul_a [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[25] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [25]),
        .Q(\alu1/mul/mul_a [25]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[26] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [26]),
        .Q(\alu1/mul/mul_a [26]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[27] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [27]),
        .Q(\alu1/mul/mul_a [27]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[28] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [28]),
        .Q(\alu1/mul/mul_a [28]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[29] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [29]),
        .Q(\alu1/mul/mul_a [29]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[2] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[2]),
        .Q(\alu1/mul/mul_a [2]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[30] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\alu1/mul_a_i [30]),
        .Q(\alu1/mul/mul_a [30]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mul_a_reg[31] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\mul_a[31]_i_1_n_0 ),
        .Q(\alu1/mul/mul_a [31]),
        .R(\<const0> ));
  FDRE \alu1/mul/mul_a_reg[32] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\mul_a[32]_i_1_n_0 ),
        .Q(\alu1/mul/mul_a [32]),
        .R(\<const0> ));
  FDRE \alu1/mul/mul_a_reg[3] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[3]),
        .Q(\alu1/mul/mul_a [3]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[4] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[4]),
        .Q(\alu1/mul/mul_a [4]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[5] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[5]),
        .Q(\alu1/mul/mul_a [5]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[6] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[6]),
        .Q(\alu1/mul/mul_a [6]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[7] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[7]),
        .Q(\alu1/mul/mul_a [7]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[8] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[8]),
        .Q(\alu1/mul/mul_a [8]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_a_reg[9] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(a1bus_0[9]),
        .Q(\alu1/mul/mul_a [9]),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[0] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[0]),
        .Q(\alu1/mul/mul_b_reg_n_0_[0] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[10] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[10]),
        .Q(\alu1/mul/mul_b_reg_n_0_[10] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[11] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[11]),
        .Q(\alu1/mul/mul_b_reg_n_0_[11] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[12] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[12]),
        .Q(\alu1/mul/mul_b_reg_n_0_[12] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[13] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[13]),
        .Q(\alu1/mul/mul_b_reg_n_0_[13] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[14] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[14]),
        .Q(\alu1/mul/mul_b_reg_n_0_[14] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[15] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[15]),
        .Q(\alu1/mul/mul_b_reg_n_0_[15] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[16] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[16]),
        .Q(\alu1/mul/mul_b_reg_n_0_[16] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[17] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[17]),
        .Q(\alu1/mul/mul_b_reg_n_0_[17] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[18] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[18]),
        .Q(\alu1/mul/mul_b_reg_n_0_[18] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[19] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[19]),
        .Q(\alu1/mul/mul_b_reg_n_0_[19] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[1] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[1]),
        .Q(\alu1/mul/mul_b_reg_n_0_[1] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[20] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[20]),
        .Q(\alu1/mul/mul_b_reg_n_0_[20] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[21] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[21]),
        .Q(\alu1/mul/mul_b_reg_n_0_[21] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[22] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[22]),
        .Q(\alu1/mul/mul_b_reg_n_0_[22] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[23] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[23]),
        .Q(\alu1/mul/mul_b_reg_n_0_[23] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[24] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[24]),
        .Q(\alu1/mul/mul_b_reg_n_0_[24] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[25] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[25]),
        .Q(\alu1/mul/mul_b_reg_n_0_[25] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[26] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[26]),
        .Q(\alu1/mul/mul_b_reg_n_0_[26] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[27] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[27]),
        .Q(\alu1/mul/mul_b_reg_n_0_[27] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[28] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[28]),
        .Q(\alu1/mul/mul_b_reg_n_0_[28] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[29] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[29]),
        .Q(\alu1/mul/mul_b_reg_n_0_[29] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[2] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[2]),
        .Q(\alu1/mul/mul_b_reg_n_0_[2] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[30] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[30]),
        .Q(\alu1/mul/mul_b_reg_n_0_[30] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[31] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\mul_b[31]_i_1__0_n_0 ),
        .Q(\alu1/mul/mul_b_reg_n_0_[31] ),
        .R(\<const0> ));
  FDRE \alu1/mul/mul_b_reg[32] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(\mul_b[32]_i_1__0_n_0 ),
        .Q(\alu1/mul/mul_b_reg_n_0_[32] ),
        .R(\<const0> ));
  FDRE \alu1/mul/mul_b_reg[3] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[3]),
        .Q(\alu1/mul/mul_b_reg_n_0_[3] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[4] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[4]),
        .Q(\alu1/mul/mul_b_reg_n_0_[4] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[5] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[5]),
        .Q(\alu1/mul/mul_b_reg_n_0_[5] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[6] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[6]),
        .Q(\alu1/mul/mul_b_reg_n_0_[6] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[7] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[7]),
        .Q(\alu1/mul/mul_b_reg_n_0_[7] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[8] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[8]),
        .Q(\alu1/mul/mul_b_reg_n_0_[8] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_b_reg[9] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(b1bus_0[9]),
        .Q(\alu1/mul/mul_b_reg_n_0_[9] ),
        .R(\mul_a[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mul_rslt_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\alu1/mul/mul_rslt0 ),
        .Q(\alu1/mul/mul_rslt ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \alu1/mul/mulh_reg[0] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[16]),
        .Q(\alu1/mul/mulh [0]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[10] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[26]),
        .Q(\alu1/mul/mulh [10]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[11] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[27]),
        .Q(\alu1/mul/mulh [11]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[12] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[28]),
        .Q(\alu1/mul/mulh [12]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[13] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[29]),
        .Q(\alu1/mul/mulh [13]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[14] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[30]),
        .Q(\alu1/mul/mulh [14]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[15] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[31]),
        .Q(\alu1/mul/mulh [15]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[1] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[17]),
        .Q(\alu1/mul/mulh [1]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[2] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[18]),
        .Q(\alu1/mul/mulh [2]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[3] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[19]),
        .Q(\alu1/mul/mulh [3]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[4] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[20]),
        .Q(\alu1/mul/mulh [4]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[5] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[21]),
        .Q(\alu1/mul/mulh [5]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[6] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[22]),
        .Q(\alu1/mul/mulh [6]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[7] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[23]),
        .Q(\alu1/mul/mulh [7]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[8] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[24]),
        .Q(\alu1/mul/mulh [8]),
        .R(\mulh[15]_i_1__0_n_0 ));
  FDRE \alu1/mul/mulh_reg[9] 
       (.C(clk),
        .CE(\alu1/mul/mul_b ),
        .D(niss_dsp_c1[25]),
        .Q(\alu1/mul/mulh [9]),
        .R(\mulh[15]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_29 
       (.I0(a0bus_0[11]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[11]),
        .O(\art/add/rgf_c0bus_wb[11]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_30 
       (.I0(a0bus_0[10]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[10]),
        .O(\art/add/rgf_c0bus_wb[11]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_31 
       (.I0(a0bus_0[9]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[9]),
        .O(\art/add/rgf_c0bus_wb[11]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[11]_i_32 
       (.I0(a0bus_0[8]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[8]),
        .O(\art/add/rgf_c0bus_wb[11]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_29 
       (.I0(a0bus_0[15]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[15]),
        .O(\art/add/rgf_c0bus_wb[15]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_30 
       (.I0(a0bus_0[14]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[14]),
        .O(\art/add/rgf_c0bus_wb[15]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_31 
       (.I0(a0bus_0[13]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[13]),
        .O(\art/add/rgf_c0bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[15]_i_32 
       (.I0(a0bus_0[12]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[12]),
        .O(\art/add/rgf_c0bus_wb[15]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[19]_i_28 
       (.I0(\alu0/mul_a_i [18]),
        .I1(b0bus_0[18]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[19]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[19]_i_29 
       (.I0(\alu0/mul_a_i [17]),
        .I1(b0bus_0[17]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[19]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \art/add/rgf_c0bus_wb[19]_i_30 
       (.I0(\alu0/asr0 ),
        .I1(\alu0/art/add/p_0_in ),
        .O(\art/add/rgf_c0bus_wb[19]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[23]_i_38 
       (.I0(\alu0/mul_a_i [21]),
        .I1(b0bus_0[21]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[23]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[23]_i_39 
       (.I0(\alu0/mul_a_i [20]),
        .I1(b0bus_0[20]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[23]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[27]_i_40 
       (.I0(\alu0/mul_a_i [27]),
        .I1(b0bus_0[27]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[27]_i_40_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[27]_i_41 
       (.I0(\alu0/mul_a_i [26]),
        .I1(b0bus_0[26]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[27]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[29]_i_29 
       (.I0(\alu0/mul_a_i [30]),
        .I1(b0bus_0[30]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[29]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c0bus_wb[29]_i_30 
       (.I0(\alu0/mul_a_i [29]),
        .I1(b0bus_0[29]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c0bus_wb[29]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_23 
       (.I0(a0bus_0[3]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c0bus_wb[3]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_24 
       (.I0(a0bus_0[2]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c0bus_wb[3]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_25 
       (.I0(a0bus_0[1]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c0bus_wb[3]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[3]_i_26 
       (.I0(a0bus_0[0]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c0bus_wb[3]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c0bus_wb[7]_i_30 
       (.I0(a0bus_0[7]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[7]),
        .O(\art/add/rgf_c0bus_wb[7]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[7]_i_31 
       (.I0(a0bus_0[6]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(\bbus_o[6]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c0bus_wb[7]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[7]_i_32 
       (.I0(a0bus_0[5]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c0bus_wb[7]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c0bus_wb[7]_i_33 
       (.I0(a0bus_0[4]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c0bus_wb[7]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_26 
       (.I0(a1bus_0[11]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[11]),
        .O(\art/add/rgf_c1bus_wb[11]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_27 
       (.I0(a1bus_0[10]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[10]),
        .O(\art/add/rgf_c1bus_wb[11]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_28 
       (.I0(a1bus_0[9]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[9]),
        .O(\art/add/rgf_c1bus_wb[11]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[11]_i_29 
       (.I0(a1bus_0[8]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[8]),
        .O(\art/add/rgf_c1bus_wb[11]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[19]_i_23 
       (.I0(\alu1/mul_a_i [19]),
        .I1(b1bus_0[19]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[19]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[19]_i_24 
       (.I0(\alu1/mul_a_i [18]),
        .I1(b1bus_0[18]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[19]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[19]_i_25 
       (.I0(\alu1/mul_a_i [17]),
        .I1(b1bus_0[17]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[19]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h1E)) 
    \art/add/rgf_c1bus_wb[19]_i_26 
       (.I0(\mul_a[16]_i_1__0_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\alu1/art/add/p_0_in ),
        .O(\art/add/rgf_c1bus_wb[19]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_35 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[15]),
        .O(\art/add/rgf_c1bus_wb[19]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_36 
       (.I0(a1bus_0[14]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[14]),
        .O(\art/add/rgf_c1bus_wb[19]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_37 
       (.I0(a1bus_0[13]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[13]),
        .O(\art/add/rgf_c1bus_wb[19]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[19]_i_38 
       (.I0(a1bus_0[12]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[12]),
        .O(\art/add/rgf_c1bus_wb[19]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[23]_i_27 
       (.I0(\alu1/mul_a_i [22]),
        .I1(b1bus_0[22]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[23]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[23]_i_28 
       (.I0(\alu1/mul_a_i [21]),
        .I1(b1bus_0[21]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[23]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[23]_i_29 
       (.I0(\alu1/mul_a_i [20]),
        .I1(b1bus_0[20]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[23]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_21 
       (.I0(\alu1/mul_a_i [27]),
        .I1(b1bus_0[27]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_22 
       (.I0(\alu1/mul_a_i [26]),
        .I1(b1bus_0[26]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_23 
       (.I0(\alu1/mul_a_i [25]),
        .I1(b1bus_0[25]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[27]_i_24 
       (.I0(\alu1/mul_a_i [24]),
        .I1(b1bus_0[24]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[27]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \art/add/rgf_c1bus_wb[31]_i_29 
       (.I0(\alu1/mul_a_i [31]),
        .I1(\alu1/art/p_0_in__0 ),
        .O(\art/add/rgf_c1bus_wb[31]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[31]_i_30 
       (.I0(\alu1/mul_a_i [30]),
        .I1(b1bus_0[30]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[31]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[31]_i_31 
       (.I0(\alu1/mul_a_i [29]),
        .I1(b1bus_0[29]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[31]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h69AA)) 
    \art/add/rgf_c1bus_wb[31]_i_32 
       (.I0(\alu1/mul_a_i [28]),
        .I1(b1bus_0[28]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\art/add/rgf_c1bus_wb[31]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_27 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c1bus_wb[3]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_28 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c1bus_wb[3]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_29 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c1bus_wb[3]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[3]_i_30 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c1bus_wb[3]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/rgf_c1bus_wb[7]_i_31 
       (.I0(a1bus_0[7]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[7]),
        .O(\art/add/rgf_c1bus_wb[7]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[7]_i_32 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c1bus_wb[7]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[7]_i_33 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\art/add/rgf_c1bus_wb[7]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h96)) 
    \art/add/rgf_c1bus_wb[7]_i_34 
       (.I0(a1bus_0[4]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\art/add/rgf_c1bus_wb[7]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \art/add/sr[6]_i_29 
       (.I0(\alu1/mul_a_i [31]),
        .I1(\alu1/art/p_0_in__0 ),
        .O(\art/add/sr[6]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[0]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[0]),
        .O(badr[0]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[0]_INST_0_i_10 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [0]),
        .O(\rgf/a0bus_sr [0]));
  LUT6 #(
    .INIT(64'h4445555544444444)) 
    \badr[0]_INST_0_i_25 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_77_n_0 ),
        .I2(\fch/ir0 [15]),
        .I3(\badr[31]_INST_0_i_78_n_0 ),
        .I4(\badr[31]_INST_0_i_79_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .O(\badr[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [0]),
        .I5(\rgf/ivec/iv [0]),
        .O(\badr[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [0]),
        .O(\badr[0]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[0]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [0]),
        .O(\badr[0]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [0]),
        .O(\badr[0]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[0]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [0]),
        .O(\badr[0]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [0]),
        .I5(\rgf/ivec/iv [0]),
        .O(\badr[0]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[10]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[10]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[10]),
        .O(badr[10]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[10]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [10]),
        .O(\rgf/a0bus_sr [10]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [10]),
        .O(\badr[10]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [10]),
        .O(\badr[10]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [10]),
        .I5(\rgf/ivec/iv [10]),
        .O(\badr[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [10]),
        .O(\badr[10]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[10]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [10]),
        .O(\badr[10]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [10]),
        .O(\badr[10]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[10]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [10]),
        .O(\badr[10]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[10]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [10]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [10]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [10]),
        .I5(\rgf/ivec/iv [10]),
        .O(\badr[10]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[11]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[11]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[11]),
        .O(badr[11]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[11]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [11]),
        .O(\rgf/a0bus_sr [11]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [11]),
        .O(\badr[11]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [11]),
        .O(\badr[11]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [11]),
        .I5(\rgf/ivec/iv [11]),
        .O(\badr[11]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [11]),
        .O(\badr[11]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[11]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [11]),
        .O(\badr[11]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [11]),
        .O(\badr[11]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[11]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [11]),
        .O(\badr[11]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[11]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [11]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [11]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [11]),
        .I5(\rgf/ivec/iv [11]),
        .O(\badr[11]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[12]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[12]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[12]),
        .O(badr[12]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[12]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [12]),
        .O(\rgf/a0bus_sr [12]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [12]),
        .O(\badr[12]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [12]),
        .O(\badr[12]_INST_0_i_21_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[12]_INST_0_i_29 
       (.CI(\badr[8]_INST_0_i_29_n_0 ),
        .CO({\badr[12]_INST_0_i_29_n_0 ,\badr[12]_INST_0_i_29_n_1 ,\badr[12]_INST_0_i_29_n_2 ,\badr[12]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [11:8]),
        .O(\rgf/sptr/data3 [12:9]),
        .S({\badr[12]_INST_0_i_46_n_0 ,\badr[12]_INST_0_i_47_n_0 ,\badr[12]_INST_0_i_48_n_0 ,\badr[12]_INST_0_i_49_n_0 }));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [12]),
        .I5(\rgf/ivec/iv [12]),
        .O(\badr[12]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_46 
       (.I0(\rgf/sptr/sp [11]),
        .I1(\rgf/sptr/sp [12]),
        .O(\badr[12]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_47 
       (.I0(\rgf/sptr/sp [10]),
        .I1(\rgf/sptr/sp [11]),
        .O(\badr[12]_INST_0_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_48 
       (.I0(\rgf/sptr/sp [9]),
        .I1(\rgf/sptr/sp [10]),
        .O(\badr[12]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_49 
       (.I0(\rgf/sptr/sp [8]),
        .I1(\rgf/sptr/sp [9]),
        .O(\badr[12]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [12]),
        .O(\badr[12]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[12]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [12]),
        .O(\badr[12]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [12]),
        .O(\badr[12]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[12]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [12]),
        .O(\badr[12]_INST_0_i_53_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[12]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [12]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [12]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [12]),
        .I5(\rgf/ivec/iv [12]),
        .O(\badr[12]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[13]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[13]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[13]),
        .O(badr[13]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[13]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [13]),
        .O(\rgf/a0bus_sr [13]));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[13]_INST_0_i_15 
       (.I0(\badr[15]_INST_0_i_14_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .O(\badr[13]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [13]),
        .O(\badr[13]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [13]),
        .O(\badr[13]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [13]),
        .I5(\rgf/ivec/iv [13]),
        .O(\badr[13]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \badr[13]_INST_0_i_46 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [8]),
        .O(\badr[13]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [13]),
        .O(\badr[13]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[13]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [13]),
        .O(\badr[13]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [13]),
        .O(\badr[13]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[13]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [13]),
        .O(\badr[13]_INST_0_i_52_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[13]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [13]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [13]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [13]),
        .I5(\rgf/ivec/iv [13]),
        .O(\badr[13]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[14]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[14]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[14]),
        .O(badr[14]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[14]_INST_0_i_10 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [14]),
        .O(\rgf/a0bus_sr [14]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [14]),
        .O(\badr[14]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[14]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [14]),
        .O(\badr[14]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [14]),
        .O(\badr[14]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[14]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [14]),
        .O(\badr[14]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [14]),
        .I5(\rgf/ivec/iv [14]),
        .O(\badr[14]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[15]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[15]),
        .O(badr[15]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_100 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [15]),
        .O(\badr[15]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_103 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [15]),
        .O(\badr[15]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[15]_INST_0_i_104 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [15]),
        .O(\badr[15]_INST_0_i_104_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[15]_INST_0_i_11 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [15]),
        .O(\rgf/a0bus_sr [15]));
  LUT6 #(
    .INIT(64'hFFFF7FFFFFDFFFFF)) 
    \badr[15]_INST_0_i_113 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [6]),
        .O(\badr[15]_INST_0_i_113_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[15]_INST_0_i_114 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [6]),
        .O(\badr[15]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000008FF)) 
    \badr[15]_INST_0_i_115 
       (.I0(\niss_dsp_b1[1]_INST_0_i_8_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [15]),
        .I3(\badr[15]_INST_0_i_133_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\badr[15]_INST_0_i_115_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000DA)) 
    \badr[15]_INST_0_i_116 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [1]),
        .I3(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I4(\fch/ir1 [2]),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\badr[15]_INST_0_i_116_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA8AAA8AAAA)) 
    \badr[15]_INST_0_i_117 
       (.I0(\sr[15]_i_6_n_0 ),
        .I1(\badr[15]_INST_0_i_134_n_0 ),
        .I2(\badr[15]_INST_0_i_135_n_0 ),
        .I3(\badr[15]_INST_0_i_136_n_0 ),
        .I4(\fch/ir1 [10]),
        .I5(\badr[15]_INST_0_i_137_n_0 ),
        .O(\badr[15]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000004F)) 
    \badr[15]_INST_0_i_118 
       (.I0(\badr[15]_INST_0_i_138_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_29_n_0 ),
        .I2(\badr[31]_INST_0_i_165_n_0 ),
        .I3(\badr[15]_INST_0_i_139_n_0 ),
        .I4(\badr[15]_INST_0_i_140_n_0 ),
        .I5(\badr[15]_INST_0_i_141_n_0 ),
        .O(\badr[15]_INST_0_i_118_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBFFFFFF3FFFFF)) 
    \badr[15]_INST_0_i_119 
       (.I0(\badr[15]_INST_0_i_142_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [10]),
        .O(\badr[15]_INST_0_i_119_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \badr[15]_INST_0_i_120 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .O(\badr[15]_INST_0_i_120_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \badr[15]_INST_0_i_121 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_121_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000005D50)) 
    \badr[15]_INST_0_i_122 
       (.I0(\badr[15]_INST_0_i_143_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_74_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\fch/ir1 [15]),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\badr[15]_INST_0_i_122_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF7FFF)) 
    \badr[15]_INST_0_i_123 
       (.I0(\niss_dsp_a1[15]_INST_0_i_17_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I2(\fch/ir1 [0]),
        .I3(fch_irq_req),
        .I4(\fch/ir1 [10]),
        .I5(\bdatw[9]_INST_0_i_10_n_0 ),
        .O(\badr[15]_INST_0_i_123_n_0 ));
  LUT5 #(
    .INIT(32'h0000007F)) 
    \badr[15]_INST_0_i_124 
       (.I0(\badr[15]_INST_0_i_144_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [0]),
        .I3(\badr[15]_INST_0_i_145_n_0 ),
        .I4(\badr[15]_INST_0_i_146_n_0 ),
        .O(\badr[15]_INST_0_i_124_n_0 ));
  LUT6 #(
    .INIT(64'hFFD0F0F0D0D0D0D0)) 
    \badr[15]_INST_0_i_125 
       (.I0(\badr[15]_INST_0_i_147_n_0 ),
        .I1(\badr[15]_INST_0_i_148_n_0 ),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [6]),
        .I5(\badr[31]_INST_0_i_165_n_0 ),
        .O(\badr[15]_INST_0_i_125_n_0 ));
  LUT6 #(
    .INIT(64'h8080808080808880)) 
    \badr[15]_INST_0_i_126 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [12]),
        .I2(\badr[15]_INST_0_i_149_n_0 ),
        .I3(\fch/ir1 [8]),
        .I4(\stat[1]_i_22_n_0 ),
        .I5(\badr[15]_INST_0_i_150_n_0 ),
        .O(\badr[15]_INST_0_i_126_n_0 ));
  LUT4 #(
    .INIT(16'h9666)) 
    \badr[15]_INST_0_i_127 
       (.I0(\fch/ir1 [11]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [7]),
        .O(\badr[15]_INST_0_i_127_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \badr[15]_INST_0_i_128 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [8]),
        .O(\badr[15]_INST_0_i_128_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDF0F0FFFFFFFF)) 
    \badr[15]_INST_0_i_129 
       (.I0(\badr[31]_INST_0_i_75_n_0 ),
        .I1(\badr[31]_INST_0_i_74_n_0 ),
        .I2(stat[2]),
        .I3(\fch/ir0 [11]),
        .I4(\badr[31]_INST_0_i_73_n_0 ),
        .I5(ctl_sela0),
        .O(\badr[15]_INST_0_i_129_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FFA2)) 
    \badr[15]_INST_0_i_130 
       (.I0(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I1(\badr[31]_INST_0_i_86_n_0 ),
        .I2(\badr[31]_INST_0_i_87_n_0 ),
        .I3(\badr[31]_INST_0_i_88_n_0 ),
        .I4(stat[2]),
        .I5(\badr[31]_INST_0_i_89_n_0 ),
        .O(ctl_sela0_rn));
  LUT6 #(
    .INIT(64'h5554555554545454)) 
    \badr[15]_INST_0_i_131 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_82_n_0 ),
        .I2(\badr[31]_INST_0_i_83_n_0 ),
        .I3(\badr[31]_INST_0_i_84_n_0 ),
        .I4(\badr[31]_INST_0_i_85_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_131_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDF0F0FFFFFFFF)) 
    \badr[15]_INST_0_i_132 
       (.I0(\badr[31]_INST_0_i_75_n_0 ),
        .I1(\badr[31]_INST_0_i_74_n_0 ),
        .I2(stat[2]),
        .I3(\fch/ir0 [11]),
        .I4(\badr[31]_INST_0_i_73_n_0 ),
        .I5(ctl_sela0),
        .O(\badr[15]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFEF)) 
    \badr[15]_INST_0_i_133 
       (.I0(\bcmd[1]_INST_0_i_14_n_0 ),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [0]),
        .O(\badr[15]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'h0080A000A0008808)) 
    \badr[15]_INST_0_i_134 
       (.I0(\bdatw[31]_INST_0_i_113_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [5]),
        .O(\badr[15]_INST_0_i_134_n_0 ));
  LUT6 #(
    .INIT(64'h4555455500000500)) 
    \badr[15]_INST_0_i_135 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(div_crdy1),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [4]),
        .O(\badr[15]_INST_0_i_135_n_0 ));
  LUT6 #(
    .INIT(64'hA2080002A0000000)) 
    \badr[15]_INST_0_i_136 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [1]),
        .O(\badr[15]_INST_0_i_136_n_0 ));
  LUT6 #(
    .INIT(64'h0140FD7F0444F777)) 
    \badr[15]_INST_0_i_137 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [7]),
        .O(\badr[15]_INST_0_i_137_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[15]_INST_0_i_138 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [1]),
        .O(\badr[15]_INST_0_i_138_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFAE00AE)) 
    \badr[15]_INST_0_i_139 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [4]),
        .I5(\stat[1]_i_22_n_0 ),
        .O(\badr[15]_INST_0_i_139_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \badr[15]_INST_0_i_14 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\badr[15]_INST_0_i_47_n_0 ),
        .I2(\badr[15]_INST_0_i_48_n_0 ),
        .I3(\badr[31]_INST_0_i_64_n_0 ),
        .I4(\fch/ir1 [9]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h5000000045004500)) 
    \badr[15]_INST_0_i_140 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(div_crdy1),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'h0404000404000000)) 
    \badr[15]_INST_0_i_141 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(div_crdy1),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [4]),
        .O(\badr[15]_INST_0_i_141_n_0 ));
  LUT6 #(
    .INIT(64'hDFFBFFFFFFFFFFFF)) 
    \badr[15]_INST_0_i_142 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [0]),
        .O(\badr[15]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \badr[15]_INST_0_i_143 
       (.I0(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [0]),
        .I5(\fch/ir1 [3]),
        .O(\badr[15]_INST_0_i_143_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[15]_INST_0_i_144 
       (.I0(\fch/ir1 [9]),
        .I1(div_crdy1),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\badr[15]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'h1001000000010000)) 
    \badr[15]_INST_0_i_145 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(div_crdy1),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [6]),
        .O(\badr[15]_INST_0_i_145_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF8A008A)) 
    \badr[15]_INST_0_i_146 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [3]),
        .I5(\stat[1]_i_22_n_0 ),
        .O(\badr[15]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFFFFFDFDFDFDF)) 
    \badr[15]_INST_0_i_147 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [8]),
        .O(\badr[15]_INST_0_i_147_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \badr[15]_INST_0_i_148 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(div_crdy1),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .O(\badr[15]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'hF4FF444444444444)) 
    \badr[15]_INST_0_i_149 
       (.I0(\fch/ir1 [10]),
        .I1(\badr[15]_INST_0_i_151_n_0 ),
        .I2(\fch/ir1 [6]),
        .I3(\bcmd[1]_INST_0_i_26_n_0 ),
        .I4(\fch/ir1 [3]),
        .I5(\niss_dsp_b1[5]_INST_0_i_65_n_0 ),
        .O(\badr[15]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h5454545544444444)) 
    \badr[15]_INST_0_i_15 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\badr[15]_INST_0_i_49_n_0 ),
        .I2(\badr[15]_INST_0_i_50_n_0 ),
        .I3(\badr[15]_INST_0_i_51_n_0 ),
        .I4(\badr[15]_INST_0_i_52_n_0 ),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\badr[15]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCFFF1F0FFF514FF5)) 
    \badr[15]_INST_0_i_150 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [5]),
        .O(\badr[15]_INST_0_i_150_n_0 ));
  LUT6 #(
    .INIT(64'hF1F4F8FCE0B07030)) 
    \badr[15]_INST_0_i_151 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [0]),
        .O(\badr[15]_INST_0_i_151_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_28 
       (.I0(\badr[15]_INST_0_i_14_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_sel_cr [1]));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_29 
       (.I0(\badr[31]_INST_0_i_58_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .O(\badr[15]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[15]_INST_0_i_44 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sel_cr [5]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_45 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sel_cr [2]));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_46 
       (.I0(\badr[31]_INST_0_i_58_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sel_cr [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFF1F110000)) 
    \badr[15]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_113_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I3(\badr[15]_INST_0_i_114_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\badr[15]_INST_0_i_115_n_0 ),
        .O(\badr[15]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \badr[15]_INST_0_i_48 
       (.I0(\fch/ir1 [15]),
        .I1(\badr[15]_INST_0_i_116_n_0 ),
        .I2(\badr[15]_INST_0_i_117_n_0 ),
        .I3(\badr[15]_INST_0_i_118_n_0 ),
        .I4(\badr[31]_INST_0_i_102_n_0 ),
        .I5(ctl_fetch1_fl_i_16_n_0),
        .O(\badr[15]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF47440000)) 
    \badr[15]_INST_0_i_49 
       (.I0(\badr[15]_INST_0_i_119_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\badr[15]_INST_0_i_120_n_0 ),
        .I3(\badr[15]_INST_0_i_121_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I5(\badr[15]_INST_0_i_122_n_0 ),
        .O(\badr[15]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_5 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_sel_cr [0]));
  LUT5 #(
    .INIT(32'hAEAEFFAE)) 
    \badr[15]_INST_0_i_50 
       (.I0(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_24_n_0 ),
        .I2(\badr[15]_INST_0_i_123_n_0 ),
        .I3(\fch/ir1 [8]),
        .I4(\badr[31]_INST_0_i_64_n_0 ),
        .O(\badr[15]_INST_0_i_50_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[15]_INST_0_i_51 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [14]),
        .O(\badr[15]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h005DFFFF005D0000)) 
    \badr[15]_INST_0_i_52 
       (.I0(\badr[31]_INST_0_i_102_n_0 ),
        .I1(\badr[15]_INST_0_i_124_n_0 ),
        .I2(\badr[15]_INST_0_i_125_n_0 ),
        .I3(\badr[15]_INST_0_i_126_n_0 ),
        .I4(\fch/ir1 [13]),
        .I5(\badr[15]_INST_0_i_127_n_0 ),
        .O(\badr[15]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_8 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [15]),
        .I5(\rgf/ivec/iv [15]),
        .O(\badr[15]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[15]_INST_0_i_99 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [15]),
        .O(\badr[15]_INST_0_i_99_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[16]_INST_0 
       (.I0(a1bus_0[16]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[16]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [0]),
        .O(badr[16]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[16]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [16]),
        .I1(\rgf/sptr/data3 [16]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [16]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [0]),
        .O(\badr[16]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [0]),
        .O(\badr[16]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\badr[16]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [0]),
        .O(\badr[16]_INST_0_i_19_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[16]_INST_0_i_21 
       (.CI(\badr[12]_INST_0_i_29_n_0 ),
        .CO({\badr[16]_INST_0_i_21_n_0 ,\badr[16]_INST_0_i_21_n_1 ,\badr[16]_INST_0_i_21_n_2 ,\badr[16]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [15:12]),
        .O(\rgf/sptr/data3 [16:13]),
        .S({\badr[16]_INST_0_i_30_n_0 ,\badr[16]_INST_0_i_31_n_0 ,\badr[16]_INST_0_i_32_n_0 ,\badr[16]_INST_0_i_33_n_0 }));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [0]),
        .O(\badr[16]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [0]),
        .O(\badr[16]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [0]),
        .O(\badr[16]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [0]),
        .O(\badr[16]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\badr[16]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[16]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [0]),
        .O(\badr[16]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [0]),
        .O(\badr[16]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[16]_INST_0_i_29 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [0]),
        .O(\badr[16]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[16]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [16]),
        .O(\badr[16]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_30 
       (.I0(\rgf/sptr/sp [15]),
        .I1(\rgf/sptr/sp [16]),
        .O(\badr[16]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_31 
       (.I0(\rgf/sptr/sp [14]),
        .I1(\rgf/sptr/sp [15]),
        .O(\badr[16]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_32 
       (.I0(\rgf/sptr/sp [13]),
        .I1(\rgf/sptr/sp [14]),
        .O(\badr[16]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_33 
       (.I0(\rgf/sptr/sp [12]),
        .I1(\rgf/sptr/sp [13]),
        .O(\badr[16]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[16]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [16]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [16]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [16]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[16]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [16]),
        .O(\badr[16]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[17]_INST_0 
       (.I0(a1bus_0[17]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[17]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [1]),
        .O(badr[17]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[17]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [17]),
        .I1(\rgf/sptr/data3 [17]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [17]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [1]),
        .O(\badr[17]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [1]),
        .O(\badr[17]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\badr[17]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\badr[17]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [1]),
        .O(\badr[17]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [1]),
        .O(\badr[17]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [1]),
        .O(\badr[17]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [1]),
        .O(\badr[17]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\badr[17]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[17]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\badr[17]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [1]),
        .O(\badr[17]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[17]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [1]),
        .O(\badr[17]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[17]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [17]),
        .O(\badr[17]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[17]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [17]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [17]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [17]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[17]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [17]),
        .O(\badr[17]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[18]_INST_0 
       (.I0(a1bus_0[18]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[18]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [2]),
        .O(badr[18]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[18]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [18]),
        .I1(\rgf/sptr/data3 [18]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [18]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [2]),
        .O(\badr[18]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [2]),
        .O(\badr[18]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\badr[18]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [2]),
        .O(\badr[18]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [2]),
        .O(\badr[18]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [2]),
        .O(\badr[18]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [2]),
        .O(\badr[18]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [2]),
        .O(\badr[18]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\badr[18]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[18]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [2]),
        .O(\badr[18]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [2]),
        .O(\badr[18]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[18]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [2]),
        .O(\badr[18]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[18]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [18]),
        .O(\badr[18]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[18]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [18]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [18]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [18]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[18]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [18]),
        .O(\badr[18]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[19]_INST_0 
       (.I0(a1bus_0[19]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[19]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [3]),
        .O(badr[19]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[19]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [19]),
        .I1(\rgf/sptr/data3 [19]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [19]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [3]),
        .O(\badr[19]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [3]),
        .O(\badr[19]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\badr[19]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\badr[19]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [3]),
        .O(\badr[19]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [3]),
        .O(\badr[19]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [3]),
        .O(\badr[19]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [3]),
        .O(\badr[19]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\badr[19]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[19]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\badr[19]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [3]),
        .O(\badr[19]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[19]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [3]),
        .O(\badr[19]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[19]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [19]),
        .O(\badr[19]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[19]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [19]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [19]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [19]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[19]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [19]),
        .O(\badr[19]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[1]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[1]),
        .O(badr[1]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[1]_INST_0_i_10 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [1]),
        .O(\rgf/a0bus_sr [1]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [1]),
        .O(\badr[1]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[1]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [1]),
        .O(\badr[1]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [1]),
        .O(\badr[1]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[1]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [1]),
        .O(\badr[1]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [1]),
        .I5(\rgf/ivec/iv [1]),
        .O(\badr[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[20]_INST_0 
       (.I0(a1bus_0[20]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[20]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [4]),
        .O(badr[20]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[20]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [20]),
        .I1(\rgf/sptr/data3 [20]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [20]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [4]),
        .O(\badr[20]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [4]),
        .O(\badr[20]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\badr[20]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [4]),
        .O(\badr[20]_INST_0_i_19_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[20]_INST_0_i_21 
       (.CI(\badr[16]_INST_0_i_21_n_0 ),
        .CO({\badr[20]_INST_0_i_21_n_0 ,\badr[20]_INST_0_i_21_n_1 ,\badr[20]_INST_0_i_21_n_2 ,\badr[20]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [19:16]),
        .O(\rgf/sptr/data3 [20:17]),
        .S({\badr[20]_INST_0_i_30_n_0 ,\badr[20]_INST_0_i_31_n_0 ,\badr[20]_INST_0_i_32_n_0 ,\badr[20]_INST_0_i_33_n_0 }));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [4]),
        .O(\badr[20]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [4]),
        .O(\badr[20]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [4]),
        .O(\badr[20]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [4]),
        .O(\badr[20]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\badr[20]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[20]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [4]),
        .O(\badr[20]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [4]),
        .O(\badr[20]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[20]_INST_0_i_29 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [4]),
        .O(\badr[20]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[20]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [20]),
        .O(\badr[20]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_30 
       (.I0(\rgf/sptr/sp [19]),
        .I1(\rgf/sptr/sp [20]),
        .O(\badr[20]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_31 
       (.I0(\rgf/sptr/sp [18]),
        .I1(\rgf/sptr/sp [19]),
        .O(\badr[20]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_32 
       (.I0(\rgf/sptr/sp [17]),
        .I1(\rgf/sptr/sp [18]),
        .O(\badr[20]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_33 
       (.I0(\rgf/sptr/sp [16]),
        .I1(\rgf/sptr/sp [17]),
        .O(\badr[20]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[20]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [20]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [20]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [20]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[20]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [20]),
        .O(\badr[20]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFE2000000E200)) 
    \badr[21]_INST_0 
       (.I0(a1bus_0[21]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(a0bus_0[21]),
        .I3(\badr[31]_INST_0_i_1_n_0 ),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [5]),
        .O(badr[21]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[21]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [21]),
        .I1(\rgf/sptr/data3 [21]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [21]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [5]),
        .O(\badr[21]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [5]),
        .O(\badr[21]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\badr[21]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [5]),
        .O(\badr[21]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [5]),
        .O(\badr[21]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [5]),
        .O(\badr[21]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [5]),
        .O(\badr[21]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [5]),
        .O(\badr[21]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\badr[21]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[21]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [5]),
        .O(\badr[21]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [5]),
        .O(\badr[21]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[21]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [5]),
        .O(\badr[21]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[21]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [21]),
        .O(\badr[21]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[21]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [21]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [21]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [21]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[21]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [21]),
        .O(\badr[21]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[22]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[22]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[22]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [6]),
        .O(badr[22]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[22]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [22]),
        .I1(\rgf/sptr/data3 [22]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [22]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [6]),
        .O(\badr[22]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [6]),
        .O(\badr[22]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [6]),
        .O(\badr[22]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [6]),
        .O(\badr[22]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [6]),
        .O(\badr[22]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [6]),
        .O(\badr[22]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [6]),
        .O(\badr[22]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [6]),
        .O(\badr[22]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [6]),
        .O(\badr[22]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[22]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [6]),
        .O(\badr[22]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [6]),
        .O(\badr[22]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[22]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [6]),
        .O(\badr[22]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[22]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [22]),
        .O(\badr[22]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[22]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [22]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [22]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [22]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[22]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [22]),
        .O(\badr[22]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[23]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[23]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[23]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [7]),
        .O(badr[23]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[23]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [23]),
        .I1(\rgf/sptr/data3 [23]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [23]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [7]),
        .O(\badr[23]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [7]),
        .O(\badr[23]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [7]),
        .O(\badr[23]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [7]),
        .O(\badr[23]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [7]),
        .O(\badr[23]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [7]),
        .O(\badr[23]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [7]),
        .O(\badr[23]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [7]),
        .O(\badr[23]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [7]),
        .O(\badr[23]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[23]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [7]),
        .O(\badr[23]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [7]),
        .O(\badr[23]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[23]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [7]),
        .O(\badr[23]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[23]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [23]),
        .O(\badr[23]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[23]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [23]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [23]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [23]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[23]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [23]),
        .O(\badr[23]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[24]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[24]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[24]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [8]),
        .O(badr[24]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[24]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [24]),
        .I1(\rgf/sptr/data3 [24]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [24]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [8]),
        .O(\badr[24]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [8]),
        .O(\badr[24]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [8]),
        .O(\badr[24]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [8]),
        .O(\badr[24]_INST_0_i_19_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[24]_INST_0_i_21 
       (.CI(\badr[20]_INST_0_i_21_n_0 ),
        .CO({\badr[24]_INST_0_i_21_n_0 ,\badr[24]_INST_0_i_21_n_1 ,\badr[24]_INST_0_i_21_n_2 ,\badr[24]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [23:20]),
        .O(\rgf/sptr/data3 [24:21]),
        .S({\badr[24]_INST_0_i_30_n_0 ,\badr[24]_INST_0_i_31_n_0 ,\badr[24]_INST_0_i_32_n_0 ,\badr[24]_INST_0_i_33_n_0 }));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [8]),
        .O(\badr[24]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [8]),
        .O(\badr[24]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [8]),
        .O(\badr[24]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [8]),
        .O(\badr[24]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [8]),
        .O(\badr[24]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[24]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [8]),
        .O(\badr[24]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [8]),
        .O(\badr[24]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[24]_INST_0_i_29 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [8]),
        .O(\badr[24]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[24]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [24]),
        .O(\badr[24]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_30 
       (.I0(\rgf/sptr/sp [23]),
        .I1(\rgf/sptr/sp [24]),
        .O(\badr[24]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_31 
       (.I0(\rgf/sptr/sp [22]),
        .I1(\rgf/sptr/sp [23]),
        .O(\badr[24]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_32 
       (.I0(\rgf/sptr/sp [21]),
        .I1(\rgf/sptr/sp [22]),
        .O(\badr[24]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_33 
       (.I0(\rgf/sptr/sp [20]),
        .I1(\rgf/sptr/sp [21]),
        .O(\badr[24]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[24]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [24]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [24]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [24]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[24]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [24]),
        .O(\badr[24]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[25]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[25]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[25]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [9]),
        .O(badr[25]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[25]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [25]),
        .I1(\rgf/sptr/data3 [25]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [25]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [9]),
        .O(\badr[25]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [9]),
        .O(\badr[25]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [9]),
        .O(\badr[25]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [9]),
        .O(\badr[25]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [9]),
        .O(\badr[25]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [9]),
        .O(\badr[25]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [9]),
        .O(\badr[25]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [9]),
        .O(\badr[25]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [9]),
        .O(\badr[25]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[25]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [9]),
        .O(\badr[25]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [9]),
        .O(\badr[25]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[25]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [9]),
        .O(\badr[25]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[25]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [25]),
        .O(\badr[25]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[25]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [25]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [25]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [25]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[25]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [25]),
        .O(\badr[25]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[26]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[26]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[26]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [10]),
        .O(badr[26]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[26]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [26]),
        .I1(\rgf/sptr/data3 [26]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [26]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [10]),
        .O(\badr[26]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [10]),
        .O(\badr[26]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [10]),
        .O(\badr[26]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [10]),
        .O(\badr[26]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [10]),
        .O(\badr[26]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [10]),
        .O(\badr[26]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [10]),
        .O(\badr[26]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [10]),
        .O(\badr[26]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [10]),
        .O(\badr[26]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[26]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [10]),
        .O(\badr[26]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [10]),
        .O(\badr[26]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[26]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [10]),
        .O(\badr[26]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[26]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [26]),
        .O(\badr[26]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[26]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [26]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [26]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [26]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[26]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [26]),
        .O(\badr[26]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[27]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[27]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[27]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [11]),
        .O(badr[27]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[27]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [27]),
        .I1(\rgf/sptr/data3 [27]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [27]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [11]),
        .O(\badr[27]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [11]),
        .O(\badr[27]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [11]),
        .O(\badr[27]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [11]),
        .O(\badr[27]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [11]),
        .O(\badr[27]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [11]),
        .O(\badr[27]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [11]),
        .O(\badr[27]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [11]),
        .O(\badr[27]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [11]),
        .O(\badr[27]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[27]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [11]),
        .O(\badr[27]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [11]),
        .O(\badr[27]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[27]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [11]),
        .O(\badr[27]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[27]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [27]),
        .O(\badr[27]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[27]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [27]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [27]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [27]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[27]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [27]),
        .O(\badr[27]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[28]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[28]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[28]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [12]),
        .O(badr[28]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[28]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [28]),
        .I1(\rgf/sptr/data3 [28]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [28]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [12]),
        .O(\badr[28]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [12]),
        .O(\badr[28]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [12]),
        .O(\badr[28]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [12]),
        .O(\badr[28]_INST_0_i_19_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[28]_INST_0_i_21 
       (.CI(\badr[24]_INST_0_i_21_n_0 ),
        .CO({\badr[28]_INST_0_i_21_n_0 ,\badr[28]_INST_0_i_21_n_1 ,\badr[28]_INST_0_i_21_n_2 ,\badr[28]_INST_0_i_21_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [27:24]),
        .O(\rgf/sptr/data3 [28:25]),
        .S({\badr[28]_INST_0_i_30_n_0 ,\badr[28]_INST_0_i_31_n_0 ,\badr[28]_INST_0_i_32_n_0 ,\badr[28]_INST_0_i_33_n_0 }));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [12]),
        .O(\badr[28]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [12]),
        .O(\badr[28]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [12]),
        .O(\badr[28]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [12]),
        .O(\badr[28]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [12]),
        .O(\badr[28]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[28]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [12]),
        .O(\badr[28]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [12]),
        .O(\badr[28]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[28]_INST_0_i_29 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [12]),
        .O(\badr[28]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[28]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [28]),
        .O(\badr[28]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_30 
       (.I0(\rgf/sptr/sp [27]),
        .I1(\rgf/sptr/sp [28]),
        .O(\badr[28]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_31 
       (.I0(\rgf/sptr/sp [26]),
        .I1(\rgf/sptr/sp [27]),
        .O(\badr[28]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_32 
       (.I0(\rgf/sptr/sp [25]),
        .I1(\rgf/sptr/sp [26]),
        .O(\badr[28]_INST_0_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_33 
       (.I0(\rgf/sptr/sp [24]),
        .I1(\rgf/sptr/sp [25]),
        .O(\badr[28]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[28]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [28]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [28]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [28]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[28]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [28]),
        .O(\badr[28]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[29]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[29]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[29]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [13]),
        .O(badr[29]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[29]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [29]),
        .I1(\rgf/sptr/data3 [29]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [29]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [13]),
        .O(\badr[29]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [13]),
        .O(\badr[29]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [13]),
        .O(\badr[29]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [13]),
        .O(\badr[29]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [13]),
        .O(\badr[29]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [13]),
        .O(\badr[29]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [13]),
        .O(\badr[29]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [13]),
        .O(\badr[29]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [13]),
        .O(\badr[29]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[29]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [13]),
        .O(\badr[29]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [13]),
        .O(\badr[29]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[29]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [13]),
        .O(\badr[29]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[29]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [29]),
        .O(\badr[29]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[29]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [29]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [29]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [29]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[29]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [29]),
        .O(\badr[29]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[2]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[2]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[2]),
        .O(badr[2]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[2]_INST_0_i_10 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [2]),
        .O(\rgf/a0bus_sr [2]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [2]),
        .O(\badr[2]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[2]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [2]),
        .O(\badr[2]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [2]),
        .O(\badr[2]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[2]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [2]),
        .O(\badr[2]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [2]),
        .I5(\rgf/ivec/iv [2]),
        .O(\badr[2]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[30]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[30]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[30]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [14]),
        .O(badr[30]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[30]_INST_0_i_14 
       (.I0(\rgf/sptr/sp [30]),
        .I1(\rgf/sptr/data3 [30]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [30]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_15 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [14]),
        .O(\badr[30]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [14]),
        .O(\badr[30]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_18 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [14]),
        .O(\badr[30]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_19 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [14]),
        .O(\badr[30]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [14]),
        .O(\badr[30]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_22 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [14]),
        .O(\badr[30]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [14]),
        .O(\badr[30]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [14]),
        .O(\badr[30]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_25 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [14]),
        .O(\badr[30]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[30]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [14]),
        .O(\badr[30]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_27 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [14]),
        .O(\badr[30]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[30]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [14]),
        .O(\badr[30]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[30]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [30]),
        .O(\badr[30]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[30]_INST_0_i_8 
       (.I0(\rgf/sptr/sp [30]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [30]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [30]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[30]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [30]),
        .O(\badr[30]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA8080000A808)) 
    \badr[31]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\badr[31]_INST_0_i_4_n_0 ),
        .I5(\rgf/treg/tr [15]),
        .O(badr[31]));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_1 
       (.I0(bcmd[0]),
        .I1(\bcmd[1]_INST_0_i_1_n_0 ),
        .O(\badr[31]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[31]_INST_0_i_10 
       (.I0(\rgf/sptr/sp [31]),
        .I1(\rgf/a1bus_sel_cr [2]),
        .I2(\rgf/sptr/data3 [31]),
        .I3(\rgf/a1bus_sel_cr [5]),
        .O(\rgf/a1bus_sp [31]));
  LUT6 #(
    .INIT(64'h888888888A888888)) 
    \badr[31]_INST_0_i_100 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\badr[31]_INST_0_i_163_n_0 ),
        .I2(\badr[31]_INST_0_i_164_n_0 ),
        .I3(\fch/ir1 [2]),
        .I4(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .O(\badr[31]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_101 
       (.I0(\rgf_selc1_rn_wb[1]_i_21_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_19_n_0 ),
        .I2(fch_irq_req),
        .I3(\fch/ir1 [0]),
        .I4(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I5(\niss_dsp_a1[15]_INST_0_i_17_n_0 ),
        .O(\badr[31]_INST_0_i_101_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_102 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [11]),
        .O(\badr[31]_INST_0_i_102_n_0 ));
  LUT6 #(
    .INIT(64'h0075007F0000007F)) 
    \badr[31]_INST_0_i_103 
       (.I0(\badr[31]_INST_0_i_165_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [6]),
        .I3(\badr[31]_INST_0_i_166_n_0 ),
        .I4(\fch/ir1 [5]),
        .I5(\badr[31]_INST_0_i_167_n_0 ),
        .O(\badr[31]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'h555555555555555D)) 
    \badr[31]_INST_0_i_104 
       (.I0(\sr[15]_i_6_n_0 ),
        .I1(\badr[31]_INST_0_i_168_n_0 ),
        .I2(\badr[31]_INST_0_i_169_n_0 ),
        .I3(\badr[31]_INST_0_i_170_n_0 ),
        .I4(\badr[31]_INST_0_i_171_n_0 ),
        .I5(\badr[31]_INST_0_i_172_n_0 ),
        .O(\badr[31]_INST_0_i_104_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF005D)) 
    \badr[31]_INST_0_i_105 
       (.I0(ctl_fetch1_fl_i_16_n_0),
        .I1(\badr[31]_INST_0_i_104_n_0 ),
        .I2(\badr[31]_INST_0_i_173_n_0 ),
        .I3(\badr[31]_INST_0_i_101_n_0 ),
        .I4(\fch/ir1 [15]),
        .I5(\badr[31]_INST_0_i_174_n_0 ),
        .O(\badr[31]_INST_0_i_105_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_106 
       (.I0(\fch/ir0 [11]),
        .I1(stat[1]),
        .O(\badr[31]_INST_0_i_106_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FBFBFBAB)) 
    \badr[31]_INST_0_i_107 
       (.I0(\ccmd[0]_INST_0_i_20_n_0 ),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [14]),
        .I3(\badr[31]_INST_0_i_175_n_0 ),
        .I4(\fch/ir0 [15]),
        .I5(\badr[31]_INST_0_i_176_n_0 ),
        .O(\badr[31]_INST_0_i_107_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFD)) 
    \badr[31]_INST_0_i_108 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [13]),
        .O(\badr[31]_INST_0_i_108_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[31]_INST_0_i_109 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [7]),
        .O(\badr[31]_INST_0_i_109_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[31]_INST_0_i_11 
       (.I0(\badr[31]_INST_0_i_38_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_40_n_0 ),
        .I3(\rgf/treg/tr [31]),
        .O(\badr[31]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF9090FF)) 
    \badr[31]_INST_0_i_110 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [11]),
        .I3(stat[1]),
        .I4(\fch/ir0 [3]),
        .I5(\badr[31]_INST_0_i_177_n_0 ),
        .O(\badr[31]_INST_0_i_110_n_0 ));
  LUT6 #(
    .INIT(64'h0404040F04040404)) 
    \badr[31]_INST_0_i_111 
       (.I0(\ccmd[4]_INST_0_i_2_n_0 ),
        .I1(\badr[31]_INST_0_i_59_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_24_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\rgf_selc0_wb[1]_i_12_n_0 ),
        .O(\badr[31]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E0000000)) 
    \badr[31]_INST_0_i_112 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [9]),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(\badr[31]_INST_0_i_59_n_0 ),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [8]),
        .O(\badr[31]_INST_0_i_112_n_0 ));
  LUT6 #(
    .INIT(64'h0000080008080800)) 
    \badr[31]_INST_0_i_113 
       (.I0(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [11]),
        .O(\badr[31]_INST_0_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hFF0A00FCFFFA00FC)) 
    \badr[31]_INST_0_i_114 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [12]),
        .I5(\badr[31]_INST_0_i_178_n_0 ),
        .O(\badr[31]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h0D0D0DFF0D0D0D0D)) 
    \badr[31]_INST_0_i_115 
       (.I0(\bbus_o[5]_INST_0_i_26_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(stat[1]),
        .I3(\ccmd[3]_INST_0_i_10_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .I5(\badr[31]_INST_0_i_179_n_0 ),
        .O(\badr[31]_INST_0_i_115_n_0 ));
  LUT5 #(
    .INIT(32'h2A028AAA)) 
    \badr[31]_INST_0_i_116 
       (.I0(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .O(\badr[31]_INST_0_i_116_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[31]_INST_0_i_117 
       (.I0(\fch/ir0 [11]),
        .I1(stat[0]),
        .O(\badr[31]_INST_0_i_117_n_0 ));
  LUT6 #(
    .INIT(64'h031033D0FFFFFFFF)) 
    \badr[31]_INST_0_i_118 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [10]),
        .O(\badr[31]_INST_0_i_118_n_0 ));
  LUT5 #(
    .INIT(32'h07000000)) 
    \badr[31]_INST_0_i_119 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(crdy),
        .I4(div_crdy0),
        .O(\badr[31]_INST_0_i_119_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF00D0)) 
    \badr[31]_INST_0_i_120 
       (.I0(\badr[31]_INST_0_i_180_n_0 ),
        .I1(\badr[31]_INST_0_i_181_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(stat[0]),
        .I4(\badr[31]_INST_0_i_182_n_0 ),
        .O(\badr[31]_INST_0_i_120_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[31]_INST_0_i_121 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [15]),
        .I4(stat[1]),
        .I5(stat[2]),
        .O(\badr[31]_INST_0_i_121_n_0 ));
  LUT6 #(
    .INIT(64'h5BFBFBFBFFFFFFFF)) 
    \badr[31]_INST_0_i_122 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [2]),
        .I4(\ccmd[0]_INST_0_i_15_n_0 ),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\badr[31]_INST_0_i_122_n_0 ));
  LUT6 #(
    .INIT(64'hF8FFF8F888888888)) 
    \badr[31]_INST_0_i_123 
       (.I0(\fch/ir0 [11]),
        .I1(\badr[31]_INST_0_i_183_n_0 ),
        .I2(\bdatw[31]_INST_0_i_138_n_0 ),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [2]),
        .I5(\stat[0]_i_16__0_n_0 ),
        .O(\badr[31]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \badr[31]_INST_0_i_124 
       (.I0(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\fch_irq_lev[1]_i_6_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_24_n_0 ),
        .I4(\ccmd[3]_INST_0_i_7_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_23_n_0 ),
        .O(\badr[31]_INST_0_i_124_n_0 ));
  LUT6 #(
    .INIT(64'h00EF0B0FABEFABEF)) 
    \badr[31]_INST_0_i_125 
       (.I0(\badr[31]_INST_0_i_184_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [8]),
        .I5(\ccmd[2]_INST_0_i_4_n_0 ),
        .O(\badr[31]_INST_0_i_125_n_0 ));
  LUT5 #(
    .INIT(32'h50303030)) 
    \badr[31]_INST_0_i_126 
       (.I0(\badr[31]_INST_0_i_185_n_0 ),
        .I1(\badr[31]_INST_0_i_186_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(div_crdy0),
        .I4(crdy),
        .O(\badr[31]_INST_0_i_126_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_127 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [12]),
        .O(\badr[31]_INST_0_i_127_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA20AAAAAAAA)) 
    \badr[31]_INST_0_i_128 
       (.I0(\sr[5]_i_8_n_0 ),
        .I1(\badr[31]_INST_0_i_187_n_0 ),
        .I2(\fch/ir0 [5]),
        .I3(\badr[31]_INST_0_i_183_n_0 ),
        .I4(\badr[31]_INST_0_i_188_n_0 ),
        .I5(\badr[31]_INST_0_i_189_n_0 ),
        .O(\badr[31]_INST_0_i_128_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \badr[31]_INST_0_i_129 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(\badr[31]_INST_0_i_134_n_0 ),
        .O(\badr[31]_INST_0_i_129_n_0 ));
  LUT6 #(
    .INIT(64'h7FFF7FFFFFFF7FFF)) 
    \badr[31]_INST_0_i_130 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [10]),
        .O(\badr[31]_INST_0_i_130_n_0 ));
  LUT6 #(
    .INIT(64'h0000C40000000000)) 
    \badr[31]_INST_0_i_131 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [9]),
        .O(\badr[31]_INST_0_i_131_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \badr[31]_INST_0_i_132 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [2]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [0]),
        .I5(\fch/ir0 [3]),
        .O(\badr[31]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[31]_INST_0_i_133 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\rgf_selc0_wb[1]_i_10_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [8]),
        .O(\badr[31]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_134 
       (.I0(\ccmd[0]_INST_0_i_24_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [2]),
        .I3(fch_irq_req),
        .I4(\fch/ir0 [0]),
        .I5(\ccmd[0]_INST_0_i_22_n_0 ),
        .O(\badr[31]_INST_0_i_134_n_0 ));
  LUT5 #(
    .INIT(32'hD000FFFF)) 
    \badr[31]_INST_0_i_135 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [15]),
        .O(\badr[31]_INST_0_i_135_n_0 ));
  LUT6 #(
    .INIT(64'h0000DD0DDD0DDD0D)) 
    \badr[31]_INST_0_i_136 
       (.I0(\badr[31]_INST_0_i_190_n_0 ),
        .I1(\badr[31]_INST_0_i_191_n_0 ),
        .I2(\badr[31]_INST_0_i_192_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(\badr[31]_INST_0_i_193_n_0 ),
        .I5(\fch/ir0 [3]),
        .O(\badr[31]_INST_0_i_136_n_0 ));
  LUT6 #(
    .INIT(64'h000000F400F700F7)) 
    \badr[31]_INST_0_i_137 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [6]),
        .I2(\badr[31]_INST_0_i_184_n_0 ),
        .I3(\badr[31]_INST_0_i_194_n_0 ),
        .I4(\badr[31]_INST_0_i_195_n_0 ),
        .I5(\fch/ir0 [3]),
        .O(\badr[31]_INST_0_i_137_n_0 ));
  LUT6 #(
    .INIT(64'hAA8A8A8AAAAA8AAA)) 
    \badr[31]_INST_0_i_138 
       (.I0(\badr[31]_INST_0_i_196_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [7]),
        .I4(\badr[31]_INST_0_i_197_n_0 ),
        .I5(\badr[31]_INST_0_i_198_n_0 ),
        .O(\badr[31]_INST_0_i_138_n_0 ));
  LUT6 #(
    .INIT(64'hF2FFF2F2F2F2F2F2)) 
    \badr[31]_INST_0_i_139 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\badr[31]_INST_0_i_199_n_0 ),
        .I2(\badr[31]_INST_0_i_200_n_0 ),
        .I3(\badr[31]_INST_0_i_184_n_0 ),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [1]),
        .O(\badr[31]_INST_0_i_139_n_0 ));
  LUT6 #(
    .INIT(64'h55455555FFFFFFFF)) 
    \badr[31]_INST_0_i_140 
       (.I0(\badr[31]_INST_0_i_195_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\fch/ir0 [4]),
        .O(\badr[31]_INST_0_i_140_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \badr[31]_INST_0_i_141 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .O(\badr[31]_INST_0_i_141_n_0 ));
  LUT3 #(
    .INIT(8'h25)) 
    \badr[31]_INST_0_i_142 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [3]),
        .O(\badr[31]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'hE0FFEEFFEEFFEEFF)) 
    \badr[31]_INST_0_i_143 
       (.I0(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\stat[0]_i_20_n_0 ),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [10]),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\badr[31]_INST_0_i_143_n_0 ));
  LUT6 #(
    .INIT(64'h5410BABA5555BABA)) 
    \badr[31]_INST_0_i_144 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [6]),
        .I3(div_crdy1),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [7]),
        .O(\badr[31]_INST_0_i_144_n_0 ));
  LUT5 #(
    .INIT(32'hFF9EDFBA)) 
    \badr[31]_INST_0_i_145 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [7]),
        .O(\badr[31]_INST_0_i_145_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_146 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .O(\badr[31]_INST_0_i_146_n_0 ));
  LUT4 #(
    .INIT(16'hF4FF)) 
    \badr[31]_INST_0_i_147 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [9]),
        .O(\badr[31]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'hFE00C200CF00CF00)) 
    \badr[31]_INST_0_i_148 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [7]),
        .O(\badr[31]_INST_0_i_148_n_0 ));
  LUT5 #(
    .INIT(32'hFAFFBFBA)) 
    \badr[31]_INST_0_i_149 
       (.I0(\badr[31]_INST_0_i_201_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [7]),
        .O(\badr[31]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEF0FEFEFEFE)) 
    \badr[31]_INST_0_i_150 
       (.I0(\bcmd[1]_INST_0_i_16_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .I2(\bdatw[31]_INST_0_i_139_n_0 ),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [6]),
        .I5(\niss_dsp_a1[32]_INST_0_i_24_n_0 ),
        .O(\badr[31]_INST_0_i_150_n_0 ));
  LUT6 #(
    .INIT(64'h444444444F444444)) 
    \badr[31]_INST_0_i_151 
       (.I0(\badr[31]_INST_0_i_202_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\bdatw[31]_INST_0_i_142_n_0 ),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(\bcmd[1]_INST_0_i_16_n_0 ),
        .O(\badr[31]_INST_0_i_151_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \badr[31]_INST_0_i_152 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [15]),
        .I2(\bdatw[31]_INST_0_i_85_n_0 ),
        .O(\badr[31]_INST_0_i_152_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFEFFFEFF)) 
    \badr[31]_INST_0_i_153 
       (.I0(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I3(\niss_dsp_a1[15]_INST_0_i_18_n_0 ),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\fch/ir1 [1]),
        .O(\badr[31]_INST_0_i_153_n_0 ));
  LUT5 #(
    .INIT(32'hF03FFFE0)) 
    \badr[31]_INST_0_i_154 
       (.I0(fch_irq_req),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [3]),
        .O(\badr[31]_INST_0_i_154_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \badr[31]_INST_0_i_155 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [11]),
        .O(\badr[31]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hFF0F4F4FFFFFFFFF)) 
    \badr[31]_INST_0_i_156 
       (.I0(\fch/ir1 [14]),
        .I1(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_5_n_0 ),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [13]),
        .O(\badr[31]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F2F2FFF2F2F2)) 
    \badr[31]_INST_0_i_157 
       (.I0(\badr[31]_INST_0_i_203_n_0 ),
        .I1(\badr[31]_INST_0_i_204_n_0 ),
        .I2(\badr[15]_INST_0_i_51_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .I4(div_crdy1),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\badr[31]_INST_0_i_157_n_0 ));
  LUT4 #(
    .INIT(16'h57FF)) 
    \badr[31]_INST_0_i_158 
       (.I0(\fch/ir1 [13]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [12]),
        .O(\badr[31]_INST_0_i_158_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_159 
       (.I0(\fch/ir1 [14]),
        .I1(\rgf/sreg/sr [7]),
        .O(\badr[31]_INST_0_i_159_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \badr[31]_INST_0_i_16 
       (.I0(\rgf/sptr/sp [31]),
        .I1(\rgf/sptr/data3 [31]),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_58_n_0 ),
        .I5(\badr[31]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_sp [31]));
  LUT5 #(
    .INIT(32'hFF400000)) 
    \badr[31]_INST_0_i_160 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .O(\badr[31]_INST_0_i_160_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D2FBF2CB)) 
    \badr[31]_INST_0_i_161 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [3]),
        .I5(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .O(\badr[31]_INST_0_i_161_n_0 ));
  LUT6 #(
    .INIT(64'h33FF0030FFFFAABA)) 
    \badr[31]_INST_0_i_162 
       (.I0(\bdatw[31]_INST_0_i_85_n_0 ),
        .I1(\fch/ir1 [14]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [13]),
        .O(\badr[31]_INST_0_i_162_n_0 ));
  LUT6 #(
    .INIT(64'hAEC0AEC0AAC0AA00)) 
    \badr[31]_INST_0_i_163 
       (.I0(\badr[31]_INST_0_i_205_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [11]),
        .I4(\badr[31]_INST_0_i_206_n_0 ),
        .I5(\bcmd[1]_INST_0_i_26_n_0 ),
        .O(\badr[31]_INST_0_i_163_n_0 ));
  LUT5 #(
    .INIT(32'hFE7FFFFF)) 
    \badr[31]_INST_0_i_164 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [3]),
        .O(\badr[31]_INST_0_i_164_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[31]_INST_0_i_165 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(div_crdy1),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .O(\badr[31]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'h0010FFFF00100010)) 
    \badr[31]_INST_0_i_166 
       (.I0(\badr[31]_INST_0_i_207_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(div_crdy1),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(\badr[31]_INST_0_i_208_n_0 ),
        .I5(\fch/ir1 [10]),
        .O(\badr[31]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF707CFFFF)) 
    \badr[31]_INST_0_i_167 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [8]),
        .I3(div_crdy1),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [9]),
        .O(\badr[31]_INST_0_i_167_n_0 ));
  LUT6 #(
    .INIT(64'h7D577FD7FDFDFFFF)) 
    \badr[31]_INST_0_i_168 
       (.I0(\bdatw[31]_INST_0_i_113_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [6]),
        .O(\badr[31]_INST_0_i_168_n_0 ));
  LUT6 #(
    .INIT(64'h5500450005004500)) 
    \badr[31]_INST_0_i_169 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [8]),
        .I5(div_crdy1),
        .O(\badr[31]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \badr[31]_INST_0_i_17 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\badr[31]_INST_0_i_59_n_0 ),
        .I2(\badr[31]_INST_0_i_60_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [11]),
        .O(\badr[31]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000CCAC0000)) 
    \badr[31]_INST_0_i_170 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [10]),
        .O(\badr[31]_INST_0_i_170_n_0 ));
  LUT6 #(
    .INIT(64'h4545404054440444)) 
    \badr[31]_INST_0_i_171 
       (.I0(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [8]),
        .O(\badr[31]_INST_0_i_171_n_0 ));
  LUT6 #(
    .INIT(64'h0000A080008AA008)) 
    \badr[31]_INST_0_i_172 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [4]),
        .O(\badr[31]_INST_0_i_172_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA20AAAAAAAA)) 
    \badr[31]_INST_0_i_173 
       (.I0(\badr[31]_INST_0_i_102_n_0 ),
        .I1(\badr[31]_INST_0_i_167_n_0 ),
        .I2(\fch/ir1 [5]),
        .I3(\badr[31]_INST_0_i_209_n_0 ),
        .I4(\badr[31]_INST_0_i_210_n_0 ),
        .I5(\badr[31]_INST_0_i_211_n_0 ),
        .O(\badr[31]_INST_0_i_173_n_0 ));
  LUT6 #(
    .INIT(64'h0888888808880888)) 
    \badr[31]_INST_0_i_174 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [11]),
        .O(\badr[31]_INST_0_i_174_n_0 ));
  LUT6 #(
    .INIT(64'h88CC000088CC8000)) 
    \badr[31]_INST_0_i_175 
       (.I0(\badr[31]_INST_0_i_212_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\badr[31]_INST_0_i_175_n_0 ));
  LUT6 #(
    .INIT(64'h3303FF47FF03FF57)) 
    \badr[31]_INST_0_i_176 
       (.I0(\badr[31]_INST_0_i_213_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\badr[31]_INST_0_i_214_n_0 ),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [14]),
        .O(\badr[31]_INST_0_i_176_n_0 ));
  LUT5 #(
    .INIT(32'h44FF44F4)) 
    \badr[31]_INST_0_i_177 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [8]),
        .O(\badr[31]_INST_0_i_177_n_0 ));
  LUT6 #(
    .INIT(64'hFF02FF022222FF22)) 
    \badr[31]_INST_0_i_178 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [10]),
        .I4(\badr[31]_INST_0_i_215_n_0 ),
        .I5(\fch/ir0 [9]),
        .O(\badr[31]_INST_0_i_178_n_0 ));
  LUT5 #(
    .INIT(32'hF03FFFE0)) 
    \badr[31]_INST_0_i_179 
       (.I0(fch_irq_req),
        .I1(stat[1]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [3]),
        .O(\badr[31]_INST_0_i_179_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_18 
       (.I0(ctl_sela1),
        .I1(\badr[31]_INST_0_i_62_n_0 ),
        .O(\badr[31]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFAEBFFFFFEFFFA)) 
    \badr[31]_INST_0_i_180 
       (.I0(\ccmd[4]_INST_0_i_2_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [6]),
        .O(\badr[31]_INST_0_i_180_n_0 ));
  LUT6 #(
    .INIT(64'h00B8FFFF00FFFF3F)) 
    \badr[31]_INST_0_i_181 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [7]),
        .O(\badr[31]_INST_0_i_181_n_0 ));
  LUT6 #(
    .INIT(64'hFF10101010101010)) 
    \badr[31]_INST_0_i_182 
       (.I0(\bdatw[31]_INST_0_i_138_n_0 ),
        .I1(\badr[31]_INST_0_i_216_n_0 ),
        .I2(\badr[31]_INST_0_i_217_n_0 ),
        .I3(stat[0]),
        .I4(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\badr[31]_INST_0_i_182_n_0 ));
  LUT5 #(
    .INIT(32'h10000000)) 
    \badr[31]_INST_0_i_183 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .O(\badr[31]_INST_0_i_183_n_0 ));
  LUT5 #(
    .INIT(32'hFFBFFFFF)) 
    \badr[31]_INST_0_i_184 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(crdy),
        .I2(div_crdy0),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .O(\badr[31]_INST_0_i_184_n_0 ));
  LUT6 #(
    .INIT(64'h007C3074FF7FFF77)) 
    \badr[31]_INST_0_i_185 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [5]),
        .O(\badr[31]_INST_0_i_185_n_0 ));
  LUT6 #(
    .INIT(64'h1D1D3F1D3FFFFF0F)) 
    \badr[31]_INST_0_i_186 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [9]),
        .O(\badr[31]_INST_0_i_186_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF04C45050FFFF)) 
    \badr[31]_INST_0_i_187 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [10]),
        .O(\badr[31]_INST_0_i_187_n_0 ));
  LUT6 #(
    .INIT(64'hDD88EC4C00000000)) 
    \badr[31]_INST_0_i_188 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [8]),
        .I5(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .O(\badr[31]_INST_0_i_188_n_0 ));
  LUT6 #(
    .INIT(64'h73FBFFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_189 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\badr[31]_INST_0_i_218_n_0 ),
        .I3(\badr[31]_INST_0_i_219_n_0 ),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [10]),
        .O(\badr[31]_INST_0_i_189_n_0 ));
  LUT6 #(
    .INIT(64'h4454555544444444)) 
    \badr[31]_INST_0_i_19 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\badr[31]_INST_0_i_63_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\badr[31]_INST_0_i_64_n_0 ),
        .I4(\badr[31]_INST_0_i_65_n_0 ),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\badr[31]_INST_0_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[31]_INST_0_i_190 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [8]),
        .O(\badr[31]_INST_0_i_190_n_0 ));
  LUT6 #(
    .INIT(64'hFF33F47D3F73F53D)) 
    \badr[31]_INST_0_i_191 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [7]),
        .O(\badr[31]_INST_0_i_191_n_0 ));
  LUT6 #(
    .INIT(64'hFEF7FBF3108040C0)) 
    \badr[31]_INST_0_i_192 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [3]),
        .O(\badr[31]_INST_0_i_192_n_0 ));
  LUT6 #(
    .INIT(64'h2022222220002222)) 
    \badr[31]_INST_0_i_193 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [6]),
        .O(\badr[31]_INST_0_i_193_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF040404)) 
    \badr[31]_INST_0_i_194 
       (.I0(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(\rgf_selc0_wb[0]_i_17_n_0 ),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\badr[31]_INST_0_i_131_n_0 ),
        .O(\badr[31]_INST_0_i_194_n_0 ));
  LUT6 #(
    .INIT(64'h4440004400400044)) 
    \badr[31]_INST_0_i_195 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [6]),
        .O(\badr[31]_INST_0_i_195_n_0 ));
  LUT6 #(
    .INIT(64'h45FF45FF45FF0000)) 
    \badr[31]_INST_0_i_196 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [8]),
        .I2(\bbus_o[5]_INST_0_i_25_n_0 ),
        .I3(\bdatw[31]_INST_0_i_158_n_0 ),
        .I4(\badr[31]_INST_0_i_220_n_0 ),
        .I5(\fch/ir0 [10]),
        .O(\badr[31]_INST_0_i_196_n_0 ));
  LUT5 #(
    .INIT(32'h5FF75F7B)) 
    \badr[31]_INST_0_i_197 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [4]),
        .O(\badr[31]_INST_0_i_197_n_0 ));
  LUT5 #(
    .INIT(32'h76108010)) 
    \badr[31]_INST_0_i_198 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [3]),
        .O(\badr[31]_INST_0_i_198_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_199 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [8]),
        .O(\badr[31]_INST_0_i_199_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[31]_INST_0_i_20 
       (.I0(\badr[15]_INST_0_i_14_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .O(\badr[31]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFF00AE000000AE00)) 
    \badr[31]_INST_0_i_200 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\ccmd[0]_INST_0_i_14_n_0 ),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [4]),
        .O(\badr[31]_INST_0_i_200_n_0 ));
  LUT4 #(
    .INIT(16'hF44F)) 
    \badr[31]_INST_0_i_201 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [3]),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .O(\badr[31]_INST_0_i_201_n_0 ));
  LUT5 #(
    .INIT(32'hFBF3FBFF)) 
    \badr[31]_INST_0_i_202 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [8]),
        .O(\badr[31]_INST_0_i_202_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888808888)) 
    \badr[31]_INST_0_i_203 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .I5(div_crdy1),
        .O(\badr[31]_INST_0_i_203_n_0 ));
  LUT4 #(
    .INIT(16'h0444)) 
    \badr[31]_INST_0_i_204 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .O(\badr[31]_INST_0_i_204_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \badr[31]_INST_0_i_205 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [6]),
        .O(\badr[31]_INST_0_i_205_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_206 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [6]),
        .O(\badr[31]_INST_0_i_206_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_207 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [8]),
        .O(\badr[31]_INST_0_i_207_n_0 ));
  LUT6 #(
    .INIT(64'h5530FFFF55FFFFFF)) 
    \badr[31]_INST_0_i_208 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [2]),
        .O(\badr[31]_INST_0_i_208_n_0 ));
  LUT6 #(
    .INIT(64'hA000A08000000080)) 
    \badr[31]_INST_0_i_209 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(\fch/ir1 [5]),
        .O(\badr[31]_INST_0_i_209_n_0 ));
  LUT6 #(
    .INIT(64'h0404000404000000)) 
    \badr[31]_INST_0_i_210 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(div_crdy1),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [5]),
        .O(\badr[31]_INST_0_i_210_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF27FFFFFF)) 
    \badr[31]_INST_0_i_211 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [5]),
        .I3(\bcmd[1]_INST_0_i_15_n_0 ),
        .I4(div_crdy1),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\badr[31]_INST_0_i_211_n_0 ));
  LUT6 #(
    .INIT(64'h3F3F8F3F0F3F4F4F)) 
    \badr[31]_INST_0_i_212 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [4]),
        .O(\badr[31]_INST_0_i_212_n_0 ));
  LUT5 #(
    .INIT(32'hA20202A2)) 
    \badr[31]_INST_0_i_213 
       (.I0(\fch/ir0 [12]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir0 [14]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\rgf/sreg/sr [7]),
        .O(\badr[31]_INST_0_i_213_n_0 ));
  LUT4 #(
    .INIT(16'hB0BB)) 
    \badr[31]_INST_0_i_214 
       (.I0(\fch/ir0 [14]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [13]),
        .I3(\rgf/sreg/sr [5]),
        .O(\badr[31]_INST_0_i_214_n_0 ));
  LUT5 #(
    .INIT(32'h707C7C7C)) 
    \badr[31]_INST_0_i_215 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(crdy),
        .I4(div_crdy0),
        .O(\badr[31]_INST_0_i_215_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_216 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [9]),
        .O(\badr[31]_INST_0_i_216_n_0 ));
  LUT3 #(
    .INIT(8'h58)) 
    \badr[31]_INST_0_i_217 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .O(\badr[31]_INST_0_i_217_n_0 ));
  LUT5 #(
    .INIT(32'h3F73F53D)) 
    \badr[31]_INST_0_i_218 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [4]),
        .O(\badr[31]_INST_0_i_218_n_0 ));
  LUT5 #(
    .INIT(32'h3020308E)) 
    \badr[31]_INST_0_i_219 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [4]),
        .O(\badr[31]_INST_0_i_219_n_0 ));
  LUT6 #(
    .INIT(64'h0E0B07031F4F8FCF)) 
    \badr[31]_INST_0_i_220 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [1]),
        .O(\badr[31]_INST_0_i_220_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_23 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [15]),
        .O(\badr[31]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_24 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [15]),
        .O(\badr[31]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_30 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\badr[31]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_31 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [15]),
        .O(\badr[31]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[31]_INST_0_i_35 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_sel_cr [2]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[31]_INST_0_i_36 
       (.CI(\badr[28]_INST_0_i_21_n_0 ),
        .CO({\badr[31]_INST_0_i_36_n_2 ,\badr[31]_INST_0_i_36_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/sptr/sp [29:28]}),
        .O(\rgf/sptr/data3 [31:29]),
        .S({\<const0> ,\badr[31]_INST_0_i_70_n_0 ,\badr[31]_INST_0_i_71_n_0 ,\badr[31]_INST_0_i_72_n_0 }));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[31]_INST_0_i_37 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAF8FAFA)) 
    \badr[31]_INST_0_i_38 
       (.I0(\badr[31]_INST_0_i_73_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(stat[2]),
        .I3(\badr[31]_INST_0_i_74_n_0 ),
        .I4(\badr[31]_INST_0_i_75_n_0 ),
        .I5(ctl_sela0),
        .O(\badr[31]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h4445555544444444)) 
    \badr[31]_INST_0_i_39 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_77_n_0 ),
        .I2(\fch/ir0 [15]),
        .I3(\badr[31]_INST_0_i_78_n_0 ),
        .I4(\badr[31]_INST_0_i_79_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .O(\badr[31]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04000000)) 
    \badr[31]_INST_0_i_4 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [10]),
        .I4(\bcmd[2]_INST_0_i_3_n_0 ),
        .I5(\badr[31]_INST_0_i_17_n_0 ),
        .O(\badr[31]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[31]_INST_0_i_40 
       (.I0(\badr[31]_INST_0_i_58_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .O(\badr[31]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_43 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr25 [15]),
        .O(\badr[31]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_44 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr26 [15]),
        .O(\badr[31]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_47 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr21 [15]),
        .O(\badr[31]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_48 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank02/bank_sel00_out ),
        .I5(\rgf/bank02/gr22 [15]),
        .O(\badr[31]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[31]_INST_0_i_5 
       (.I0(\badr[31]_INST_0_i_18_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_20_n_0 ),
        .I3(\rgf/treg/tr [31]),
        .O(\badr[31]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_51 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\badr[31]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_52 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr26 [15]),
        .O(\badr[31]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_55 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr21 [15]),
        .O(\badr[31]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[31]_INST_0_i_56 
       (.I0(\badr[31]_INST_0_i_80_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\rgf/bank13/bank_sel00_out ),
        .I5(\rgf/bank13/gr22 [15]),
        .O(\badr[31]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h5554555554545454)) 
    \badr[31]_INST_0_i_57 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_82_n_0 ),
        .I2(\badr[31]_INST_0_i_83_n_0 ),
        .I3(\badr[31]_INST_0_i_84_n_0 ),
        .I4(\badr[31]_INST_0_i_85_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .O(\badr[31]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FFA2)) 
    \badr[31]_INST_0_i_58 
       (.I0(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I1(\badr[31]_INST_0_i_86_n_0 ),
        .I2(\badr[31]_INST_0_i_87_n_0 ),
        .I3(\badr[31]_INST_0_i_88_n_0 ),
        .I4(stat[2]),
        .I5(\badr[31]_INST_0_i_89_n_0 ),
        .O(\badr[31]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \badr[31]_INST_0_i_59 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [14]),
        .O(\badr[31]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[31]_INST_0_i_60 
       (.I0(stat[1]),
        .I1(stat[2]),
        .I2(stat[0]),
        .I3(\fch/ir0 [15]),
        .O(\badr[31]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBAAAAAAAA)) 
    \badr[31]_INST_0_i_61 
       (.I0(\badr[31]_INST_0_i_90_n_0 ),
        .I1(\badr[31]_INST_0_i_91_n_0 ),
        .I2(\niss_dsp_a1[15]_INST_0_i_10_n_0 ),
        .I3(\badr[31]_INST_0_i_92_n_0 ),
        .I4(\badr[31]_INST_0_i_93_n_0 ),
        .I5(\badr[31]_INST_0_i_94_n_0 ),
        .O(ctl_sela1));
  LUT6 #(
    .INIT(64'h4540454545404540)) 
    \badr[31]_INST_0_i_62 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\badr[31]_INST_0_i_95_n_0 ),
        .I2(\badr[31]_INST_0_i_96_n_0 ),
        .I3(\badr[31]_INST_0_i_97_n_0 ),
        .I4(\badr[31]_INST_0_i_98_n_0 ),
        .I5(\badr[31]_INST_0_i_99_n_0 ),
        .O(\badr[31]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAEAEAEAEAEFE)) 
    \badr[31]_INST_0_i_63 
       (.I0(\badr[31]_INST_0_i_100_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_2_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [15]),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\badr[31]_INST_0_i_63_n_0 ));
  LUT5 #(
    .INIT(32'hD000FFFF)) 
    \badr[31]_INST_0_i_64 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [15]),
        .O(\badr[31]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hBBABAAAABBBBBBBB)) 
    \badr[31]_INST_0_i_65 
       (.I0(\fch/ir1 [15]),
        .I1(\badr[31]_INST_0_i_101_n_0 ),
        .I2(\badr[31]_INST_0_i_102_n_0 ),
        .I3(\badr[31]_INST_0_i_103_n_0 ),
        .I4(\badr[31]_INST_0_i_104_n_0 ),
        .I5(ctl_fetch1_fl_i_16_n_0),
        .O(\badr[31]_INST_0_i_65_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_66 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .O(\rgf/bank02/bank_sel00_out ));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[31]_INST_0_i_67 
       (.I0(\badr[31]_INST_0_i_62_n_0 ),
        .I1(ctl_sela1),
        .O(\badr[31]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h00F2FFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_68 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\badr[31]_INST_0_i_105_n_0 ),
        .I2(\badr[31]_INST_0_i_63_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[2] ),
        .I4(ctl_sela1),
        .I5(\badr[31]_INST_0_i_62_n_0 ),
        .O(\badr[31]_INST_0_i_68_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[31]_INST_0_i_69 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .O(\rgf/bank13/bank_sel00_out ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_70 
       (.I0(\rgf/sptr/sp [30]),
        .I1(\rgf/sptr/sp [31]),
        .O(\badr[31]_INST_0_i_70_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_71 
       (.I0(\rgf/sptr/sp [29]),
        .I1(\rgf/sptr/sp [30]),
        .O(\badr[31]_INST_0_i_71_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_72 
       (.I0(\rgf/sptr/sp [28]),
        .I1(\rgf/sptr/sp [29]),
        .O(\badr[31]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFF0FFFFFDDDDDDDD)) 
    \badr[31]_INST_0_i_73 
       (.I0(\badr[31]_INST_0_i_106_n_0 ),
        .I1(\badr[31]_INST_0_i_107_n_0 ),
        .I2(\ccmd[1]_INST_0_i_5_n_0 ),
        .I3(\badr[31]_INST_0_i_108_n_0 ),
        .I4(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I5(\badr[31]_INST_0_i_74_n_0 ),
        .O(\badr[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h888888888888A8AA)) 
    \badr[31]_INST_0_i_74 
       (.I0(stat[0]),
        .I1(\badr[31]_INST_0_i_109_n_0 ),
        .I2(\badr[31]_INST_0_i_110_n_0 ),
        .I3(\badr[31]_INST_0_i_111_n_0 ),
        .I4(\badr[31]_INST_0_i_112_n_0 ),
        .I5(\badr[31]_INST_0_i_113_n_0 ),
        .O(\badr[31]_INST_0_i_74_n_0 ));
  LUT5 #(
    .INIT(32'h03770044)) 
    \badr[31]_INST_0_i_75 
       (.I0(\badr[31]_INST_0_i_114_n_0 ),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [1]),
        .I3(stat[1]),
        .I4(\badr[31]_INST_0_i_115_n_0 ),
        .O(\badr[31]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEEAEAAAAAAAA)) 
    \badr[31]_INST_0_i_76 
       (.I0(\badr[31]_INST_0_i_116_n_0 ),
        .I1(\badr[31]_INST_0_i_117_n_0 ),
        .I2(\badr[31]_INST_0_i_118_n_0 ),
        .I3(\badr[31]_INST_0_i_119_n_0 ),
        .I4(\badr[31]_INST_0_i_120_n_0 ),
        .I5(\badr[31]_INST_0_i_121_n_0 ),
        .O(ctl_sela0));
  LUT6 #(
    .INIT(64'hFFD0FFD0FFFFFFD0)) 
    \badr[31]_INST_0_i_77 
       (.I0(\badr[31]_INST_0_i_122_n_0 ),
        .I1(\badr[31]_INST_0_i_123_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I3(\badr[31]_INST_0_i_124_n_0 ),
        .I4(\ccmd[1]_INST_0_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .O(\badr[31]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555FF5D)) 
    \badr[31]_INST_0_i_78 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\badr[31]_INST_0_i_125_n_0 ),
        .I2(\badr[31]_INST_0_i_126_n_0 ),
        .I3(\badr[31]_INST_0_i_127_n_0 ),
        .I4(\badr[31]_INST_0_i_128_n_0 ),
        .I5(\badr[31]_INST_0_i_129_n_0 ),
        .O(\badr[31]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'hD555D5D5FFFFFFFF)) 
    \badr[31]_INST_0_i_79 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\badr[31]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDF0F0FFFFFFFF)) 
    \badr[31]_INST_0_i_80 
       (.I0(\badr[31]_INST_0_i_75_n_0 ),
        .I1(\badr[31]_INST_0_i_74_n_0 ),
        .I2(stat[2]),
        .I3(\fch/ir0 [11]),
        .I4(\badr[31]_INST_0_i_73_n_0 ),
        .I5(ctl_sela0),
        .O(\badr[31]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h4445555544444444)) 
    \badr[31]_INST_0_i_81 
       (.I0(stat[2]),
        .I1(\badr[31]_INST_0_i_77_n_0 ),
        .I2(\fch/ir0 [15]),
        .I3(\badr[31]_INST_0_i_78_n_0 ),
        .I4(\badr[31]_INST_0_i_79_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .O(\badr[31]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h00A2AAAA00A200A2)) 
    \badr[31]_INST_0_i_82 
       (.I0(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\ccmd[0]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_130_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\badr[31]_INST_0_i_131_n_0 ),
        .O(\badr[31]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h00000000CDC00000)) 
    \badr[31]_INST_0_i_83 
       (.I0(\rgf_selc0_rn_wb[1]_i_19_n_0 ),
        .I1(\badr[31]_INST_0_i_132_n_0 ),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\bdatw[31]_INST_0_i_24_n_0 ),
        .I5(\badr[31]_INST_0_i_133_n_0 ),
        .O(\badr[31]_INST_0_i_83_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF22F2)) 
    \badr[31]_INST_0_i_84 
       (.I0(\rgf_selc0_wb[1]_i_12_n_0 ),
        .I1(\badr[31]_INST_0_i_134_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\badr[31]_INST_0_i_135_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .O(\badr[31]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDFFFFDFFDDFF)) 
    \badr[31]_INST_0_i_85 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [12]),
        .I4(\badr[31]_INST_0_i_136_n_0 ),
        .I5(\badr[31]_INST_0_i_137_n_0 ),
        .O(\badr[31]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB3F7B3B3)) 
    \badr[31]_INST_0_i_86 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [12]),
        .I2(\badr[31]_INST_0_i_138_n_0 ),
        .I3(\badr[31]_INST_0_i_139_n_0 ),
        .I4(\badr[31]_INST_0_i_140_n_0 ),
        .I5(\badr[31]_INST_0_i_141_n_0 ),
        .O(\badr[31]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h444444444444444F)) 
    \badr[31]_INST_0_i_87 
       (.I0(\badr[31]_INST_0_i_135_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\badr[31]_INST_0_i_142_n_0 ),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [12]),
        .I5(\stat[1]_i_8__0_n_0 ),
        .O(\badr[31]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hF4FF444444444444)) 
    \badr[31]_INST_0_i_88 
       (.I0(\badr[31]_INST_0_i_143_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_7_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_23_n_0 ),
        .I4(\ccmd[1]_INST_0_i_6_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .O(\badr[31]_INST_0_i_88_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \badr[31]_INST_0_i_89 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(\fch/ir0 [15]),
        .I3(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .O(\badr[31]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h0880888808080888)) 
    \badr[31]_INST_0_i_90 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [11]),
        .O(\badr[31]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF5515FFFFFFFF)) 
    \badr[31]_INST_0_i_91 
       (.I0(\badr[31]_INST_0_i_144_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\badr[31]_INST_0_i_145_n_0 ),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\fch/ir1 [11]),
        .O(\badr[31]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h000F000F4F004400)) 
    \badr[31]_INST_0_i_92 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\badr[31]_INST_0_i_146_n_0 ),
        .I2(\badr[31]_INST_0_i_147_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [10]),
        .O(\badr[31]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h1010111011101110)) 
    \badr[31]_INST_0_i_93 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [11]),
        .I2(\badr[31]_INST_0_i_148_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [8]),
        .O(\badr[31]_INST_0_i_93_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \badr[31]_INST_0_i_94 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [15]),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\ctl1/stat_reg_n_0_[1] ),
        .O(\badr[31]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \badr[31]_INST_0_i_95 
       (.I0(\niss_dsp_a1[32]_INST_0_i_26_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [0]),
        .I5(\niss_dsp_a1[32]_INST_0_i_24_n_0 ),
        .O(\badr[31]_INST_0_i_95_n_0 ));
  LUT6 #(
    .INIT(64'h00A8AAAA00A800A8)) 
    \badr[31]_INST_0_i_96 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\badr[31]_INST_0_i_149_n_0 ),
        .I2(\badr[31]_INST_0_i_150_n_0 ),
        .I3(\badr[31]_INST_0_i_151_n_0 ),
        .I4(\bcmd[3]_INST_0_i_13_n_0 ),
        .I5(\bdatw[9]_INST_0_i_11_n_0 ),
        .O(\badr[31]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h7500FFFF75007500)) 
    \badr[31]_INST_0_i_97 
       (.I0(\badr[31]_INST_0_i_152_n_0 ),
        .I1(\badr[31]_INST_0_i_153_n_0 ),
        .I2(\badr[31]_INST_0_i_154_n_0 ),
        .I3(\badr[31]_INST_0_i_155_n_0 ),
        .I4(\badr[31]_INST_0_i_156_n_0 ),
        .I5(\badr[31]_INST_0_i_157_n_0 ),
        .O(\badr[31]_INST_0_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEEAAEA)) 
    \badr[31]_INST_0_i_98 
       (.I0(\badr[31]_INST_0_i_158_n_0 ),
        .I1(\badr[31]_INST_0_i_159_n_0 ),
        .I2(\badr[31]_INST_0_i_160_n_0 ),
        .I3(\badr[31]_INST_0_i_161_n_0 ),
        .I4(\fch/ir1 [15]),
        .I5(\badr[31]_INST_0_i_162_n_0 ),
        .O(\badr[31]_INST_0_i_98_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_99 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .O(\badr[31]_INST_0_i_99_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[3]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[3]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[3]),
        .O(badr[3]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[3]_INST_0_i_10 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [3]),
        .O(\rgf/a0bus_sr [3]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_43 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [3]),
        .O(\badr[3]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[3]_INST_0_i_44 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [3]),
        .O(\badr[3]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [3]),
        .O(\badr[3]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[3]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [3]),
        .O(\badr[3]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [3]),
        .I5(\rgf/ivec/iv [3]),
        .O(\badr[3]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[4]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[4]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[4]),
        .O(badr[4]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[4]_INST_0_i_10 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [4]),
        .O(\rgf/a0bus_sr [4]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[4]_INST_0_i_25 
       (.CI(\<const0> ),
        .CO({\badr[4]_INST_0_i_25_n_0 ,\badr[4]_INST_0_i_25_n_1 ,\badr[4]_INST_0_i_25_n_2 ,\badr[4]_INST_0_i_25_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf/sptr/sp [3],\badr[4]_INST_0_i_44_n_0 ,\badr[4]_INST_0_i_45_n_0 ,\<const0> }),
        .O(\rgf/sptr/data3 [4:1]),
        .S({\badr[4]_INST_0_i_46_n_0 ,\badr[4]_INST_0_i_47_n_0 ,\badr[4]_INST_0_i_48_n_0 ,\badr[4]_INST_0_i_49_n_0 }));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[4]_INST_0_i_44 
       (.I0(\rgf/sptr/sp [2]),
        .I1(\rgf/sptr/ctl_sp_id4 ),
        .O(\badr[4]_INST_0_i_44_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[4]_INST_0_i_45 
       (.I0(\rgf/sptr/sp [1]),
        .I1(\rgf/sptr/ctl_sp_id4 ),
        .O(\badr[4]_INST_0_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_46 
       (.I0(\rgf/sptr/sp [3]),
        .I1(\rgf/sptr/sp [4]),
        .O(\badr[4]_INST_0_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_47 
       (.I0(\rgf/sptr/sp [2]),
        .I1(\rgf/sptr/ctl_sp_id4 ),
        .I2(\rgf/sptr/sp [3]),
        .O(\badr[4]_INST_0_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_48 
       (.I0(\rgf/sptr/sp [1]),
        .I1(\rgf/sptr/ctl_sp_id4 ),
        .I2(\rgf/sptr/sp [2]),
        .O(\badr[4]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_49 
       (.I0(\rgf/sptr/sp [1]),
        .I1(\rgf/sptr/ctl_sp_id4 ),
        .O(\badr[4]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [4]),
        .O(\badr[4]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[4]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [4]),
        .O(\badr[4]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [4]),
        .O(\badr[4]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[4]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [4]),
        .O(\badr[4]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hBBAAAAAAAAAAABBB)) 
    \badr[4]_INST_0_i_54 
       (.I0(ctl_sp_id40),
        .I1(\badr[4]_INST_0_i_56_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [9]),
        .O(\rgf/sptr/ctl_sp_id4 ));
  LUT6 #(
    .INIT(64'h0000000040014005)) 
    \badr[4]_INST_0_i_55 
       (.I0(\badr[4]_INST_0_i_57_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(brdy),
        .I5(\badr[4]_INST_0_i_58_n_0 ),
        .O(ctl_sp_id40));
  LUT6 #(
    .INIT(64'hFFFFFFFF19007900)) 
    \badr[4]_INST_0_i_56 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [6]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\badr[4]_INST_0_i_59_n_0 ),
        .O(\badr[4]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAD00FD00)) 
    \badr[4]_INST_0_i_57 
       (.I0(stat[1]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [0]),
        .I3(\bcmd[3]_INST_0_i_19_n_0 ),
        .I4(brdy),
        .I5(\badr[4]_INST_0_i_60_n_0 ),
        .O(\badr[4]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hF1FFFFFFFFFFFFF0)) 
    \badr[4]_INST_0_i_58 
       (.I0(\bdatw[31]_INST_0_i_168_n_0 ),
        .I1(\badr[4]_INST_0_i_61_n_0 ),
        .I2(\badr[4]_INST_0_i_62_n_0 ),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [9]),
        .O(\badr[4]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45415551)) 
    \badr[4]_INST_0_i_59 
       (.I0(\bcmd[3]_INST_0_i_15_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [1]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\badr[4]_INST_0_i_63_n_0 ),
        .O(\badr[4]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF1)) 
    \badr[4]_INST_0_i_60 
       (.I0(\bcmd[3]_INST_0_i_19_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [15]),
        .I3(stat[0]),
        .I4(stat[2]),
        .I5(\fch/ir0 [7]),
        .O(\badr[4]_INST_0_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    \badr[4]_INST_0_i_61 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [4]),
        .I2(brdy),
        .O(\badr[4]_INST_0_i_61_n_0 ));
  LUT5 #(
    .INIT(32'hFFFE7FFE)) 
    \badr[4]_INST_0_i_62 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(stat[1]),
        .O(\badr[4]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF7F7E)) 
    \badr[4]_INST_0_i_63 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [9]),
        .I3(\bcmd[3]_INST_0_i_15_n_0 ),
        .I4(\badr[4]_INST_0_i_64_n_0 ),
        .O(\badr[4]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBC)) 
    \badr[4]_INST_0_i_64 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [7]),
        .I4(\badr[4]_INST_0_i_65_n_0 ),
        .I5(\bcmd[0]_INST_0_i_2_n_0 ),
        .O(\badr[4]_INST_0_i_64_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[4]_INST_0_i_65 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\fch/ir1 [15]),
        .O(\badr[4]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [4]),
        .I5(\rgf/ivec/iv [4]),
        .O(\badr[4]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[5]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[5]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[5]),
        .O(badr[5]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[5]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [5]),
        .O(\rgf/a0bus_sr [5]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [5]),
        .O(\badr[5]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [5]),
        .O(\badr[5]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [5]),
        .I5(\rgf/ivec/iv [5]),
        .O(\badr[5]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [5]),
        .O(\badr[5]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[5]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [5]),
        .O(\badr[5]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [5]),
        .O(\badr[5]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[5]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [5]),
        .O(\badr[5]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[5]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [5]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [5]),
        .I5(\rgf/ivec/iv [5]),
        .O(\badr[5]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[6]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[6]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[6]),
        .O(badr[6]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[6]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf/a0bus_sr [6]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [6]),
        .O(\badr[6]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [6]),
        .O(\badr[6]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [6]),
        .I5(\rgf/ivec/iv [6]),
        .O(\badr[6]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [6]),
        .O(\badr[6]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[6]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [6]),
        .O(\badr[6]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [6]),
        .O(\badr[6]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[6]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [6]),
        .O(\badr[6]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[6]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [6]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [6]),
        .I5(\rgf/ivec/iv [6]),
        .O(\badr[6]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[7]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[7]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[7]),
        .O(badr[7]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[7]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [7]),
        .O(\rgf/a0bus_sr [7]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [7]),
        .O(\badr[7]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [7]),
        .O(\badr[7]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [7]),
        .I5(\rgf/ivec/iv [7]),
        .O(\badr[7]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [7]),
        .O(\badr[7]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[7]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [7]),
        .O(\badr[7]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [7]),
        .O(\badr[7]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[7]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [7]),
        .O(\badr[7]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[7]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [7]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [7]),
        .I5(\rgf/ivec/iv [7]),
        .O(\badr[7]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[8]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[8]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[8]),
        .O(badr[8]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[8]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf/a0bus_sr [8]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [8]),
        .O(\badr[8]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [8]),
        .O(\badr[8]_INST_0_i_21_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[8]_INST_0_i_29 
       (.CI(\badr[4]_INST_0_i_25_n_0 ),
        .CO({\badr[8]_INST_0_i_29_n_0 ,\badr[8]_INST_0_i_29_n_1 ,\badr[8]_INST_0_i_29_n_2 ,\badr[8]_INST_0_i_29_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\rgf/sptr/sp [7:4]),
        .O(\rgf/sptr/data3 [8:5]),
        .S({\badr[8]_INST_0_i_46_n_0 ,\badr[8]_INST_0_i_47_n_0 ,\badr[8]_INST_0_i_48_n_0 ,\badr[8]_INST_0_i_49_n_0 }));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [8]),
        .I5(\rgf/ivec/iv [8]),
        .O(\badr[8]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_46 
       (.I0(\rgf/sptr/sp [7]),
        .I1(\rgf/sptr/sp [8]),
        .O(\badr[8]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_47 
       (.I0(\rgf/sptr/sp [6]),
        .I1(\rgf/sptr/sp [7]),
        .O(\badr[8]_INST_0_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_48 
       (.I0(\rgf/sptr/sp [5]),
        .I1(\rgf/sptr/sp [6]),
        .O(\badr[8]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_49 
       (.I0(\rgf/sptr/sp [4]),
        .I1(\rgf/sptr/sp [5]),
        .O(\badr[8]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_50 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [8]),
        .O(\badr[8]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[8]_INST_0_i_51 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [8]),
        .O(\badr[8]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_52 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [8]),
        .O(\badr[8]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[8]_INST_0_i_53 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [8]),
        .O(\badr[8]_INST_0_i_53_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[8]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [8]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [8]),
        .I5(\rgf/ivec/iv [8]),
        .O(\badr[8]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    \badr[9]_INST_0 
       (.I0(\badr[31]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[9]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(a0bus_0[9]),
        .O(badr[9]));
  LUT5 #(
    .INIT(32'h00010000)) 
    \badr[9]_INST_0_i_12 
       (.I0(\badr[31]_INST_0_i_39_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_38_n_0 ),
        .I4(\rgf/sreg/sr [9]),
        .O(\rgf/a0bus_sr [9]));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_17 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr01 [9]),
        .O(\badr[9]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [9]),
        .O(\badr[9]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_20_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[31]_INST_0_i_18_n_0 ),
        .I3(\badr[13]_INST_0_i_15_n_0 ),
        .I4(\rgf/treg/tr [9]),
        .I5(\rgf/ivec/iv [9]),
        .O(\badr[9]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_45 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [9]),
        .O(\badr[9]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0010000000000000)) 
    \badr[9]_INST_0_i_46 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr02 [9]),
        .O(\badr[9]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_47 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [9]),
        .O(\badr[9]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[9]_INST_0_i_48 
       (.I0(\badr[15]_INST_0_i_132_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [9]),
        .O(\badr[9]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[9]_INST_0_i_6 
       (.I0(\rgf/sreg/sr [9]),
        .I1(\rgf/a1bus_sel_cr [0]),
        .O(\rgf/a1bus_sr [9]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_9 
       (.I0(\badr[31]_INST_0_i_40_n_0 ),
        .I1(\badr[31]_INST_0_i_39_n_0 ),
        .I2(\badr[31]_INST_0_i_38_n_0 ),
        .I3(\badr[15]_INST_0_i_29_n_0 ),
        .I4(\rgf/treg/tr [9]),
        .I5(\rgf/ivec/iv [9]),
        .O(\badr[9]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[0]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(bbus_o[0]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bbus_o[0]_INST_0_i_1 
       (.I0(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I1(\rgf/b0bus_out/bbus_o[0]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/p_1_in3_in [0]),
        .I3(\rgf/bank02/p_0_in2_in [0]),
        .I4(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I5(p_2_in1_in[0]),
        .O(\bbus_o[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB9BB5755FFFFFFFF)) 
    \bbus_o[0]_INST_0_i_2 
       (.I0(ctl_selb0_0),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [1]),
        .I3(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_2_n_0 ),
        .O(\bbus_o[0]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[0]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_sr ));
  LUT3 #(
    .INIT(8'h08)) 
    \bbus_o[0]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [0]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[0]));
  LUT2 #(
    .INIT(4'h1)) 
    \bbus_o[0]_INST_0_i_8 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .O(\bbus_o[0]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[10]_INST_0 
       (.I0(b0bus_0[10]),
        .I1(ccmd[4]),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[11]_INST_0 
       (.I0(b0bus_0[11]),
        .I1(ccmd[4]),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[12]_INST_0 
       (.I0(b0bus_0[12]),
        .I1(ccmd[4]),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[13]_INST_0 
       (.I0(b0bus_0[13]),
        .I1(ccmd[4]),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[14]_INST_0 
       (.I0(b0bus_0[14]),
        .I1(ccmd[4]),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[15]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(ccmd[4]),
        .O(bbus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[16]_INST_0 
       (.I0(b0bus_0[16]),
        .I1(ccmd[4]),
        .O(bbus_o[16]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[17]_INST_0 
       (.I0(b0bus_0[17]),
        .I1(ccmd[4]),
        .O(bbus_o[17]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[18]_INST_0 
       (.I0(b0bus_0[18]),
        .I1(ccmd[4]),
        .O(bbus_o[18]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[19]_INST_0 
       (.I0(b0bus_0[19]),
        .I1(ccmd[4]),
        .O(bbus_o[19]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[1]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(bbus_o[1]));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bbus_o[1]_INST_0_i_1 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[1]_INST_0_i_3_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[1]_INST_0_i_4_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[1]_INST_0_i_5_n_0 ),
        .I5(p_2_in1_in[1]),
        .O(\bbus_o[1]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAA90A0AAAAA5F5F)) 
    \bbus_o[1]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [2]),
        .I4(ctl_selb0_0),
        .I5(\fch/ir0 [0]),
        .O(\bbus_o[1]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bbus_o[1]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [1]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[20]_INST_0 
       (.I0(b0bus_0[20]),
        .I1(ccmd[4]),
        .O(bbus_o[20]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[21]_INST_0 
       (.I0(b0bus_0[21]),
        .I1(ccmd[4]),
        .O(bbus_o[21]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[22]_INST_0 
       (.I0(b0bus_0[22]),
        .I1(ccmd[4]),
        .O(bbus_o[22]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[23]_INST_0 
       (.I0(b0bus_0[23]),
        .I1(ccmd[4]),
        .O(bbus_o[23]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[24]_INST_0 
       (.I0(b0bus_0[24]),
        .I1(ccmd[4]),
        .O(bbus_o[24]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[25]_INST_0 
       (.I0(b0bus_0[25]),
        .I1(ccmd[4]),
        .O(bbus_o[25]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[26]_INST_0 
       (.I0(b0bus_0[26]),
        .I1(ccmd[4]),
        .O(bbus_o[26]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[27]_INST_0 
       (.I0(b0bus_0[27]),
        .I1(ccmd[4]),
        .O(bbus_o[27]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[28]_INST_0 
       (.I0(b0bus_0[28]),
        .I1(ccmd[4]),
        .O(bbus_o[28]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[29]_INST_0 
       (.I0(b0bus_0[29]),
        .I1(ccmd[4]),
        .O(bbus_o[29]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[2]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(bbus_o[2]));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bbus_o[2]_INST_0_i_1 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[2]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[2]_INST_0_i_3_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[2]_INST_0_i_4_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[2]_INST_0_i_5_n_0 ),
        .I5(p_2_in1_in[2]),
        .O(\bbus_o[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAA900AAAAAA55FF)) 
    \bbus_o[2]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [2]),
        .I4(ctl_selb0_0),
        .I5(\fch/ir0 [1]),
        .O(\bbus_o[2]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bbus_o[2]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [2]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[30]_INST_0 
       (.I0(b0bus_0[30]),
        .I1(ccmd[4]),
        .O(bbus_o[30]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[31]_INST_0 
       (.I0(b0bus_0[31]),
        .I1(ccmd[4]),
        .O(bbus_o[31]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[3]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(bbus_o[3]));
  LUT5 #(
    .INIT(32'h00000002)) 
    \bbus_o[3]_INST_0_i_1 
       (.I0(\bbus_o[3]_INST_0_i_2_n_0 ),
        .I1(\rgf/b0bus_out/bbus_o[3]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[3]_INST_0_i_4_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[3]_INST_0_i_5_n_0 ),
        .I4(p_2_in1_in[3]),
        .O(\bbus_o[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h37F7333337F7FF3F)) 
    \bbus_o[3]_INST_0_i_2 
       (.I0(\fch/ir0 [3]),
        .I1(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I2(ctl_selb0_0),
        .I3(\bbus_o[3]_INST_0_i_7_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(\fch/ir0 [2]),
        .O(\bbus_o[3]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bbus_o[3]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [3]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[3]));
  LUT4 #(
    .INIT(16'h0040)) 
    \bbus_o[3]_INST_0_i_7 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [2]),
        .O(\bbus_o[3]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[4]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(bbus_o[4]));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bbus_o[4]_INST_0_i_1 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[4]_INST_0_i_3_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[4]_INST_0_i_4_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[4]_INST_0_i_5_n_0 ),
        .I5(p_2_in1_in[4]),
        .O(\bbus_o[4]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC3CCC44447777)) 
    \bbus_o[4]_INST_0_i_2 
       (.I0(\fch/ir0 [4]),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(\fch/ir0 [2]),
        .I3(\bdatw[12]_INST_0_i_23_n_0 ),
        .I4(\fch/ir0 [3]),
        .I5(ctl_selb0_0),
        .O(\bbus_o[4]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bbus_o[4]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [4]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[4]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(bbus_o[5]));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \bbus_o[5]_INST_0_i_1 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[5]_INST_0_i_4_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[5]_INST_0_i_5_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[5]_INST_0_i_6_n_0 ),
        .I5(p_2_in1_in[5]),
        .O(\bbus_o[5]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h5FFF5FFF5FFDF5FD)) 
    \bbus_o[5]_INST_0_i_10 
       (.I0(\fch/ir0 [13]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [12]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\fch/ir0 [14]),
        .O(\bbus_o[5]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0D05050505050505)) 
    \bbus_o[5]_INST_0_i_11 
       (.I0(\fch/ir0 [14]),
        .I1(\bbus_o[5]_INST_0_i_24_n_0 ),
        .I2(\fch/ir0 [15]),
        .I3(\bbus_o[5]_INST_0_i_25_n_0 ),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\fch/ir0 [8]),
        .O(\bbus_o[5]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hC8CCFFFFFFFFC8CC)) 
    \bbus_o[5]_INST_0_i_12 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\rgf/sreg/sr [6]),
        .I4(\bbus_o[5]_INST_0_i_26_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\bbus_o[5]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0_i_13 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .O(\bbus_o[5]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h20AA2020AAAAAAAA)) 
    \bbus_o[5]_INST_0_i_2 
       (.I0(\bbus_o[5]_INST_0_i_8_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I2(\fch/ir0 [15]),
        .I3(\bbus_o[5]_INST_0_i_10_n_0 ),
        .I4(\bbus_o[5]_INST_0_i_11_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_12_n_0 ),
        .O(\bbus_o[5]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \bbus_o[5]_INST_0_i_23 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[2]),
        .I5(ctl_selb0_rn[0]),
        .O(\rgf/b0bus_sel_cr [1]));
  LUT2 #(
    .INIT(4'h6)) 
    \bbus_o[5]_INST_0_i_24 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [5]),
        .O(\bbus_o[5]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[5]_INST_0_i_25 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .O(\bbus_o[5]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h5ACCF0FF)) 
    \bbus_o[5]_INST_0_i_26 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [12]),
        .O(\bbus_o[5]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h33CCCCCC47474747)) 
    \bbus_o[5]_INST_0_i_3 
       (.I0(\fch/ir0 [5]),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(\fch/ir0 [4]),
        .I3(\bdatw[9]_INST_0_i_17_n_0 ),
        .I4(\bbus_o[5]_INST_0_i_13_n_0 ),
        .I5(ctl_selb0_0),
        .O(\bbus_o[5]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bbus_o[5]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [5]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[5]));
  LUT3 #(
    .INIT(8'h01)) 
    \bbus_o[5]_INST_0_i_8 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(stat[2]),
        .O(\bbus_o[5]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bbus_o[5]_INST_0_i_9 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .O(\bbus_o[5]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[6]_INST_0 
       (.I0(ccmd[4]),
        .I1(\bbus_o[6]_INST_0_i_1_n_0 ),
        .O(bbus_o[6]));
  LUT6 #(
    .INIT(64'h0202020200020202)) 
    \bbus_o[6]_INST_0_i_1 
       (.I0(\bbus_o[6]_INST_0_i_2_n_0 ),
        .I1(\rgf/b0bus_out/bbus_o[6]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[6]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [6]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bbus_o[6]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \bbus_o[6]_INST_0_i_2 
       (.I0(\fch/ir0 [5]),
        .I1(ctl_selb0_0),
        .I2(\bbus_o[6]_INST_0_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(\fch/ir0 [6]),
        .I5(\bbus_o[5]_INST_0_i_2_n_0 ),
        .O(\bbus_o[6]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \bbus_o[6]_INST_0_i_5 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [2]),
        .O(\bbus_o[6]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[7]_INST_0 
       (.I0(b0bus_0[7]),
        .I1(ccmd[4]),
        .O(bbus_o[7]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bbus_o[7]_INST_0_i_1 
       (.I0(\bbus_o[7]_INST_0_i_2_n_0 ),
        .I1(\rgf/b0bus_out/bbus_o[7]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [7]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[7]));
  LUT6 #(
    .INIT(64'hAA0A08A8A00008A8)) 
    \bbus_o[7]_INST_0_i_2 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(ctl_selb0_0),
        .I3(\bbus_o[7]_INST_0_i_5_n_0 ),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(\fch/ir0 [7]),
        .O(\bbus_o[7]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bbus_o[7]_INST_0_i_5 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [2]),
        .O(\bbus_o[7]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[8]_INST_0 
       (.I0(b0bus_0[8]),
        .I1(ccmd[4]),
        .O(bbus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[9]_INST_0 
       (.I0(b0bus_0[9]),
        .I1(ccmd[4]),
        .O(bbus_o[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFF01000000)) 
    \bcmd[0]_INST_0 
       (.I0(\bcmd[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_2_n_0 ),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\bcmd[0]_INST_0_i_4_n_0 ),
        .I4(\bcmd[0]_INST_0_i_5_n_0 ),
        .I5(\bcmd[0]_INST_0_i_6_n_0 ),
        .O(bcmd[0]));
  LUT6 #(
    .INIT(64'h5501FFFFFF55FFAA)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(\fch/ir1 [11]),
        .I1(div_crdy1),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [10]),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  MUXF7 \bcmd[0]_INST_0_i_10 
       (.I0(\bcmd[0]_INST_0_i_15_n_0 ),
        .I1(\bcmd[0]_INST_0_i_16_n_0 ),
        .O(\bcmd[0]_INST_0_i_10_n_0 ),
        .S(\fch/ir0 [9]));
  LUT5 #(
    .INIT(32'hDFFFFFFD)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\bcmd[0]_INST_0_i_17_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [14]),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [8]),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \bcmd[0]_INST_0_i_13 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [5]),
        .I4(\bcmd[0]_INST_0_i_18_n_0 ),
        .O(\bcmd[0]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h9A000000)) 
    \bcmd[0]_INST_0_i_14 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [3]),
        .O(\bcmd[0]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8000000088040804)) 
    \bcmd[0]_INST_0_i_15 
       (.I0(\fch/ir0 [11]),
        .I1(\rgf_selc0_wb[1]_i_11_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [10]),
        .I4(stat[0]),
        .I5(\bcmd[0]_INST_0_i_19_n_0 ),
        .O(\bcmd[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h232300003232C030)) 
    \bcmd[0]_INST_0_i_16 
       (.I0(\bcmd[0]_INST_0_i_20_n_0 ),
        .I1(stat[0]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [11]),
        .O(\bcmd[0]_INST_0_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[0]_INST_0_i_17 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(\fch/ir0 [15]),
        .O(\bcmd[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h44D0)) 
    \bcmd[0]_INST_0_i_18 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [3]),
        .O(\bcmd[0]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \bcmd[0]_INST_0_i_19 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [4]),
        .I4(\bcmd[0]_INST_0_i_21_n_0 ),
        .O(\bcmd[0]_INST_0_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [13]),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h88000880)) 
    \bcmd[0]_INST_0_i_20 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [7]),
        .O(\bcmd[0]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h08AC)) 
    \bcmd[0]_INST_0_i_21 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(stat[0]),
        .O(\bcmd[0]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h8CBF)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(\bcmd[0]_INST_0_i_7_n_0 ),
        .I1(\mem/bctl/fch_term_fl ),
        .I2(fch_memacc1),
        .I3(\mem/bctl/ctl/p_0_in [4]),
        .O(\bcmd[0]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\fch/ir1 [15]),
        .O(\bcmd[0]_INST_0_i_4_n_0 ));
  MUXF7 \bcmd[0]_INST_0_i_5 
       (.I0(\bcmd[0]_INST_0_i_8_n_0 ),
        .I1(\bcmd[0]_INST_0_i_9_n_0 ),
        .O(\bcmd[0]_INST_0_i_5_n_0 ),
        .S(\fch/ir1 [9]));
  LUT6 #(
    .INIT(64'h2202000002000002)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(\bcmd[0]_INST_0_i_10_n_0 ),
        .I1(\bcmd[0]_INST_0_i_11_n_0 ),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .I5(\fch/ir0 [10]),
        .O(\bcmd[0]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hA8FFA8A8)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(fch_memacc1),
        .I1(\fch/fch_irq_req_fl ),
        .I2(\ir0_id_fl[21]_i_1_n_0 ),
        .I3(\mem/bctl/ctl/p_0_in [4]),
        .I4(\mem/bctl/ctl/p_0_in [5]),
        .O(\bcmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h8000000080008484)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(\fch/ir1 [11]),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [7]),
        .I5(\bcmd[0]_INST_0_i_13_n_0 ),
        .O(\bcmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0A0F00000F0AC300)) 
    \bcmd[0]_INST_0_i_9 
       (.I0(\bcmd[0]_INST_0_i_14_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [11]),
        .O(\bcmd[0]_INST_0_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \bcmd[1]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .O(bcmd[1]));
  LUT6 #(
    .INIT(64'hBBBBFFFFBBBB00F0)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(\bcmd[1]_INST_0_i_2_n_0 ),
        .I1(\bcmd[1]_INST_0_i_3_n_0 ),
        .I2(\bcmd[1]_INST_0_i_4_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\bcmd[3]_INST_0_i_4_n_0 ),
        .O(\bcmd[1]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hD5F5D5F575D5D5F5)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(\bcmd[1]_INST_0_i_22_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [7]),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(\fch/ir1 [13]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [12]),
        .O(\bcmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AAAE)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(\bcmd[1]_INST_0_i_23_n_0 ),
        .I1(\bcmd[1]_INST_0_i_24_n_0 ),
        .I2(\bcmd[1]_INST_0_i_25_n_0 ),
        .I3(\sr[6]_i_7_n_0 ),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .O(\bcmd[1]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .O(\bcmd[1]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [13]),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF7F)) 
    \bcmd[1]_INST_0_i_17 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [11]),
        .O(\bcmd[1]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBF004B00FDFFFFFF)) 
    \bcmd[1]_INST_0_i_18 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [6]),
        .O(\bcmd[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h8888888F88888888)) 
    \bcmd[1]_INST_0_i_19 
       (.I0(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I1(fch_heir_nir_i_6_n_0),
        .I2(\ccmd[1]_INST_0_i_7_n_0 ),
        .I3(\ccmd[0]_INST_0_i_24_n_0 ),
        .I4(\bcmd[1]_INST_0_i_27_n_0 ),
        .I5(\bcmd[1]_INST_0_i_28_n_0 ),
        .O(\bcmd[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF9FFF)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(\fch/ir0 [9]),
        .I1(stat[0]),
        .I2(\bcmd[1]_INST_0_i_6_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\bcmd[1]_INST_0_i_7_n_0 ),
        .I5(\bcmd[1]_INST_0_i_8_n_0 ),
        .O(\bcmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFFFFFFFFFFFFF)) 
    \bcmd[1]_INST_0_i_20 
       (.I0(\fch/ir0 [9]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\fch/ir0 [8]),
        .I4(\ccmd[2]_INST_0_i_5_n_0 ),
        .I5(\badr[31]_INST_0_i_59_n_0 ),
        .O(\bcmd[1]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \bcmd[1]_INST_0_i_21 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [4]),
        .O(\bcmd[1]_INST_0_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_22 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .O(\bcmd[1]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \bcmd[1]_INST_0_i_23 
       (.I0(\fch/ir1 [12]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(ctl_fetch1_fl_i_16_n_0),
        .I3(\bcmd[1]_INST_0_i_29_n_0 ),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [10]),
        .O(\bcmd[1]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h050000E0)) 
    \bcmd[1]_INST_0_i_24 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(fch_irq_req),
        .I2(\fch/ir1 [0]),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\fch/ir1 [3]),
        .O(\bcmd[1]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bcmd[1]_INST_0_i_25 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [14]),
        .O(\bcmd[1]_INST_0_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_26 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .O(\bcmd[1]_INST_0_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[1]_INST_0_i_27 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .O(\bcmd[1]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h050000E0)) 
    \bcmd[1]_INST_0_i_28 
       (.I0(stat[0]),
        .I1(fch_irq_req),
        .I2(\fch/ir0 [0]),
        .I3(stat[1]),
        .I4(\fch/ir0 [3]),
        .O(\bcmd[1]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_29 
       (.I0(\fch/ir1 [9]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .O(\bcmd[1]_INST_0_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(\fch/ir0 [15]),
        .I1(stat[2]),
        .O(\bcmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF44FFFFFFFFF)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(\bcmd[1]_INST_0_i_9_n_0 ),
        .I1(\bcmd[1]_INST_0_i_10_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [9]),
        .I4(\bcmd[1]_INST_0_i_11_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\bcmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAEAAAAAAAAAA)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(\bcmd[1]_INST_0_i_12_n_0 ),
        .I1(\bcmd[1]_INST_0_i_13_n_0 ),
        .I2(\bcmd[1]_INST_0_i_14_n_0 ),
        .I3(\bcmd[1]_INST_0_i_15_n_0 ),
        .I4(\bcmd[1]_INST_0_i_16_n_0 ),
        .I5(\bcmd[1]_INST_0_i_17_n_0 ),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(stat[1]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [12]),
        .O(\bcmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFAAFFFF3FFFFF)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(\bcmd[1]_INST_0_i_18_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [9]),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D0FFD0D0)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\bcmd[1]_INST_0_i_19_n_0 ),
        .I3(\bcmd[1]_INST_0_i_20_n_0 ),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\bcmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0300800000000000)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(\bcmd[1]_INST_0_i_21_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [10]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04400000)) 
    \bcmd[2]_INST_0 
       (.I0(\bcmd[2]_INST_0_i_1_n_0 ),
        .I1(\bcmd[2]_INST_0_i_2_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [10]),
        .I4(\bcmd[2]_INST_0_i_3_n_0 ),
        .I5(\bcmd[2]_INST_0_i_4_n_0 ),
        .O(bcmd[2]));
  LUT6 #(
    .INIT(64'hFDFFFFFFFFFFFFFF)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\fch/ir1 [15]),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [12]),
        .O(\bcmd[2]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .O(\bcmd[2]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h00E0)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(div_crdy1),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(\bcmd[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000220)) 
    \bcmd[2]_INST_0_i_4 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [10]),
        .I4(\ccmd[4]_INST_0_i_2_n_0 ),
        .I5(\bcmd[2]_INST_0_i_7_n_0 ),
        .O(\bcmd[2]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[2]_INST_0_i_5 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .O(\bcmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \bcmd[2]_INST_0_i_6 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [13]),
        .O(\bcmd[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    \bcmd[2]_INST_0_i_7 
       (.I0(\fch/ir0 [15]),
        .I1(stat[1]),
        .I2(stat[2]),
        .I3(\fch/ir0 [12]),
        .I4(stat[0]),
        .I5(\bcmd[2]_INST_0_i_8_n_0 ),
        .O(\bcmd[2]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bcmd[2]_INST_0_i_8 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .O(\bcmd[2]_INST_0_i_8_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \bcmd[3]_INST_0 
       (.I0(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bcmd[3]));
  LUT6 #(
    .INIT(64'h5555555155555555)) 
    \bcmd[3]_INST_0_i_1 
       (.I0(\bcmd[3]_INST_0_i_2_n_0 ),
        .I1(\bcmd[3]_INST_0_i_3_n_0 ),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\bcmd[3]_INST_0_i_4_n_0 ),
        .I4(\bcmd[3]_INST_0_i_5_n_0 ),
        .I5(\bcmd[3]_INST_0_i_6_n_0 ),
        .O(\bcmd[3]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF54550000)) 
    \bcmd[3]_INST_0_i_10 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\bcmd[3]_INST_0_i_19_n_0 ),
        .I4(\bcmd[3]_INST_0_i_20_n_0 ),
        .I5(\bcmd[3]_INST_0_i_21_n_0 ),
        .O(\bcmd[3]_INST_0_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[3]_INST_0_i_11 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [2]),
        .O(\bcmd[3]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[3]_INST_0_i_12 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [3]),
        .O(\bcmd[3]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[3]_INST_0_i_13 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [9]),
        .O(\bcmd[3]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFB7B)) 
    \bcmd[3]_INST_0_i_14 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .O(\bcmd[3]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \bcmd[3]_INST_0_i_15 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [2]),
        .O(\bcmd[3]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hBEFEFFFF)) 
    \bcmd[3]_INST_0_i_16 
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [10]),
        .O(\bcmd[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \bcmd[3]_INST_0_i_17 
       (.I0(\bcmd[3]_INST_0_i_22_n_0 ),
        .I1(\fch/ir1 [13]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\bcmd[0]_INST_0_i_12_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [10]),
        .O(\bcmd[3]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h7FFFFF5F)) 
    \bcmd[3]_INST_0_i_18 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [6]),
        .I2(\bcmd[1]_INST_0_i_6_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [8]),
        .O(\bcmd[3]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \bcmd[3]_INST_0_i_19 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [2]),
        .O(\bcmd[3]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00AE000000000000)) 
    \bcmd[3]_INST_0_i_2 
       (.I0(\bcmd[3]_INST_0_i_7_n_0 ),
        .I1(\bcmd[3]_INST_0_i_8_n_0 ),
        .I2(\bcmd[3]_INST_0_i_9_n_0 ),
        .I3(\bcmd[3]_INST_0_i_10_n_0 ),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(\bcmd[1]_INST_0_i_3_n_0 ),
        .O(\bcmd[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBFBBBBBBBBFFBBBB)) 
    \bcmd[3]_INST_0_i_20 
       (.I0(stat[0]),
        .I1(\ccmd[0]_INST_0_i_14_n_0 ),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [4]),
        .O(\bcmd[3]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00FFFFFF00004040)) 
    \bcmd[3]_INST_0_i_21 
       (.I0(\bcmd[3]_INST_0_i_23_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\bcmd[3]_INST_0_i_24_n_0 ),
        .I3(stat[0]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [7]),
        .O(\bcmd[3]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[3]_INST_0_i_22 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [14]),
        .O(\bcmd[3]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[3]_INST_0_i_23 
       (.I0(\fch/ir0 [0]),
        .I1(stat[1]),
        .O(\bcmd[3]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0101010101010001)) 
    \bcmd[3]_INST_0_i_24 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [2]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(stat[1]),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [0]),
        .O(\bcmd[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFABFA)) 
    \bcmd[3]_INST_0_i_3 
       (.I0(\bcmd[3]_INST_0_i_11_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [0]),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\bcmd[3]_INST_0_i_12_n_0 ),
        .I5(\bcmd[3]_INST_0_i_13_n_0 ),
        .O(\bcmd[3]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[3]_INST_0_i_4 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .O(\bcmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00FFFFFFFF5FFCFC)) 
    \bcmd[3]_INST_0_i_5 
       (.I0(\bcmd[3]_INST_0_i_14_n_0 ),
        .I1(\bcmd[3]_INST_0_i_15_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [7]),
        .O(\bcmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04550454)) 
    \bcmd[3]_INST_0_i_6 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(div_crdy1),
        .I5(\bcmd[3]_INST_0_i_17_n_0 ),
        .O(\bcmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FFF0F08)) 
    \bcmd[3]_INST_0_i_7 
       (.I0(crdy),
        .I1(div_crdy0),
        .I2(stat[0]),
        .I3(\fch/ir0 [11]),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(\bcmd[3]_INST_0_i_18_n_0 ),
        .O(\bcmd[3]_INST_0_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[3]_INST_0_i_8 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .O(\bcmd[3]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bcmd[3]_INST_0_i_9 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(stat[0]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [6]),
        .O(\bcmd[3]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h07)) 
    \bdatw[0]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[8]_INST_0_i_1_n_0 ),
        .O(bdatw[0]));
  LUT6 #(
    .INIT(64'h5404FFFF54045404)) 
    \bdatw[10]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(b1bus_0[10]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(b0bus_0[10]),
        .I4(\bdatw[10]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(bdatw[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAE)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(\bdatw[10]_INST_0_i_4_n_0 ),
        .I1(\bdatw[15]_INST_0_i_7_n_0 ),
        .I2(\bdatw[10]_INST_0_i_5_n_0 ),
        .I3(p_2_in4_in[10]),
        .I4(\rgf/b1bus_out/bdatw[10]_INST_0_i_7_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[10]_INST_0_i_8_n_0 ),
        .O(b1bus_0[10]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_12 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [2]),
        .O(\bdatw[10]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_13 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .O(\bdatw[10]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[10]_INST_0_i_19 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [0]),
        .O(\bdatw[10]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(\bdatw[10]_INST_0_i_9_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[10]_INST_0_i_10_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[10]_INST_0_i_11_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [10]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .O(\bdatw[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h070007000F000000)) 
    \bdatw[10]_INST_0_i_4 
       (.I0(\bdatw[10]_INST_0_i_12_n_0 ),
        .I1(\bdatw[10]_INST_0_i_13_n_0 ),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_0[2]),
        .I4(\fch/ir1 [9]),
        .I5(ctl_selb1_0[1]),
        .O(\bdatw[10]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFF7FFFF)) 
    \bdatw[10]_INST_0_i_5 
       (.I0(ctl_selb1_0[1]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [1]),
        .O(\bdatw[10]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[10]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [10]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[10]));
  LUT6 #(
    .INIT(64'hA000000008A8A8A8)) 
    \bdatw[10]_INST_0_i_9 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(ctl_selb0_0),
        .I3(\bdatw[10]_INST_0_i_19_n_0 ),
        .I4(\bdatw[11]_INST_0_i_19_n_0 ),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[10]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5404FFFF54045404)) 
    \bdatw[11]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(b1bus_0[11]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(b0bus_0[11]),
        .I4(\bdatw[11]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(bdatw[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF4)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(\bdatw[11]_INST_0_i_4_n_0 ),
        .I1(\bdatw[31]_INST_0_i_8_n_0 ),
        .I2(\bdatw[11]_INST_0_i_5_n_0 ),
        .I3(p_2_in4_in[11]),
        .I4(\rgf/b1bus_out/bdatw[11]_INST_0_i_7_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[11]_INST_0_i_8_n_0 ),
        .O(b1bus_0[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_12 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [1]),
        .O(\bdatw[11]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[11]_INST_0_i_18 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [0]),
        .O(\bdatw[11]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_19 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [2]),
        .O(\bdatw[11]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(\bdatw[11]_INST_0_i_9_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[11]_INST_0_i_10_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[11]_INST_0_i_11_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [11]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[11]_INST_0_i_3 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .O(\bdatw[11]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00008000)) 
    \bdatw[11]_INST_0_i_4 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .I2(ctl_selb1_0[1]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [2]),
        .O(\bdatw[11]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00008000AAAAAAAA)) 
    \bdatw[11]_INST_0_i_5 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(\bdatw[11]_INST_0_i_12_n_0 ),
        .I2(ctl_selb1_0[1]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [2]),
        .I5(\bdatw[31]_INST_0_i_30_n_0 ),
        .O(\bdatw[11]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[11]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [11]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[11]));
  LUT6 #(
    .INIT(64'h800080002AAA0888)) 
    \bdatw[11]_INST_0_i_9 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[11]_INST_0_i_18_n_0 ),
        .I3(\bdatw[11]_INST_0_i_19_n_0 ),
        .I4(\fch/ir0 [10]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[11]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[12]_INST_0 
       (.I0(\bdatw[12]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(b1bus_0[12]),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(b0bus_0[12]),
        .O(bdatw[12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\bdatw[12]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h55F5FF575FFFFF57)) 
    \bdatw[12]_INST_0_i_11 
       (.I0(ctl_selb1_0[2]),
        .I1(\fch/ir1 [3]),
        .I2(ctl_selb1_0[1]),
        .I3(\bdatw[12]_INST_0_i_29_n_0 ),
        .I4(\bdatw[31]_INST_0_i_12_n_0 ),
        .I5(\fch/ir1 [4]),
        .O(\bdatw[12]_INST_0_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[12]_INST_0_i_16 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [4]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[4]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(\bdatw[12]_INST_0_i_5_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[12]_INST_0_i_6_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[12]_INST_0_i_7_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [12]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_22 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [3]),
        .O(\bdatw[12]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[12]_INST_0_i_23 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [0]),
        .O(\bdatw[12]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[12]_INST_0_i_29 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [3]),
        .O(\bdatw[12]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(\bdatw[12]_INST_0_i_8_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[12]_INST_0_i_9_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[12]_INST_0_i_10_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [12]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_33 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [4]),
        .O(\bdatw[12]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \bdatw[12]_INST_0_i_34 
       (.I0(\rgf/b1bus_sel_0 [6]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/bank02/gr26 [4]),
        .O(\bdatw[12]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(\bdatw[12]_INST_0_i_11_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[12]_INST_0_i_12_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14_n_0 ),
        .I4(\rgf/b1bus_out/bdatw[12]_INST_0_i_15_n_0 ),
        .I5(p_2_in4_in[4]),
        .O(\bdatw[12]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \bdatw[12]_INST_0_i_43 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\rgf/sreg/sr [4]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sr [4]));
  LUT6 #(
    .INIT(64'h44444444444444C0)) 
    \bdatw[12]_INST_0_i_5 
       (.I0(\bdatw[31]_INST_0_i_30_n_0 ),
        .I1(ctl_selb1_0[2]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [1]),
        .I5(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[12]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_60 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr03 [4]),
        .O(\bdatw[12]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_61 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [4]),
        .O(\bdatw[12]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[12]_INST_0_i_62 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr07 [4]),
        .O(\bdatw[12]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_63 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [4]),
        .O(\bdatw[12]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_64 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr23 [4]),
        .O(\bdatw[12]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_65 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr21 [4]),
        .O(\bdatw[12]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \bdatw[12]_INST_0_i_66 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr27 [4]),
        .O(\bdatw[12]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \bdatw[12]_INST_0_i_67 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\bdatw[12]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h800080002AAA0888)) 
    \bdatw[12]_INST_0_i_8 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[12]_INST_0_i_22_n_0 ),
        .I3(\bdatw[12]_INST_0_i_23_n_0 ),
        .I4(\fch/ir0 [10]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[13]_INST_0 
       (.I0(\bdatw[13]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(b1bus_0[13]),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(b0bus_0[13]),
        .O(bdatw[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\bdatw[13]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13]_INST_0_i_4_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[13]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[13]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [13]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[13]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(\bdatw[13]_INST_0_i_7_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[13]_INST_0_i_8_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[13]_INST_0_i_9_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [13]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[13]));
  LUT6 #(
    .INIT(64'h444444444444C044)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_30_n_0 ),
        .I1(ctl_selb1_0[2]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [1]),
        .I5(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[13]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h101010101010A010)) 
    \bdatw[13]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [1]),
        .I5(\bdatw[15]_INST_0_i_22_n_0 ),
        .O(\bdatw[13]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h5404FFFF54045404)) 
    \bdatw[14]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(b1bus_0[14]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(b0bus_0[14]),
        .I4(\bdatw[14]_INST_0_i_3_n_0 ),
        .I5(\bdatw[15]_INST_0_i_4_n_0 ),
        .O(bdatw[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAC)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\bdatw[15]_INST_0_i_7_n_0 ),
        .I2(\bdatw[14]_INST_0_i_4_n_0 ),
        .I3(p_2_in4_in[14]),
        .I4(\rgf/b1bus_out/bdatw[14]_INST_0_i_6_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[14]_INST_0_i_7_n_0 ),
        .O(b1bus_0[14]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(\bdatw[14]_INST_0_i_8_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[14]_INST_0_i_9_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[14]_INST_0_i_10_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [14]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .O(\bdatw[14]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \bdatw[14]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_14_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [1]),
        .O(\bdatw[14]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[14]_INST_0_i_5 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [14]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[14]));
  LUT6 #(
    .INIT(64'h1010101010A01010)) 
    \bdatw[14]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_22_n_0 ),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [0]),
        .O(\bdatw[14]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF540454045404)) 
    \bdatw[15]_INST_0 
       (.I0(\bdatw[15]_INST_0_i_1_n_0 ),
        .I1(b1bus_0[15]),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(b0bus_0[15]),
        .I4(\bdatw[15]_INST_0_i_4_n_0 ),
        .I5(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[15]));
  LUT3 #(
    .INIT(8'hF8)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(bcmd[2]),
        .O(\bdatw[15]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h10A0101010101010)) 
    \bdatw[15]_INST_0_i_11 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I3(\bdatw[15]_INST_0_i_22_n_0 ),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [0]),
        .O(\bdatw[15]_INST_0_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \bdatw[15]_INST_0_i_14 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [2]),
        .I2(ctl_selb1_0[1]),
        .O(\bdatw[15]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .O(\rgf/b1bus_sel_cr [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFE2)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\bdatw[15]_INST_0_i_6_n_0 ),
        .I2(\bdatw[15]_INST_0_i_7_n_0 ),
        .I3(p_2_in4_in[15]),
        .I4(\rgf/b1bus_out/bdatw[15]_INST_0_i_9_n_0 ),
        .I5(\rgf/b1bus_out/bdatw[15]_INST_0_i_10_n_0 ),
        .O(b1bus_0[15]));
  LUT4 #(
    .INIT(16'h0008)) 
    \bdatw[15]_INST_0_i_21 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .O(\rgf/b1bus_sel_cr [3]));
  LUT3 #(
    .INIT(8'h7F)) 
    \bdatw[15]_INST_0_i_22 
       (.I0(ctl_selb0_0),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [2]),
        .O(\bdatw[15]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \bdatw[15]_INST_0_i_25 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[2]),
        .O(\rgf/b0bus_sel_cr [3]));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[15]_INST_0_i_29 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_cr [0]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_11_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[15]_INST_0_i_12_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[15]_INST_0_i_13_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [15]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[15]));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \bdatw[15]_INST_0_i_30 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[2]),
        .I2(ctl_selb1_rn[0]),
        .I3(ctl_selb1_0[1]),
        .I4(\bdatw[31]_INST_0_i_12_n_0 ),
        .I5(ctl_selb1_0[2]),
        .O(\rgf/b1bus_sel_cr [1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(bcmd[2]),
        .I1(\bcmd[1]_INST_0_i_1_n_0 ),
        .O(\bdatw[15]_INST_0_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[15]_INST_0_i_5 
       (.I0(b0bus_0[7]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[7]),
        .O(\bdatw[15]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[15]_INST_0_i_6 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .I2(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[15]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFAFBFAFAAAAAAAA)) 
    \bdatw[15]_INST_0_i_63 
       (.I0(\bdatw[15]_INST_0_i_90_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_48_n_0 ),
        .I2(\niss_dsp_b1[2]_INST_0_i_37_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_54_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_49_n_0 ),
        .O(\bdatw[15]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h44F5F4F5FFFFFFFF)) 
    \bdatw[15]_INST_0_i_64 
       (.I0(\bdatw[15]_INST_0_i_90_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_48_n_0 ),
        .I2(\niss_dsp_b1[2]_INST_0_i_37_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_54_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_49_n_0 ),
        .O(\bdatw[15]_INST_0_i_64_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_12_n_0 ),
        .I1(ctl_selb1_0[2]),
        .O(\bdatw[15]_INST_0_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \bdatw[15]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [15]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[15]));
  LUT6 #(
    .INIT(64'h80008080A020A0A0)) 
    \bdatw[15]_INST_0_i_90 
       (.I0(\niss_dsp_b1[5]_INST_0_i_53_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [12]),
        .I3(\bdatw[15]_INST_0_i_91_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_67_n_0 ),
        .I5(\bdatw[15]_INST_0_i_92_n_0 ),
        .O(\bdatw[15]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF44444F44)) 
    \bdatw[15]_INST_0_i_91 
       (.I0(\bdatw[15]_INST_0_i_93_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [3]),
        .I3(\bdatw[31]_INST_0_i_139_n_0 ),
        .I4(\bdatw[15]_INST_0_i_94_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_80_n_0 ),
        .O(\bdatw[15]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h88888088AAAAAAAA)) 
    \bdatw[15]_INST_0_i_92 
       (.I0(\bdatw[15]_INST_0_i_95_n_0 ),
        .I1(\badr[31]_INST_0_i_167_n_0 ),
        .I2(\bdatw[15]_INST_0_i_96_n_0 ),
        .I3(div_crdy1),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(\fch/ir1 [1]),
        .O(\bdatw[15]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hD0DCD3D3C2C2C0C0)) 
    \bdatw[15]_INST_0_i_93 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(div_crdy1),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_93_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FFFFFFFFFFFFF)) 
    \bdatw[15]_INST_0_i_94 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h7FFF7FFF777F7FFF)) 
    \bdatw[15]_INST_0_i_95 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [8]),
        .O(\bdatw[15]_INST_0_i_95_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \bdatw[15]_INST_0_i_96 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [6]),
        .O(\bdatw[15]_INST_0_i_96_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[16]_INST_0 
       (.I0(b0bus_0[16]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[16]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[16]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[16]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[16]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[16]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [16]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[16]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [0]),
        .I5(\rgf/bank02/gr25 [0]),
        .O(\bdatw[16]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [0]),
        .I5(\rgf/bank02/gr23 [0]),
        .O(\bdatw[16]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [0]),
        .I5(\rgf/bank02/gr21 [0]),
        .O(\bdatw[16]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [0]),
        .I5(\rgf/bank02/gr27 [0]),
        .O(\bdatw[16]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [0]),
        .I5(\rgf/bank02/gr25 [0]),
        .O(\bdatw[16]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [0]),
        .I5(\rgf/bank13/gr21 [0]),
        .O(\bdatw[16]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[16]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[16]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[16]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [16]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[16]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [0]),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\bdatw[16]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [0]),
        .I5(\rgf/bank13/gr21 [0]),
        .O(\bdatw[16]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [0]),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\bdatw[16]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [0]),
        .I5(\rgf/bank02/gr23 [0]),
        .O(\bdatw[16]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [0]),
        .I5(\rgf/bank02/gr21 [0]),
        .O(\bdatw[16]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [0]),
        .I5(\rgf/bank02/gr27 [0]),
        .O(\bdatw[16]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[17]_INST_0 
       (.I0(b0bus_0[17]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[17]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[17]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[17]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[17]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[17]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [17]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[17]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [1]),
        .I5(\rgf/bank02/gr25 [1]),
        .O(\bdatw[17]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [1]),
        .I5(\rgf/bank02/gr23 [1]),
        .O(\bdatw[17]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [1]),
        .I5(\rgf/bank02/gr21 [1]),
        .O(\bdatw[17]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [1]),
        .I5(\rgf/bank02/gr27 [1]),
        .O(\bdatw[17]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [1]),
        .I5(\rgf/bank02/gr25 [1]),
        .O(\bdatw[17]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [1]),
        .I5(\rgf/bank13/gr21 [1]),
        .O(\bdatw[17]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[17]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[17]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[17]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [17]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[17]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [1]),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\bdatw[17]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [1]),
        .I5(\rgf/bank13/gr21 [1]),
        .O(\bdatw[17]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [1]),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\bdatw[17]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [1]),
        .I5(\rgf/bank02/gr23 [1]),
        .O(\bdatw[17]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [1]),
        .I5(\rgf/bank02/gr21 [1]),
        .O(\bdatw[17]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [1]),
        .I5(\rgf/bank02/gr27 [1]),
        .O(\bdatw[17]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[18]_INST_0 
       (.I0(b0bus_0[18]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[18]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[18]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[18]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[18]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[18]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [18]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[18]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [2]),
        .I5(\rgf/bank02/gr25 [2]),
        .O(\bdatw[18]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [2]),
        .I5(\rgf/bank02/gr23 [2]),
        .O(\bdatw[18]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [2]),
        .I5(\rgf/bank02/gr21 [2]),
        .O(\bdatw[18]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [2]),
        .I5(\rgf/bank02/gr27 [2]),
        .O(\bdatw[18]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [2]),
        .I5(\rgf/bank02/gr25 [2]),
        .O(\bdatw[18]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [2]),
        .I5(\rgf/bank13/gr21 [2]),
        .O(\bdatw[18]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[18]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[18]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[18]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [18]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[18]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [2]),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\bdatw[18]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [2]),
        .I5(\rgf/bank13/gr21 [2]),
        .O(\bdatw[18]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [2]),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\bdatw[18]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [2]),
        .I5(\rgf/bank02/gr23 [2]),
        .O(\bdatw[18]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [2]),
        .I5(\rgf/bank02/gr21 [2]),
        .O(\bdatw[18]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [2]),
        .I5(\rgf/bank02/gr27 [2]),
        .O(\bdatw[18]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[19]_INST_0 
       (.I0(b0bus_0[19]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[19]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[19]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[19]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[19]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[19]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [19]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[19]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [3]),
        .I5(\rgf/bank02/gr25 [3]),
        .O(\bdatw[19]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [3]),
        .I5(\rgf/bank02/gr23 [3]),
        .O(\bdatw[19]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [3]),
        .I5(\rgf/bank02/gr21 [3]),
        .O(\bdatw[19]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [3]),
        .I5(\rgf/bank02/gr27 [3]),
        .O(\bdatw[19]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [3]),
        .I5(\rgf/bank02/gr25 [3]),
        .O(\bdatw[19]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [3]),
        .I5(\rgf/bank13/gr21 [3]),
        .O(\bdatw[19]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[19]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[19]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[19]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [19]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[19]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [3]),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\bdatw[19]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [3]),
        .I5(\rgf/bank13/gr21 [3]),
        .O(\bdatw[19]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [3]),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\bdatw[19]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [3]),
        .I5(\rgf/bank02/gr23 [3]),
        .O(\bdatw[19]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [3]),
        .I5(\rgf/bank02/gr21 [3]),
        .O(\bdatw[19]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [3]),
        .I5(\rgf/bank02/gr27 [3]),
        .O(\bdatw[19]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h07)) 
    \bdatw[1]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[9]_INST_0_i_1_n_0 ),
        .O(bdatw[1]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[20]_INST_0 
       (.I0(b0bus_0[20]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[20]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[20]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[20]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[20]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[20]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [20]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[20]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [4]),
        .I5(\rgf/bank02/gr25 [4]),
        .O(\bdatw[20]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [4]),
        .I5(\rgf/bank02/gr23 [4]),
        .O(\bdatw[20]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [4]),
        .I5(\rgf/bank02/gr21 [4]),
        .O(\bdatw[20]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [4]),
        .I5(\rgf/bank02/gr27 [4]),
        .O(\bdatw[20]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [4]),
        .I5(\rgf/bank02/gr25 [4]),
        .O(\bdatw[20]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [4]),
        .I5(\rgf/bank13/gr21 [4]),
        .O(\bdatw[20]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[20]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[20]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[20]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [20]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[20]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [4]),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\bdatw[20]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [4]),
        .I5(\rgf/bank13/gr21 [4]),
        .O(\bdatw[20]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [4]),
        .I5(\rgf/bank13/gr25 [4]),
        .O(\bdatw[20]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [4]),
        .I5(\rgf/bank02/gr23 [4]),
        .O(\bdatw[20]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [4]),
        .I5(\rgf/bank02/gr21 [4]),
        .O(\bdatw[20]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [4]),
        .I5(\rgf/bank02/gr27 [4]),
        .O(\bdatw[20]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[21]_INST_0 
       (.I0(b0bus_0[21]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[21]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[21]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[21]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[21]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[21]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [21]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[21]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [5]),
        .I5(\rgf/bank02/gr25 [5]),
        .O(\bdatw[21]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [5]),
        .I5(\rgf/bank02/gr23 [5]),
        .O(\bdatw[21]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [5]),
        .I5(\rgf/bank02/gr21 [5]),
        .O(\bdatw[21]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [5]),
        .I5(\rgf/bank02/gr27 [5]),
        .O(\bdatw[21]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [5]),
        .I5(\rgf/bank02/gr25 [5]),
        .O(\bdatw[21]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [5]),
        .I5(\rgf/bank13/gr21 [5]),
        .O(\bdatw[21]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[21]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[21]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[21]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [21]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[21]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [5]),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\bdatw[21]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [5]),
        .I5(\rgf/bank13/gr21 [5]),
        .O(\bdatw[21]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [5]),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\bdatw[21]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [5]),
        .I5(\rgf/bank02/gr23 [5]),
        .O(\bdatw[21]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [5]),
        .I5(\rgf/bank02/gr21 [5]),
        .O(\bdatw[21]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [5]),
        .I5(\rgf/bank02/gr27 [5]),
        .O(\bdatw[21]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[22]_INST_0 
       (.I0(b0bus_0[22]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[22]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[22]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[22]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[22]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[22]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [22]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[22]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [6]),
        .I5(\rgf/bank02/gr25 [6]),
        .O(\bdatw[22]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [6]),
        .I5(\rgf/bank02/gr23 [6]),
        .O(\bdatw[22]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [6]),
        .I5(\rgf/bank02/gr21 [6]),
        .O(\bdatw[22]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [6]),
        .I5(\rgf/bank02/gr27 [6]),
        .O(\bdatw[22]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [6]),
        .I5(\rgf/bank02/gr25 [6]),
        .O(\bdatw[22]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [6]),
        .I5(\rgf/bank13/gr21 [6]),
        .O(\bdatw[22]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[22]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[22]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[22]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [22]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[22]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [6]),
        .I5(\rgf/bank13/gr25 [6]),
        .O(\bdatw[22]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [6]),
        .I5(\rgf/bank13/gr21 [6]),
        .O(\bdatw[22]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [6]),
        .I5(\rgf/bank13/gr25 [6]),
        .O(\bdatw[22]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [6]),
        .I5(\rgf/bank02/gr23 [6]),
        .O(\bdatw[22]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [6]),
        .I5(\rgf/bank02/gr21 [6]),
        .O(\bdatw[22]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [6]),
        .I5(\rgf/bank02/gr27 [6]),
        .O(\bdatw[22]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[23]_INST_0 
       (.I0(b0bus_0[23]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[23]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[23]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[23]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[23]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[23]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [23]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[23]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [7]),
        .I5(\rgf/bank02/gr25 [7]),
        .O(\bdatw[23]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [7]),
        .I5(\rgf/bank02/gr23 [7]),
        .O(\bdatw[23]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [7]),
        .I5(\rgf/bank02/gr21 [7]),
        .O(\bdatw[23]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [7]),
        .I5(\rgf/bank02/gr27 [7]),
        .O(\bdatw[23]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [7]),
        .I5(\rgf/bank02/gr25 [7]),
        .O(\bdatw[23]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [7]),
        .I5(\rgf/bank13/gr21 [7]),
        .O(\bdatw[23]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[23]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[23]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[23]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [23]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[23]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [7]),
        .I5(\rgf/bank13/gr25 [7]),
        .O(\bdatw[23]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [7]),
        .I5(\rgf/bank13/gr21 [7]),
        .O(\bdatw[23]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [7]),
        .I5(\rgf/bank13/gr25 [7]),
        .O(\bdatw[23]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [7]),
        .I5(\rgf/bank02/gr23 [7]),
        .O(\bdatw[23]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [7]),
        .I5(\rgf/bank02/gr21 [7]),
        .O(\bdatw[23]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [7]),
        .I5(\rgf/bank02/gr27 [7]),
        .O(\bdatw[23]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[24]_INST_0 
       (.I0(b0bus_0[24]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[24]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[24]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[24]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[24]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[24]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [24]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[24]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [8]),
        .I5(\rgf/bank02/gr25 [8]),
        .O(\bdatw[24]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [8]),
        .I5(\rgf/bank02/gr23 [8]),
        .O(\bdatw[24]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [8]),
        .I5(\rgf/bank02/gr21 [8]),
        .O(\bdatw[24]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [8]),
        .I5(\rgf/bank02/gr27 [8]),
        .O(\bdatw[24]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [8]),
        .I5(\rgf/bank02/gr25 [8]),
        .O(\bdatw[24]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [8]),
        .I5(\rgf/bank13/gr21 [8]),
        .O(\bdatw[24]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[24]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[24]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[24]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [24]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[24]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [8]),
        .I5(\rgf/bank13/gr25 [8]),
        .O(\bdatw[24]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [8]),
        .I5(\rgf/bank13/gr21 [8]),
        .O(\bdatw[24]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [8]),
        .I5(\rgf/bank13/gr25 [8]),
        .O(\bdatw[24]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [8]),
        .I5(\rgf/bank02/gr23 [8]),
        .O(\bdatw[24]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [8]),
        .I5(\rgf/bank02/gr21 [8]),
        .O(\bdatw[24]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [8]),
        .I5(\rgf/bank02/gr27 [8]),
        .O(\bdatw[24]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[25]_INST_0 
       (.I0(b0bus_0[25]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[25]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[25]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[25]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[25]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[25]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [25]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[25]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [9]),
        .I5(\rgf/bank02/gr25 [9]),
        .O(\bdatw[25]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [9]),
        .I5(\rgf/bank02/gr23 [9]),
        .O(\bdatw[25]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [9]),
        .I5(\rgf/bank02/gr21 [9]),
        .O(\bdatw[25]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [9]),
        .I5(\rgf/bank02/gr27 [9]),
        .O(\bdatw[25]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [9]),
        .I5(\rgf/bank02/gr25 [9]),
        .O(\bdatw[25]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [9]),
        .I5(\rgf/bank13/gr21 [9]),
        .O(\bdatw[25]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[25]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[25]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[25]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [25]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[25]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [9]),
        .I5(\rgf/bank13/gr25 [9]),
        .O(\bdatw[25]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [9]),
        .I5(\rgf/bank13/gr21 [9]),
        .O(\bdatw[25]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [9]),
        .I5(\rgf/bank13/gr25 [9]),
        .O(\bdatw[25]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [9]),
        .I5(\rgf/bank02/gr23 [9]),
        .O(\bdatw[25]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [9]),
        .I5(\rgf/bank02/gr21 [9]),
        .O(\bdatw[25]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [9]),
        .I5(\rgf/bank02/gr27 [9]),
        .O(\bdatw[25]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[26]_INST_0 
       (.I0(b0bus_0[26]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[26]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[26]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[26]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[26]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[26]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [26]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[26]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [10]),
        .I5(\rgf/bank02/gr25 [10]),
        .O(\bdatw[26]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [10]),
        .I5(\rgf/bank02/gr23 [10]),
        .O(\bdatw[26]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [10]),
        .I5(\rgf/bank02/gr21 [10]),
        .O(\bdatw[26]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [10]),
        .I5(\rgf/bank02/gr27 [10]),
        .O(\bdatw[26]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [10]),
        .I5(\rgf/bank02/gr25 [10]),
        .O(\bdatw[26]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [10]),
        .I5(\rgf/bank13/gr21 [10]),
        .O(\bdatw[26]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[26]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[26]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[26]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [26]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[26]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [10]),
        .I5(\rgf/bank13/gr25 [10]),
        .O(\bdatw[26]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [10]),
        .I5(\rgf/bank13/gr21 [10]),
        .O(\bdatw[26]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [10]),
        .I5(\rgf/bank13/gr25 [10]),
        .O(\bdatw[26]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [10]),
        .I5(\rgf/bank02/gr23 [10]),
        .O(\bdatw[26]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [10]),
        .I5(\rgf/bank02/gr21 [10]),
        .O(\bdatw[26]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [10]),
        .I5(\rgf/bank02/gr27 [10]),
        .O(\bdatw[26]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[27]_INST_0 
       (.I0(b0bus_0[27]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[27]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[27]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[27]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[27]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[27]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [27]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[27]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [11]),
        .I5(\rgf/bank02/gr25 [11]),
        .O(\bdatw[27]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [11]),
        .I5(\rgf/bank02/gr23 [11]),
        .O(\bdatw[27]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [11]),
        .I5(\rgf/bank02/gr21 [11]),
        .O(\bdatw[27]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [11]),
        .I5(\rgf/bank02/gr27 [11]),
        .O(\bdatw[27]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [11]),
        .I5(\rgf/bank02/gr25 [11]),
        .O(\bdatw[27]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [11]),
        .I5(\rgf/bank13/gr21 [11]),
        .O(\bdatw[27]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[27]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[27]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[27]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [27]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[27]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [11]),
        .I5(\rgf/bank13/gr25 [11]),
        .O(\bdatw[27]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [11]),
        .I5(\rgf/bank13/gr21 [11]),
        .O(\bdatw[27]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [11]),
        .I5(\rgf/bank13/gr25 [11]),
        .O(\bdatw[27]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [11]),
        .I5(\rgf/bank02/gr23 [11]),
        .O(\bdatw[27]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [11]),
        .I5(\rgf/bank02/gr21 [11]),
        .O(\bdatw[27]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [11]),
        .I5(\rgf/bank02/gr27 [11]),
        .O(\bdatw[27]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[28]_INST_0 
       (.I0(b0bus_0[28]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[28]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[28]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[28]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[28]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[28]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [28]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[28]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [12]),
        .I5(\rgf/bank02/gr25 [12]),
        .O(\bdatw[28]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [12]),
        .I5(\rgf/bank02/gr23 [12]),
        .O(\bdatw[28]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [12]),
        .I5(\rgf/bank02/gr21 [12]),
        .O(\bdatw[28]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [12]),
        .I5(\rgf/bank02/gr27 [12]),
        .O(\bdatw[28]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [12]),
        .I5(\rgf/bank02/gr25 [12]),
        .O(\bdatw[28]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [12]),
        .I5(\rgf/bank13/gr21 [12]),
        .O(\bdatw[28]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[28]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[28]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[28]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [28]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[28]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [12]),
        .I5(\rgf/bank13/gr25 [12]),
        .O(\bdatw[28]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [12]),
        .I5(\rgf/bank13/gr21 [12]),
        .O(\bdatw[28]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [12]),
        .I5(\rgf/bank13/gr25 [12]),
        .O(\bdatw[28]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [12]),
        .I5(\rgf/bank02/gr23 [12]),
        .O(\bdatw[28]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [12]),
        .I5(\rgf/bank02/gr21 [12]),
        .O(\bdatw[28]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [12]),
        .I5(\rgf/bank02/gr27 [12]),
        .O(\bdatw[28]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[29]_INST_0 
       (.I0(b0bus_0[29]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[29]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[29]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[29]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[29]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[29]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [29]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[29]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [13]),
        .I5(\rgf/bank02/gr25 [13]),
        .O(\bdatw[29]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [13]),
        .I5(\rgf/bank02/gr23 [13]),
        .O(\bdatw[29]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [13]),
        .I5(\rgf/bank02/gr21 [13]),
        .O(\bdatw[29]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [13]),
        .I5(\rgf/bank02/gr27 [13]),
        .O(\bdatw[29]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [13]),
        .I5(\rgf/bank02/gr25 [13]),
        .O(\bdatw[29]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [13]),
        .I5(\rgf/bank13/gr21 [13]),
        .O(\bdatw[29]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[29]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[29]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[29]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [29]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[29]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [13]),
        .I5(\rgf/bank13/gr25 [13]),
        .O(\bdatw[29]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [13]),
        .I5(\rgf/bank13/gr21 [13]),
        .O(\bdatw[29]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [13]),
        .I5(\rgf/bank13/gr25 [13]),
        .O(\bdatw[29]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [13]),
        .I5(\rgf/bank02/gr23 [13]),
        .O(\bdatw[29]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [13]),
        .I5(\rgf/bank02/gr21 [13]),
        .O(\bdatw[29]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [13]),
        .I5(\rgf/bank02/gr27 [13]),
        .O(\bdatw[29]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h07)) 
    \bdatw[2]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[10]_INST_0_i_3_n_0 ),
        .O(bdatw[2]));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[30]_INST_0 
       (.I0(b0bus_0[30]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[30]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[30]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[30]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[30]_INST_0_i_3_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[30]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [30]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[30]));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [14]),
        .I5(\rgf/bank02/gr25 [14]),
        .O(\bdatw[30]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [14]),
        .I5(\rgf/bank02/gr23 [14]),
        .O(\bdatw[30]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [14]),
        .I5(\rgf/bank02/gr21 [14]),
        .O(\bdatw[30]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [14]),
        .I5(\rgf/bank02/gr27 [14]),
        .O(\bdatw[30]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [14]),
        .I5(\rgf/bank02/gr25 [14]),
        .O(\bdatw[30]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_19 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [14]),
        .I5(\rgf/bank13/gr21 [14]),
        .O(\bdatw[30]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[30]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[30]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[30]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [30]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[30]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [14]),
        .I5(\rgf/bank13/gr25 [14]),
        .O(\bdatw[30]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [14]),
        .I5(\rgf/bank13/gr21 [14]),
        .O(\bdatw[30]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_22 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [14]),
        .I5(\rgf/bank13/gr25 [14]),
        .O(\bdatw[30]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [14]),
        .I5(\rgf/bank02/gr23 [14]),
        .O(\bdatw[30]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_8 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [14]),
        .I5(\rgf/bank02/gr21 [14]),
        .O(\bdatw[30]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [14]),
        .I5(\rgf/bank02/gr27 [14]),
        .O(\bdatw[30]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \bdatw[31]_INST_0 
       (.I0(b0bus_0[31]),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(b1bus_0[31]),
        .I3(\bcmd[3]_INST_0_i_1_n_0 ),
        .O(bdatw[31]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[31]_INST_0_i_1 
       (.I0(\bdatw[31]_INST_0_i_3_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[31]_INST_0_i_4_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[31]_INST_0_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [31]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[31]));
  LUT6 #(
    .INIT(64'hFFFFDFFFDDDDDDDD)) 
    \bdatw[31]_INST_0_i_100 
       (.I0(\fch/ir1 [13]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\bdatw[31]_INST_0_i_141_n_0 ),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(\bdatw[31]_INST_0_i_142_n_0 ),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\bdatw[31]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFFFDDCFCFCCCC)) 
    \bdatw[31]_INST_0_i_101 
       (.I0(\bdatw[31]_INST_0_i_143_n_0 ),
        .I1(\bdatw[31]_INST_0_i_144_n_0 ),
        .I2(\bdatw[31]_INST_0_i_145_n_0 ),
        .I3(\bdatw[31]_INST_0_i_146_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\bdatw[31]_INST_0_i_147_n_0 ),
        .O(\bdatw[31]_INST_0_i_101_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \bdatw[31]_INST_0_i_102 
       (.I0(\bcmd[1]_INST_0_i_24_n_0 ),
        .I1(\bdatw[31]_INST_0_i_148_n_0 ),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [11]),
        .O(\bdatw[31]_INST_0_i_102_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_103 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [2]),
        .O(\bdatw[31]_INST_0_i_103_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_104 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [14]),
        .O(\bdatw[31]_INST_0_i_104_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1400)) 
    \bdatw[31]_INST_0_i_105 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [6]),
        .I3(\bdatw[31]_INST_0_i_149_n_0 ),
        .I4(\bdatw[31]_INST_0_i_150_n_0 ),
        .O(\bdatw[31]_INST_0_i_105_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7FDFF77)) 
    \bdatw[31]_INST_0_i_106 
       (.I0(\bdatw[31]_INST_0_i_151_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [4]),
        .I5(\bdatw[31]_INST_0_i_152_n_0 ),
        .O(\bdatw[31]_INST_0_i_106_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_107 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [8]),
        .O(\bdatw[31]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8AFA8A8)) 
    \bdatw[31]_INST_0_i_108 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(div_crdy1),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\bdatw[31]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hAAEAFFAEAAFAFFBF)) 
    \bdatw[31]_INST_0_i_109 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [6]),
        .I5(div_crdy1),
        .O(\bdatw[31]_INST_0_i_109_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_11 
       (.I0(ctl_selb1_0[1]),
        .I1(ctl_selb1_0[2]),
        .O(\bdatw[31]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h15404015)) 
    \bdatw[31]_INST_0_i_110 
       (.I0(\fch/ir1 [13]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\fch/ir1 [11]),
        .O(\bdatw[31]_INST_0_i_110_n_0 ));
  LUT6 #(
    .INIT(64'h0000400040000000)) 
    \bdatw[31]_INST_0_i_111 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [9]),
        .O(\bdatw[31]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFDFFFFFF)) 
    \bdatw[31]_INST_0_i_112 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [3]),
        .I3(\bdatw[31]_INST_0_i_153_n_0 ),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [4]),
        .O(\bdatw[31]_INST_0_i_112_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \bdatw[31]_INST_0_i_113 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [10]),
        .O(\bdatw[31]_INST_0_i_113_n_0 ));
  LUT5 #(
    .INIT(32'h8A80202A)) 
    \bdatw[31]_INST_0_i_114 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [13]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir1 [11]),
        .O(\bdatw[31]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FFFEFFFE)) 
    \bdatw[31]_INST_0_i_115 
       (.I0(\bdatw[31]_INST_0_i_154_n_0 ),
        .I1(\bdatw[31]_INST_0_i_155_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_19_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch_irq_lev[1]_i_7_n_0 ),
        .I5(\fch/ir1 [13]),
        .O(\bdatw[31]_INST_0_i_115_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_116 
       (.I0(\fch/ir1 [13]),
        .I1(\rgf/sreg/sr [6]),
        .O(\bdatw[31]_INST_0_i_116_n_0 ));
  LUT6 #(
    .INIT(64'h000F2F2F0F2F2F2F)) 
    \bdatw[31]_INST_0_i_117 
       (.I0(\bdatw[31]_INST_0_i_156_n_0 ),
        .I1(\badr[31]_INST_0_i_195_n_0 ),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [6]),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\bdatw[31]_INST_0_i_138_n_0 ),
        .O(\bdatw[31]_INST_0_i_117_n_0 ));
  LUT5 #(
    .INIT(32'h00002A22)) 
    \bdatw[31]_INST_0_i_118 
       (.I0(\bdatw[31]_INST_0_i_157_n_0 ),
        .I1(\fch/ir0 [1]),
        .I2(\bdatw[31]_INST_0_i_158_n_0 ),
        .I3(\bdatw[31]_INST_0_i_159_n_0 ),
        .I4(\bdatw[31]_INST_0_i_160_n_0 ),
        .O(\bdatw[31]_INST_0_i_118_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \bdatw[31]_INST_0_i_119 
       (.I0(stat[0]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .I3(stat[2]),
        .I4(stat[1]),
        .I5(\fch/ir0 [15]),
        .O(\bdatw[31]_INST_0_i_119_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF0DFF0DFF0D)) 
    \bdatw[31]_INST_0_i_12 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\bdatw[31]_INST_0_i_41_n_0 ),
        .I2(\bdatw[31]_INST_0_i_42_n_0 ),
        .I3(\bdatw[31]_INST_0_i_43_n_0 ),
        .I4(\bdatw[31]_INST_0_i_44_n_0 ),
        .I5(\bdatw[31]_INST_0_i_45_n_0 ),
        .O(\bdatw[31]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000048000000)) 
    \bdatw[31]_INST_0_i_120 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [1]),
        .I4(\badr[31]_INST_0_i_121_n_0 ),
        .I5(\bdatw[31]_INST_0_i_161_n_0 ),
        .O(\bdatw[31]_INST_0_i_120_n_0 ));
  LUT6 #(
    .INIT(64'hD0DDDDDDFFFFFFFF)) 
    \bdatw[31]_INST_0_i_121 
       (.I0(\fch/ir0 [0]),
        .I1(\bdatw[31]_INST_0_i_162_n_0 ),
        .I2(\bdatw[31]_INST_0_i_163_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\sr[5]_i_8_n_0 ),
        .O(\bdatw[31]_INST_0_i_121_n_0 ));
  LUT5 #(
    .INIT(32'h00A20000)) 
    \bdatw[31]_INST_0_i_122 
       (.I0(\fch/ir0 [0]),
        .I1(\bdatw[31]_INST_0_i_156_n_0 ),
        .I2(\bdatw[31]_INST_0_i_164_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .O(\bdatw[31]_INST_0_i_122_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \bdatw[31]_INST_0_i_123 
       (.I0(\bdatw[31]_INST_0_i_165_n_0 ),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [7]),
        .I4(stat[2]),
        .I5(stat[1]),
        .O(\bdatw[31]_INST_0_i_123_n_0 ));
  LUT6 #(
    .INIT(64'hD500FFFFFFFFFFFF)) 
    \bdatw[31]_INST_0_i_124 
       (.I0(\fch/ir0 [2]),
        .I1(\bdatw[31]_INST_0_i_159_n_0 ),
        .I2(\bdatw[31]_INST_0_i_166_n_0 ),
        .I3(\bdatw[31]_INST_0_i_167_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [12]),
        .O(\bdatw[31]_INST_0_i_124_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDFDDDF)) 
    \bdatw[31]_INST_0_i_125 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [11]),
        .I2(\bdatw[31]_INST_0_i_164_n_0 ),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(ctl_fetch0_fl_i_28_n_0),
        .I5(\bdatw[31]_INST_0_i_128_n_0 ),
        .O(\bdatw[31]_INST_0_i_125_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFFFFFFF)) 
    \bdatw[31]_INST_0_i_126 
       (.I0(\bdatw[31]_INST_0_i_165_n_0 ),
        .I1(stat[1]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [6]),
        .I5(\badr[31]_INST_0_i_124_n_0 ),
        .O(\bdatw[31]_INST_0_i_126_n_0 ));
  LUT4 #(
    .INIT(16'hA415)) 
    \bdatw[31]_INST_0_i_127 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\bdatw[31]_INST_0_i_127_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_128 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [9]),
        .O(\bdatw[31]_INST_0_i_128_n_0 ));
  LUT6 #(
    .INIT(64'h1505050510101010)) 
    \bdatw[31]_INST_0_i_129 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(crdy),
        .I4(div_crdy0),
        .I5(\fch/ir0 [10]),
        .O(\bdatw[31]_INST_0_i_129_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_13 
       (.I0(ctl_selb0_0),
        .I1(\fch/ir0 [10]),
        .O(\bdatw[31]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0C3C8C3F003C003F)) 
    \bdatw[31]_INST_0_i_130 
       (.I0(\bdatw[31]_INST_0_i_168_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [6]),
        .O(\bdatw[31]_INST_0_i_130_n_0 ));
  LUT5 #(
    .INIT(32'h8C004004)) 
    \bdatw[31]_INST_0_i_131 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [3]),
        .O(\bdatw[31]_INST_0_i_131_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_132 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .O(\bdatw[31]_INST_0_i_132_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[31]_INST_0_i_133 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .O(\bdatw[31]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'h00000F0F00000222)) 
    \bdatw[31]_INST_0_i_134 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [6]),
        .I4(ctl_fetch0_fl_i_29_n_0),
        .I5(\fch/ir0 [10]),
        .O(\bdatw[31]_INST_0_i_134_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[31]_INST_0_i_135 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [12]),
        .O(\bdatw[31]_INST_0_i_135_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[31]_INST_0_i_136 
       (.I0(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\ccmd[1]_INST_0_i_13_n_0 ),
        .I3(\fch/ir0 [1]),
        .I4(\fch/ir0 [6]),
        .I5(\bdatw[31]_INST_0_i_135_n_0 ),
        .O(\bdatw[31]_INST_0_i_136_n_0 ));
  LUT6 #(
    .INIT(64'h0131D80003332000)) 
    \bdatw[31]_INST_0_i_137 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [6]),
        .O(\bdatw[31]_INST_0_i_137_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_138 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .O(\bdatw[31]_INST_0_i_138_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[31]_INST_0_i_139 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [5]),
        .O(\bdatw[31]_INST_0_i_139_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [15]),
        .I5(\rgf/bank02/gr23 [15]),
        .O(\bdatw[31]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF77FF7FD5)) 
    \bdatw[31]_INST_0_i_140 
       (.I0(\bdatw[31]_INST_0_i_84_n_0 ),
        .I1(\fch/ir1 [12]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [15]),
        .O(\bdatw[31]_INST_0_i_140_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000800080)) 
    \bdatw[31]_INST_0_i_141 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [11]),
        .O(\bdatw[31]_INST_0_i_141_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_142 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .O(\bdatw[31]_INST_0_i_142_n_0 ));
  LUT5 #(
    .INIT(32'hFFEEFEEE)) 
    \bdatw[31]_INST_0_i_143 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .O(\bdatw[31]_INST_0_i_143_n_0 ));
  LUT6 #(
    .INIT(64'h60000000FFFFFFFF)) 
    \bdatw[31]_INST_0_i_144 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [11]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\bcmd[1]_INST_0_i_13_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_31_n_0 ),
        .I5(\badr[15]_INST_0_i_147_n_0 ),
        .O(\bdatw[31]_INST_0_i_144_n_0 ));
  LUT6 #(
    .INIT(64'h0E0E0E0E0E0E000E)) 
    \bdatw[31]_INST_0_i_145 
       (.I0(\bdatw[31]_INST_0_i_169_n_0 ),
        .I1(\bdatw[31]_INST_0_i_170_n_0 ),
        .I2(\bdatw[31]_INST_0_i_171_n_0 ),
        .I3(\bdatw[31]_INST_0_i_172_n_0 ),
        .I4(\badr[31]_INST_0_i_146_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .O(\bdatw[31]_INST_0_i_145_n_0 ));
  LUT6 #(
    .INIT(64'hEC30A333A000A000)) 
    \bdatw[31]_INST_0_i_146 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(\fch/ir1 [7]),
        .O(\bdatw[31]_INST_0_i_146_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \bdatw[31]_INST_0_i_147 
       (.I0(\fch/ir1 [10]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(div_crdy1),
        .O(\bdatw[31]_INST_0_i_147_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \bdatw[31]_INST_0_i_148 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\bdatw[31]_INST_0_i_173_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .O(\bdatw[31]_INST_0_i_148_n_0 ));
  LUT5 #(
    .INIT(32'h20004040)) 
    \bdatw[31]_INST_0_i_149 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .I2(div_crdy1),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [8]),
        .O(\bdatw[31]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_15 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [15]),
        .I5(\rgf/bank02/gr21 [15]),
        .O(\bdatw[31]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0002000F0A020A0A)) 
    \bdatw[31]_INST_0_i_150 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [10]),
        .O(\bdatw[31]_INST_0_i_150_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_151 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [9]),
        .O(\bdatw[31]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'h00FFAFF0C000AFF0)) 
    \bdatw[31]_INST_0_i_152 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [6]),
        .O(\bdatw[31]_INST_0_i_152_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_153 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .O(\bdatw[31]_INST_0_i_153_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFBFFFD)) 
    \bdatw[31]_INST_0_i_154 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [1]),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\ctl1/stat_reg_n_0_[1] ),
        .O(\bdatw[31]_INST_0_i_154_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[31]_INST_0_i_155 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .O(\bdatw[31]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFBFFFB)) 
    \bdatw[31]_INST_0_i_156 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [9]),
        .O(\bdatw[31]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'hBF7F4F7FFFFFFFFF)) 
    \bdatw[31]_INST_0_i_157 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [3]),
        .I5(\stat[2]_i_15_n_0 ),
        .O(\bdatw[31]_INST_0_i_157_n_0 ));
  LUT6 #(
    .INIT(64'h080F0F0F00000000)) 
    \bdatw[31]_INST_0_i_158 
       (.I0(div_crdy0),
        .I1(crdy),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [10]),
        .O(\bdatw[31]_INST_0_i_158_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFFFFFF)) 
    \bdatw[31]_INST_0_i_159 
       (.I0(\rgf_selc0_rn_wb[0]_i_31_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [10]),
        .I4(\bbus_o[5]_INST_0_i_24_n_0 ),
        .I5(\bdatw[31]_INST_0_i_174_n_0 ),
        .O(\bdatw[31]_INST_0_i_159_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_16 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [15]),
        .I5(\rgf/bank02/gr27 [15]),
        .O(\bdatw[31]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \bdatw[31]_INST_0_i_160 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [10]),
        .O(\bdatw[31]_INST_0_i_160_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \bdatw[31]_INST_0_i_161 
       (.I0(stat[0]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .O(\bdatw[31]_INST_0_i_161_n_0 ));
  LUT6 #(
    .INIT(64'hF350F0CCF30FF000)) 
    \bdatw[31]_INST_0_i_162 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [7]),
        .O(\bdatw[31]_INST_0_i_162_n_0 ));
  LUT6 #(
    .INIT(64'h9AFF6B7F3DFDFFFF)) 
    \bdatw[31]_INST_0_i_163 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [6]),
        .O(\bdatw[31]_INST_0_i_163_n_0 ));
  LUT6 #(
    .INIT(64'hF03000C0C0B000B0)) 
    \bdatw[31]_INST_0_i_164 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [9]),
        .O(\bdatw[31]_INST_0_i_164_n_0 ));
  LUT6 #(
    .INIT(64'h0004000004000000)) 
    \bdatw[31]_INST_0_i_165 
       (.I0(\fch/ir0 [8]),
        .I1(stat[0]),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [11]),
        .O(\bdatw[31]_INST_0_i_165_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF33B3FFFFF3B3)) 
    \bdatw[31]_INST_0_i_166 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\bdatw[31]_INST_0_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hB7FF3F77FFFFFFFF)) 
    \bdatw[31]_INST_0_i_167 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [3]),
        .I5(\stat[2]_i_15_n_0 ),
        .O(\bdatw[31]_INST_0_i_167_n_0 ));
  LUT3 #(
    .INIT(8'h94)) 
    \bdatw[31]_INST_0_i_168 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .O(\bdatw[31]_INST_0_i_168_n_0 ));
  LUT4 #(
    .INIT(16'h6FFF)) 
    \bdatw[31]_INST_0_i_169 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [7]),
        .O(\bdatw[31]_INST_0_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_17 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [15]),
        .I5(\rgf/bank02/gr25 [15]),
        .O(\bdatw[31]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h84C10000)) 
    \bdatw[31]_INST_0_i_170 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [9]),
        .O(\bdatw[31]_INST_0_i_170_n_0 ));
  LUT6 #(
    .INIT(64'h0F3000BC0FF30FFF)) 
    \bdatw[31]_INST_0_i_171 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [8]),
        .O(\bdatw[31]_INST_0_i_171_n_0 ));
  LUT3 #(
    .INIT(8'h94)) 
    \bdatw[31]_INST_0_i_172 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .O(\bdatw[31]_INST_0_i_172_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_173 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [4]),
        .O(\bdatw[31]_INST_0_i_173_n_0 ));
  LUT5 #(
    .INIT(32'h00F9003B)) 
    \bdatw[31]_INST_0_i_174 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [6]),
        .O(\bdatw[31]_INST_0_i_174_n_0 ));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \bdatw[31]_INST_0_i_18 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[2]),
        .O(\rgf/b0bus_sel_cr [4]));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \bdatw[31]_INST_0_i_19 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[31]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[31]_INST_0_i_9_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[31]_INST_0_i_10_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [31]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[31]));
  LUT6 #(
    .INIT(64'h0000004000000000)) 
    \bdatw[31]_INST_0_i_20 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_n_0 ),
        .I2(ctl_selb0_0),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_cr [2]));
  LUT6 #(
    .INIT(64'h00000000FFFF5551)) 
    \bdatw[31]_INST_0_i_23 
       (.I0(\bdatw[31]_INST_0_i_63_n_0 ),
        .I1(\bdatw[31]_INST_0_i_64_n_0 ),
        .I2(\bdatw[31]_INST_0_i_65_n_0 ),
        .I3(\bdatw[31]_INST_0_i_66_n_0 ),
        .I4(\bdatw[31]_INST_0_i_67_n_0 ),
        .I5(\bdatw[31]_INST_0_i_68_n_0 ),
        .O(ctl_selb0_0));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_24 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [15]),
        .O(\bdatw[31]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h8888B888BBBBBBBB)) 
    \bdatw[31]_INST_0_i_25 
       (.I0(\bdatw[31]_INST_0_i_69_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\ccmd[1]_INST_0_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_70_n_0 ),
        .I4(\bdatw[31]_INST_0_i_71_n_0 ),
        .I5(\bdatw[31]_INST_0_i_72_n_0 ),
        .O(\bdatw[31]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004440404)) 
    \bdatw[31]_INST_0_i_26 
       (.I0(\bdatw[31]_INST_0_i_73_n_0 ),
        .I1(\bdatw[31]_INST_0_i_74_n_0 ),
        .I2(\ccmd[0]_INST_0_i_13_n_0 ),
        .I3(\bdatw[31]_INST_0_i_75_n_0 ),
        .I4(\bdatw[31]_INST_0_i_76_n_0 ),
        .I5(\bdatw[31]_INST_0_i_77_n_0 ),
        .O(\bdatw[31]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0030AA000000AA00)) 
    \bdatw[31]_INST_0_i_27 
       (.I0(\bdatw[31]_INST_0_i_78_n_0 ),
        .I1(\bdatw[31]_INST_0_i_79_n_0 ),
        .I2(\bdatw[31]_INST_0_i_80_n_0 ),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .O(\bdatw[31]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hF000440000004400)) 
    \bdatw[31]_INST_0_i_28 
       (.I0(\bdatw[31]_INST_0_i_81_n_0 ),
        .I1(\badr[31]_INST_0_i_60_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [12]),
        .O(\bdatw[31]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA8A8A8A8A8AA)) 
    \bdatw[31]_INST_0_i_29 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\bdatw[31]_INST_0_i_82_n_0 ),
        .I2(\bdatw[31]_INST_0_i_83_n_0 ),
        .I3(\bdatw[31]_INST_0_i_84_n_0 ),
        .I4(\bdatw[31]_INST_0_i_85_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(ctl_selb1_0[2]));
  LUT3 #(
    .INIT(8'h10)) 
    \bdatw[31]_INST_0_i_3 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[31]_INST_0_i_13_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_2_n_0 ),
        .O(\bdatw[31]_INST_0_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \bdatw[31]_INST_0_i_30 
       (.I0(\bdatw[31]_INST_0_i_12_n_0 ),
        .I1(ctl_selb1_0[1]),
        .I2(\fch/ir1 [10]),
        .O(\bdatw[31]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_31 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .I4(\rgf/bank02/gr24 [15]),
        .I5(\rgf/bank02/gr23 [15]),
        .O(\bdatw[31]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_32 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank02/gr22 [15]),
        .I5(\rgf/bank02/gr21 [15]),
        .O(\bdatw[31]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_33 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .I3(\rgf/b1bus_sel_0 [0]),
        .I4(\rgf/bank02/gr20 [15]),
        .I5(\rgf/bank02/gr27 [15]),
        .O(\bdatw[31]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_34 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank02/gr26 [15]),
        .I5(\rgf/bank02/gr25 [15]),
        .O(\bdatw[31]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[31]_INST_0_i_35 
       (.I0(ctl_selb1_rn[1]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .O(\rgf/b1bus_sel_cr [4]));
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \bdatw[31]_INST_0_i_36 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_0[1]),
        .I4(\bdatw[31]_INST_0_i_12_n_0 ),
        .I5(ctl_selb1_0[2]),
        .O(\rgf/b1bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \bdatw[31]_INST_0_i_37 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_0[1]),
        .I4(\bdatw[31]_INST_0_i_12_n_0 ),
        .I5(ctl_selb1_0[2]),
        .O(\rgf/b1bus_sel_cr [2]));
  LUT6 #(
    .INIT(64'h00000000F4F4F000)) 
    \bdatw[31]_INST_0_i_40 
       (.I0(\bdatw[31]_INST_0_i_100_n_0 ),
        .I1(\bdatw[31]_INST_0_i_101_n_0 ),
        .I2(\bdatw[31]_INST_0_i_102_n_0 ),
        .I3(\bdatw[31]_INST_0_i_103_n_0 ),
        .I4(\bdatw[31]_INST_0_i_104_n_0 ),
        .I5(\bcmd[3]_INST_0_i_4_n_0 ),
        .O(ctl_selb1_0[1]));
  LUT6 #(
    .INIT(64'h0000000045450045)) 
    \bdatw[31]_INST_0_i_41 
       (.I0(\bdatw[31]_INST_0_i_105_n_0 ),
        .I1(\bdatw[31]_INST_0_i_106_n_0 ),
        .I2(\bdatw[31]_INST_0_i_107_n_0 ),
        .I3(\bdatw[31]_INST_0_i_108_n_0 ),
        .I4(\bdatw[31]_INST_0_i_109_n_0 ),
        .I5(\bdatw[31]_INST_0_i_110_n_0 ),
        .O(\bdatw[31]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'h40FF4040)) 
    \bdatw[31]_INST_0_i_42 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\bdatw[31]_INST_0_i_111_n_0 ),
        .I3(\bdatw[31]_INST_0_i_112_n_0 ),
        .I4(\bdatw[31]_INST_0_i_113_n_0 ),
        .O(\bdatw[31]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF00FFFFFF7F)) 
    \bdatw[31]_INST_0_i_43 
       (.I0(\bdatw[31]_INST_0_i_110_n_0 ),
        .I1(\fch/ir1 [14]),
        .I2(\bcmd[2]_INST_0_i_5_n_0 ),
        .I3(\fch/ir1 [15]),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\rgf_selc1_wb[0]_i_4_n_0 ),
        .O(\bdatw[31]_INST_0_i_43_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_44 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [14]),
        .O(\bdatw[31]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBB8B8B8B88)) 
    \bdatw[31]_INST_0_i_45 
       (.I0(\bdatw[31]_INST_0_i_114_n_0 ),
        .I1(\fch/ir1 [12]),
        .I2(\bdatw[31]_INST_0_i_115_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\bdatw[31]_INST_0_i_116_n_0 ),
        .I5(\stat[1]_i_12__0_n_0 ),
        .O(\bdatw[31]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_46 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_0 [3]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_47 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[0]),
        .I4(ctl_selb0_rn[2]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_0 [4]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_48 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_0 [1]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_49 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[1]),
        .I5(ctl_selb0_rn[0]),
        .O(\rgf/b0bus_sel_0 [2]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_50 
       (.I0(ctl_selb0_rn[2]),
        .I1(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I2(ctl_selb0_0),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_0 [7]));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \bdatw[31]_INST_0_i_51 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[2]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[1]),
        .O(\rgf/b0bus_sel_0 [0]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_52 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[1]),
        .I4(ctl_selb0_rn[0]),
        .I5(ctl_selb0_rn[2]),
        .O(\rgf/b0bus_sel_0 [5]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_53 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .I3(ctl_selb0_rn[0]),
        .I4(ctl_selb0_rn[1]),
        .I5(ctl_selb0_rn[2]),
        .O(\rgf/b0bus_sel_0 [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFF30500000)) 
    \bdatw[31]_INST_0_i_54 
       (.I0(\bdatw[31]_INST_0_i_117_n_0 ),
        .I1(\bdatw[31]_INST_0_i_118_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(\bdatw[31]_INST_0_i_119_n_0 ),
        .I5(\bdatw[31]_INST_0_i_120_n_0 ),
        .O(ctl_selb0_rn[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFA20000)) 
    \bdatw[31]_INST_0_i_55 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\bdatw[31]_INST_0_i_121_n_0 ),
        .I2(\bdatw[31]_INST_0_i_122_n_0 ),
        .I3(\badr[31]_INST_0_i_129_n_0 ),
        .I4(\badr[31]_INST_0_i_60_n_0 ),
        .I5(\bdatw[31]_INST_0_i_123_n_0 ),
        .O(ctl_selb0_rn[0]));
  LUT6 #(
    .INIT(64'h750075007500FFFF)) 
    \bdatw[31]_INST_0_i_56 
       (.I0(\bdatw[31]_INST_0_i_124_n_0 ),
        .I1(\bdatw[31]_INST_0_i_125_n_0 ),
        .I2(\fch/ir0 [2]),
        .I3(\bdatw[31]_INST_0_i_119_n_0 ),
        .I4(\bdatw[31]_INST_0_i_126_n_0 ),
        .I5(stat[2]),
        .O(ctl_selb0_rn[2]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_59 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [15]),
        .I5(\rgf/bank13/gr21 [15]),
        .O(\bdatw[31]_INST_0_i_59_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_6 
       (.I0(ctl_selb0_0),
        .I1(\bbus_o[5]_INST_0_i_2_n_0 ),
        .O(\bdatw[31]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_62 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [5]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [15]),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\bdatw[31]_INST_0_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hBBFB)) 
    \bdatw[31]_INST_0_i_63 
       (.I0(stat[1]),
        .I1(\fch/ir0 [13]),
        .I2(stat[0]),
        .I3(\bdatw[31]_INST_0_i_78_n_0 ),
        .O(\bdatw[31]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hABAFAFAFBBBFFFFF)) 
    \bdatw[31]_INST_0_i_64 
       (.I0(\fch/ir0 [11]),
        .I1(\bdatw[31]_INST_0_i_127_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\fch/ir0 [7]),
        .I5(\bdatw[31]_INST_0_i_128_n_0 ),
        .O(\bdatw[31]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8A8A8AAA8A8)) 
    \bdatw[31]_INST_0_i_65 
       (.I0(\fch/ir0 [11]),
        .I1(\bdatw[31]_INST_0_i_129_n_0 ),
        .I2(\bdatw[31]_INST_0_i_130_n_0 ),
        .I3(\bdatw[31]_INST_0_i_131_n_0 ),
        .I4(\bdatw[31]_INST_0_i_132_n_0 ),
        .I5(\bdatw[31]_INST_0_i_133_n_0 ),
        .O(\bdatw[31]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEEEEEEFEEEEEE)) 
    \bdatw[31]_INST_0_i_66 
       (.I0(\bdatw[31]_INST_0_i_134_n_0 ),
        .I1(\bdatw[31]_INST_0_i_78_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .I5(\ccmd[2]_INST_0_i_5_n_0 ),
        .O(\bdatw[31]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \bdatw[31]_INST_0_i_67 
       (.I0(\bcmd[1]_INST_0_i_28_n_0 ),
        .I1(\bdatw[31]_INST_0_i_135_n_0 ),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [1]),
        .I4(\ccmd[1]_INST_0_i_13_n_0 ),
        .I5(\bdatw[31]_INST_0_i_79_n_0 ),
        .O(\bdatw[31]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h77747777FFFFFFFF)) 
    \bdatw[31]_INST_0_i_68 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [2]),
        .I3(\bdatw[31]_INST_0_i_136_n_0 ),
        .I4(\bcmd[1]_INST_0_i_28_n_0 ),
        .I5(\bcmd[1]_INST_0_i_3_n_0 ),
        .O(\bdatw[31]_INST_0_i_68_n_0 ));
  LUT5 #(
    .INIT(32'h8A80202A)) 
    \bdatw[31]_INST_0_i_69 
       (.I0(\bbus_o[5]_INST_0_i_8_n_0 ),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [13]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir0 [11]),
        .O(\bdatw[31]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h0000770777777777)) 
    \bdatw[31]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_24_n_0 ),
        .I1(\bdatw[31]_INST_0_i_25_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I3(\bdatw[31]_INST_0_i_26_n_0 ),
        .I4(\bdatw[31]_INST_0_i_27_n_0 ),
        .I5(\bdatw[31]_INST_0_i_28_n_0 ),
        .O(\bdatw[31]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[31]_INST_0_i_70 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [2]),
        .I2(stat[0]),
        .I3(\fch/ir0 [13]),
        .O(\bdatw[31]_INST_0_i_70_n_0 ));
  LUT4 #(
    .INIT(16'hF9EF)) 
    \bdatw[31]_INST_0_i_71 
       (.I0(stat[2]),
        .I1(stat[1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .O(\bdatw[31]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF2FFFD)) 
    \bdatw[31]_INST_0_i_72 
       (.I0(\fch/ir0 [13]),
        .I1(\rgf/sreg/sr [6]),
        .I2(stat[0]),
        .I3(stat[1]),
        .I4(\fch/ir0 [11]),
        .I5(stat[2]),
        .O(\bdatw[31]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAABAAAAAAAAA)) 
    \bdatw[31]_INST_0_i_73 
       (.I0(\bdatw[31]_INST_0_i_137_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(ctl_fetch0_fl_i_28_n_0),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [9]),
        .O(\bdatw[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hFBAABBAAFBFBFBFB)) 
    \bdatw[31]_INST_0_i_74 
       (.I0(\ccmd[1]_INST_0_i_13_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\bdatw[31]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h2FCF20CF0FC00FC0)) 
    \bdatw[31]_INST_0_i_75 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\fch/ir0 [7]),
        .O(\bdatw[31]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFB79FFFFFFFFFFFF)) 
    \bdatw[31]_INST_0_i_76 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [6]),
        .O(\bdatw[31]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'h15404015)) 
    \bdatw[31]_INST_0_i_77 
       (.I0(\fch/ir0 [13]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [12]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\fch/ir0 [11]),
        .O(\bdatw[31]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h2800000000000000)) 
    \bdatw[31]_INST_0_i_78 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [6]),
        .I5(\bdatw[31]_INST_0_i_138_n_0 ),
        .O(\bdatw[31]_INST_0_i_78_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bdatw[31]_INST_0_i_79 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [4]),
        .O(\bdatw[31]_INST_0_i_79_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_8 
       (.I0(ctl_selb1_0[2]),
        .I1(\bdatw[31]_INST_0_i_30_n_0 ),
        .O(\bdatw[31]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0_i_80 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [3]),
        .O(\bdatw[31]_INST_0_i_80_n_0 ));
  LUT4 #(
    .INIT(16'h9666)) 
    \bdatw[31]_INST_0_i_81 
       (.I0(\fch/ir0 [11]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [12]),
        .I3(\rgf/sreg/sr [7]),
        .O(\bdatw[31]_INST_0_i_81_n_0 ));
  LUT4 #(
    .INIT(16'h2AAA)) 
    \bdatw[31]_INST_0_i_82 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [14]),
        .O(\bdatw[31]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055D55555)) 
    \bdatw[31]_INST_0_i_83 
       (.I0(\fch/ir1 [14]),
        .I1(\bdatw[31]_INST_0_i_139_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I3(\stat[1]_i_22_n_0 ),
        .I4(\fch/ir1 [8]),
        .I5(\bdatw[31]_INST_0_i_140_n_0 ),
        .O(\bdatw[31]_INST_0_i_83_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \bdatw[31]_INST_0_i_84 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\rgf/sreg/sr [6]),
        .O(\bdatw[31]_INST_0_i_84_n_0 ));
  LUT5 #(
    .INIT(32'h5FA0CFCF)) 
    \bdatw[31]_INST_0_i_85 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\fch/ir1 [14]),
        .O(\bdatw[31]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_86 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sel_0 [3]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_87 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_rn[0]),
        .I4(ctl_selb1_rn[2]),
        .I5(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sel_0 [4]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_88 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sel_0 [1]));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \bdatw[31]_INST_0_i_89 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[1]),
        .I5(ctl_selb1_rn[0]),
        .O(\rgf/b1bus_sel_0 [2]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_90 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(ctl_selb1_0[1]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sel_0 [7]));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \bdatw[31]_INST_0_i_91 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_rn[2]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sel_0 [0]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_92 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_rn[1]),
        .I4(ctl_selb1_rn[0]),
        .I5(ctl_selb1_rn[2]),
        .O(\rgf/b1bus_sel_0 [5]));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \bdatw[31]_INST_0_i_93 
       (.I0(ctl_selb1_0[2]),
        .I1(ctl_selb1_0[1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_rn[0]),
        .I4(ctl_selb1_rn[1]),
        .I5(ctl_selb1_rn[2]),
        .O(\rgf/b1bus_sel_0 [6]));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_96 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [1]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .I4(\rgf/bank13/gr22 [15]),
        .I5(\rgf/bank13/gr21 [15]),
        .O(\bdatw[31]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_99 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [5]),
        .I3(\rgf/b1bus_sel_0 [6]),
        .I4(\rgf/bank13/gr26 [15]),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\bdatw[31]_INST_0_i_99_n_0 ));
  LUT3 #(
    .INIT(8'h07)) 
    \bdatw[3]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[11]_INST_0_i_3_n_0 ),
        .O(bdatw[3]));
  LUT3 #(
    .INIT(8'h07)) 
    \bdatw[4]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[12]_INST_0_i_1_n_0 ),
        .O(bdatw[4]));
  LUT3 #(
    .INIT(8'h07)) 
    \bdatw[5]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[13]_INST_0_i_1_n_0 ),
        .O(bdatw[5]));
  LUT3 #(
    .INIT(8'h07)) 
    \bdatw[6]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[14]_INST_0_i_3_n_0 ),
        .O(bdatw[6]));
  LUT3 #(
    .INIT(8'h70)) 
    \bdatw[7]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_1_n_0 ),
        .I2(\bdatw[15]_INST_0_i_5_n_0 ),
        .O(bdatw[7]));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[8]_INST_0 
       (.I0(\bdatw[8]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(b1bus_0[8]),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(b0bus_0[8]),
        .O(bdatw[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\bdatw[8]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_10 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [0]),
        .O(\bdatw[8]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_4_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[8]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[8]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [8]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[8]));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[8]_INST_0_i_21 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [1]),
        .O(\bdatw[8]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_22 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [0]),
        .O(\bdatw[8]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEEFEEE)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(\rgf/b0bus_out/bdatw[8]_INST_0_i_7_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[8]_INST_0_i_8_n_0 ),
        .I2(\bdatw[31]_INST_0_i_6_n_0 ),
        .I3(\fch/eir [8]),
        .I4(\bdatw[31]_INST_0_i_7_n_0 ),
        .I5(\bdatw[8]_INST_0_i_9_n_0 ),
        .O(b0bus_0[8]));
  LUT6 #(
    .INIT(64'h0C000000C0CC8888)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(\fch/ir1 [7]),
        .I1(ctl_selb1_0[2]),
        .I2(\bdatw[9]_INST_0_i_10_n_0 ),
        .I3(\bdatw[8]_INST_0_i_10_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(\bdatw[8]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0C000000C0CC8888)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(\fch/ir0 [7]),
        .I1(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I2(\bdatw[8]_INST_0_i_21_n_0 ),
        .I3(\bdatw[8]_INST_0_i_22_n_0 ),
        .I4(ctl_selb0_0),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[8]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444F44)) 
    \bdatw[9]_INST_0 
       (.I0(\bdatw[9]_INST_0_i_1_n_0 ),
        .I1(\bdatw[15]_INST_0_i_4_n_0 ),
        .I2(\bdatw[15]_INST_0_i_1_n_0 ),
        .I3(b1bus_0[9]),
        .I4(\bcmd[0]_INST_0_i_3_n_0 ),
        .I5(b0bus_0[9]),
        .O(bdatw[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .O(\bdatw[9]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[9]_INST_0_i_10 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [1]),
        .O(\bdatw[9]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[9]_INST_0_i_11 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [0]),
        .O(\bdatw[9]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[9]_INST_0_i_17 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .O(\bdatw[9]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(\bdatw[9]_INST_0_i_4_n_0 ),
        .I1(\rgf/b1bus_out/bdatw[9]_INST_0_i_5_n_0 ),
        .I2(\rgf/b1bus_out/bdatw[9]_INST_0_i_6_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [9]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[9]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(\bdatw[9]_INST_0_i_7_n_0 ),
        .I1(\rgf/b0bus_out/bdatw[9]_INST_0_i_8_n_0 ),
        .I2(\rgf/b0bus_out/bdatw[9]_INST_0_i_9_n_0 ),
        .I3(\bdatw[31]_INST_0_i_6_n_0 ),
        .I4(\fch/eir [9]),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(b0bus_0[9]));
  LUT6 #(
    .INIT(64'h00A00000A808A8A8)) 
    \bdatw[9]_INST_0_i_4 
       (.I0(ctl_selb1_0[2]),
        .I1(\fch/ir1 [8]),
        .I2(ctl_selb1_0[1]),
        .I3(\bdatw[9]_INST_0_i_10_n_0 ),
        .I4(\bdatw[9]_INST_0_i_11_n_0 ),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(\bdatw[9]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hA000000008A8A8A8)) 
    \bdatw[9]_INST_0_i_7 
       (.I0(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(ctl_selb0_0),
        .I3(\bdatw[9]_INST_0_i_17_n_0 ),
        .I4(\bdatw[11]_INST_0_i_19_n_0 ),
        .I5(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(\bdatw[9]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(ccmd[0]));
  LUT6 #(
    .INIT(64'hBBBBBBBBABABABAA)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(stat[2]),
        .I1(\ccmd[0]_INST_0_i_2_n_0 ),
        .I2(\ccmd[0]_INST_0_i_3_n_0 ),
        .I3(\ccmd[0]_INST_0_i_4_n_0 ),
        .I4(\ccmd[0]_INST_0_i_5_n_0 ),
        .I5(\ccmd[0]_INST_0_i_6_n_0 ),
        .O(\ccmd[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0011010000110000)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(stat[1]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [15]),
        .I5(\rgf/sreg/sr [6]),
        .O(\ccmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(\fch/ir0 [14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\fch/ir0 [12]),
        .I4(\rgf/sreg/sr [6]),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hAA2A0A0AAA2AA020)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(\ccmd[0]_INST_0_i_25_n_0 ),
        .I1(\ccmd[3]_INST_0_i_15_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [14]),
        .I5(\rgf/sreg/sr [7]),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [8]),
        .O(\ccmd[0]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[0]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h40000020)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [4]),
        .O(\ccmd[0]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFD0DFD)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .O(\ccmd[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h77CD77DD73DC73DC)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(stat[1]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\fch/ir0 [6]),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h600C)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[0]_INST_0_i_19 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFEFEFE00FEFE)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(\ccmd[0]_INST_0_i_7_n_0 ),
        .I1(\ccmd[0]_INST_0_i_8_n_0 ),
        .I2(\ccmd[0]_INST_0_i_9_n_0 ),
        .I3(\ccmd[0]_INST_0_i_10_n_0 ),
        .I4(\fch/ir0 [13]),
        .I5(\ccmd[0]_INST_0_i_11_n_0 ),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_20 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .O(\ccmd[0]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \ccmd[0]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir0 [12]),
        .I2(\rgf/sreg/sr [5]),
        .O(\ccmd[0]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \ccmd[0]_INST_0_i_22 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .O(\ccmd[0]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \ccmd[0]_INST_0_i_23 
       (.I0(\ccmd[2]_INST_0_i_18_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [8]),
        .I3(\fadr[15]_INST_0_i_12_n_0 ),
        .I4(\fch/ir0 [9]),
        .I5(stat[1]),
        .O(\ccmd[0]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[0]_INST_0_i_24 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [10]),
        .O(\ccmd[0]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF70FFFFFF)) 
    \ccmd[0]_INST_0_i_25 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [9]),
        .O(\ccmd[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0C05000500050005)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(\ccmd[0]_INST_0_i_12_n_0 ),
        .I1(\ccmd[0]_INST_0_i_13_n_0 ),
        .I2(stat[1]),
        .I3(stat[0]),
        .I4(\ccmd[0]_INST_0_i_14_n_0 ),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFFFCF3A0AFACA)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(\ccmd[0]_INST_0_i_16_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [10]),
        .I3(\ccmd[0]_INST_0_i_17_n_0 ),
        .I4(\ccmd[0]_INST_0_i_18_n_0 ),
        .I5(stat[1]),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEEFAAAABFAEAAAA)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(stat[0]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [6]),
        .I4(\ccmd[0]_INST_0_i_19_n_0 ),
        .I5(\fch/ir0 [3]),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEEFFFFFEF)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(\ccmd[0]_INST_0_i_20_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [14]),
        .O(\ccmd[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000020002020002)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(\fch/ir0 [14]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\ccmd[0]_INST_0_i_21_n_0 ),
        .I4(\fch/ir0 [15]),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF80)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(\ccmd[0]_INST_0_i_22_n_0 ),
        .I1(\bdatw[8]_INST_0_i_22_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I3(\ccmd[0]_INST_0_i_23_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(\ccmd[0]_INST_0_i_24_n_0 ),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4444404040044040)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(\fch/ir0 [14]),
        .I1(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir0 [12]),
        .I5(\fch/ir0 [15]),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'h2222222202222222)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_2_n_0 ),
        .I1(\ccmd[1]_INST_0_i_3_n_0 ),
        .I2(\ccmd[1]_INST_0_i_4_n_0 ),
        .I3(\ccmd[1]_INST_0_i_5_n_0 ),
        .I4(\ccmd[1]_INST_0_i_6_n_0 ),
        .I5(\ccmd[1]_INST_0_i_7_n_0 ),
        .O(\ccmd[1]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [7]),
        .O(\ccmd[1]_INST_0_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(div_crdy0),
        .I1(crdy),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [11]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(\ccmd[1]_INST_0_i_16_n_0 ),
        .I1(\ccmd[1]_INST_0_i_17_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\bbus_o[5]_INST_0_i_9_n_0 ),
        .O(\ccmd[1]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h3302C0F302028002)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [11]),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0002280808000800)) 
    \ccmd[1]_INST_0_i_15 
       (.I0(\ccmd[0]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [6]),
        .O(\ccmd[1]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \ccmd[1]_INST_0_i_16 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [8]),
        .O(\ccmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBFFFFF)) 
    \ccmd[1]_INST_0_i_17 
       (.I0(stat[0]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(stat[2]),
        .I4(stat[1]),
        .I5(\fch/ir0 [15]),
        .O(\ccmd[1]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBABFBABFBABFAAAA)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(\bcmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[1]_INST_0_i_8_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\ccmd[1]_INST_0_i_9_n_0 ),
        .I4(\ccmd[1]_INST_0_i_10_n_0 ),
        .I5(\ccmd[1]_INST_0_i_11_n_0 ),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF73CF0000)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [14]),
        .I4(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I5(\ccmd[1]_INST_0_i_12_n_0 ),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0024)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .I2(stat[2]),
        .I3(\fch/ir0 [1]),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(\ccmd[1]_INST_0_i_13_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [7]),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(\fch/ir0 [15]),
        .I1(stat[0]),
        .I2(stat[1]),
        .O(\ccmd[1]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [14]),
        .O(\ccmd[1]_INST_0_i_7_n_0 ));
  MUXF7 \ccmd[1]_INST_0_i_8 
       (.I0(\ccmd[1]_INST_0_i_14_n_0 ),
        .I1(\ccmd[1]_INST_0_i_15_n_0 ),
        .O(\ccmd[1]_INST_0_i_8_n_0 ),
        .S(\fch/ir0 [9]));
  LUT6 #(
    .INIT(64'h25252F0515002A00)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [11]),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(ccmd[2]));
  LUT6 #(
    .INIT(64'h00000000EAEAAAEA)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(\ccmd[2]_INST_0_i_2_n_0 ),
        .I1(\ccmd[2]_INST_0_i_3_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\ccmd[2]_INST_0_i_4_n_0 ),
        .I4(\ccmd[2]_INST_0_i_5_n_0 ),
        .I5(\ccmd[2]_INST_0_i_6_n_0 ),
        .O(\ccmd[2]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(crdy),
        .I1(div_crdy0),
        .O(\ccmd[2]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFAFAFBEBFABAFBEB)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(\fch/ir0 [7]),
        .I1(stat[1]),
        .I2(\fch/ir0 [9]),
        .I3(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [3]),
        .O(\ccmd[2]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h020AA20A)) 
    \ccmd[2]_INST_0_i_13 
       (.I0(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [14]),
        .O(\ccmd[2]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF07A7FF0F)) 
    \ccmd[2]_INST_0_i_14 
       (.I0(\fch/ir0 [7]),
        .I1(\ccmd[4]_INST_0_i_1_n_0 ),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [6]),
        .I5(\ccmd[2]_INST_0_i_19_n_0 ),
        .O(\ccmd[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABAAAAAAAAAA)) 
    \ccmd[2]_INST_0_i_15 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [11]),
        .I3(stat[1]),
        .I4(\fch/ir0 [9]),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\ccmd[2]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h5444)) 
    \ccmd[2]_INST_0_i_16 
       (.I0(\fch/ir0 [11]),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(crdy),
        .I3(div_crdy0),
        .O(\ccmd[2]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h40004444)) 
    \ccmd[2]_INST_0_i_17 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(crdy),
        .I3(div_crdy0),
        .I4(\fch/ir0 [7]),
        .O(\ccmd[2]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[2]_INST_0_i_18 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .O(\ccmd[2]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[2]_INST_0_i_19 
       (.I0(stat[1]),
        .I1(\fch/ir0 [10]),
        .O(\ccmd[2]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFEE)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(\ccmd[2]_INST_0_i_7_n_0 ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(stat[1]),
        .I4(stat[2]),
        .I5(stat[0]),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h777F0000FFFFFFFF)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(\ccmd[2]_INST_0_i_9_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\ccmd[2]_INST_0_i_11_n_0 ),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\ccmd[2]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(\fch/ir0 [9]),
        .I1(crdy),
        .I2(div_crdy0),
        .I3(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAAAAAAAAAAA)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(\ccmd[2]_INST_0_i_13_n_0 ),
        .I1(\fch/ir0 [1]),
        .I2(stat[2]),
        .I3(stat[1]),
        .I4(\rgf_selc0_wb[1]_i_5_n_0 ),
        .I5(\ccmd[1]_INST_0_i_5_n_0 ),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h2222222222220222)) 
    \ccmd[2]_INST_0_i_7 
       (.I0(\ccmd[2]_INST_0_i_14_n_0 ),
        .I1(\ccmd[2]_INST_0_i_15_n_0 ),
        .I2(\ccmd[2]_INST_0_i_16_n_0 ),
        .I3(\ccmd[2]_INST_0_i_17_n_0 ),
        .I4(stat[1]),
        .I5(\ccmd[2]_INST_0_i_18_n_0 ),
        .O(\ccmd[2]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h37BF3F33)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [4]),
        .O(\ccmd[2]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(\fch/ir0 [7]),
        .I1(stat[1]),
        .O(\ccmd[2]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0 
       (.I0(ccmd[4]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(ccmd[3]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBAABA)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(stat[2]),
        .I1(\ccmd[3]_INST_0_i_2_n_0 ),
        .I2(stat[1]),
        .I3(\fch/ir0 [10]),
        .I4(\ccmd[3]_INST_0_i_3_n_0 ),
        .I5(\ccmd[3]_INST_0_i_4_n_0 ),
        .O(\ccmd[3]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(\fch/ir0 [2]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [12]),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [1]),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(stat[0]),
        .I1(\fch/ir0 [8]),
        .O(\ccmd[3]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h80808000FFFFFFFF)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [6]),
        .I2(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\ccmd[3]_INST_0_i_19_n_0 ),
        .O(\ccmd[3]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[3]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0800314000202010)) 
    \ccmd[3]_INST_0_i_17 
       (.I0(\fch/ir0 [4]),
        .I1(stat[0]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [3]),
        .O(\ccmd[3]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAEAAAAAAAA)) 
    \ccmd[3]_INST_0_i_18 
       (.I0(\ccmd[3]_INST_0_i_20_n_0 ),
        .I1(\bdatw[31]_INST_0_i_138_n_0 ),
        .I2(stat[0]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [6]),
        .O(\ccmd[3]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDDDDDFFFFFFF)) 
    \ccmd[3]_INST_0_i_19 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(\ccmd[3]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABAAAAABAAAA)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(\ccmd[3]_INST_0_i_5_n_0 ),
        .I1(\ccmd[3]_INST_0_i_6_n_0 ),
        .I2(\ccmd[3]_INST_0_i_7_n_0 ),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [3]),
        .I5(stat[1]),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h6200000022003300)) 
    \ccmd[3]_INST_0_i_20 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\ccmd[3]_INST_0_i_21_n_0 ),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [10]),
        .O(\ccmd[3]_INST_0_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_21 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[3]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [15]),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  MUXF7 \ccmd[3]_INST_0_i_4 
       (.I0(\ccmd[3]_INST_0_i_8_n_0 ),
        .I1(\ccmd[3]_INST_0_i_9_n_0 ),
        .O(\ccmd[3]_INST_0_i_4_n_0 ),
        .S(\fch/ir0 [11]));
  LUT6 #(
    .INIT(64'h0080880008880000)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I1(\fch/ir0 [15]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [13]),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFFFFFFF)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(\ccmd[3]_INST_0_i_10_n_0 ),
        .I1(\ccmd[3]_INST_0_i_11_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [13]),
        .I4(\ccmd[3]_INST_0_i_12_n_0 ),
        .I5(\ccmd[3]_INST_0_i_13_n_0 ),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [4]),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7777777077777777)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(\ccmd[3]_INST_0_i_14_n_0 ),
        .I1(\ccmd[3]_INST_0_i_15_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(stat[0]),
        .I4(\ccmd[3]_INST_0_i_16_n_0 ),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\ccmd[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BFFFFFFF)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(stat[1]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [10]),
        .I4(\ccmd[3]_INST_0_i_17_n_0 ),
        .I5(\ccmd[3]_INST_0_i_18_n_0 ),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000AAAA08)) 
    \ccmd[4]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(stat[0]),
        .I4(stat[1]),
        .I5(\ccmd[4]_INST_0_i_3_n_0 ),
        .O(ccmd[4]));
  LUT3 #(
    .INIT(8'h08)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(div_crdy0),
        .I1(crdy),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\ccmd[4]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .O(\ccmd[4]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(stat[2]),
        .I1(\fch/ir0 [11]),
        .O(\ccmd[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFF)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [12]),
        .I5(\fch/ir0 [13]),
        .O(\ccmd[4]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h82FF8200)) 
    chg_quo_sgn_i_1
       (.I0(\alu0/div/dctl/dctl_sign ),
        .I1(chg_quo_sgn_i_2_n_0),
        .I2(\alu0/div/den2 ),
        .I3(\alu0/div/dctl/fsm/set_sgn ),
        .I4(\alu0/div/chg_quo_sgn ),
        .O(chg_quo_sgn_i_1_n_0));
  LUT5 #(
    .INIT(32'h82FF8200)) 
    chg_quo_sgn_i_1__0
       (.I0(\alu1/div/dctl/dctl_sign ),
        .I1(chg_quo_sgn_i_2__0_n_0),
        .I2(\alu1/div/den2 ),
        .I3(\alu1/div/dctl/fsm/set_sgn ),
        .I4(\alu1/div/chg_quo_sgn ),
        .O(chg_quo_sgn_i_1__0_n_0));
  LUT5 #(
    .INIT(32'h4540757F)) 
    chg_quo_sgn_i_2
       (.I0(\alu0/div/dso_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(div_crdy0),
        .I3(\alu0/div/dctl/dctl_long_f ),
        .I4(\alu0/div/dso_0 [15]),
        .O(chg_quo_sgn_i_2_n_0));
  LUT5 #(
    .INIT(32'h4540757F)) 
    chg_quo_sgn_i_2__0
       (.I0(\alu1/div/dso_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(div_crdy1),
        .I3(\alu1/div/dctl/dctl_long_f ),
        .I4(\alu1/div/dso_0 [15]),
        .O(chg_quo_sgn_i_2__0_n_0));
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    chg_rem_sgn_i_1
       (.I0(\alu0/div/dctl/fsm/chg_rem_sgn0 ),
        .I1(\alu0/div/dctl_stat [1]),
        .I2(\alu0/div/dctl_stat [2]),
        .I3(\alu0/div/dctl_stat [0]),
        .I4(\alu0/div/dctl_stat [3]),
        .I5(\alu0/div/chg_rem_sgn ),
        .O(chg_rem_sgn_i_1_n_0));
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    chg_rem_sgn_i_1__0
       (.I0(\alu1/div/dctl/fsm/chg_rem_sgn0 ),
        .I1(\alu1/div/dctl_stat [1]),
        .I2(\alu1/div/dctl_stat [2]),
        .I3(\alu1/div/dctl_stat [0]),
        .I4(\alu1/div/dctl_stat [3]),
        .I5(\alu1/div/chg_rem_sgn ),
        .O(chg_rem_sgn_i_1__0_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    chg_rem_sgn_i_2
       (.I0(\alu0/div/den2 ),
        .I1(\alu0/div/dctl/dctl_sign ),
        .O(\alu0/div/dctl/fsm/chg_rem_sgn0 ));
  LUT2 #(
    .INIT(4'h8)) 
    chg_rem_sgn_i_2__0
       (.I0(\alu1/div/den2 ),
        .I1(\alu1/div/dctl/dctl_sign ),
        .O(\alu1/div/dctl/fsm/chg_rem_sgn0 ));
  FDRE \ctl0/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl0/stat_nx [0]),
        .Q(stat[0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \ctl0/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl0/stat_nx [1]),
        .Q(stat[1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \ctl0/stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat[2]_i_1__1_n_0 ),
        .Q(stat[2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \ctl1/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl1/stat_nx [0]),
        .Q(\ctl1/stat_reg_n_0_[0] ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \ctl1/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl1/stat_nx [1]),
        .Q(\ctl1/stat_reg_n_0_[1] ),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \ctl1/stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ctl1/stat_nx [2]),
        .Q(\ctl1/stat_reg_n_0_[2] ),
        .R(\alu1/div/p_0_in__0 ));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_bcc_take0_fl_i_1
       (.I0(fch_term),
        .I1(rst_n),
        .O(ctl_bcc_take0_fl_i_1_n_0));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take0_fl_i_2
       (.I0(stat[0]),
        .I1(stat[2]),
        .I2(stat[1]),
        .I3(\fch/ctl_bcc_take0_fl ),
        .O(ctl_bcc_take0_fl_i_2_n_0));
  LUT4 #(
    .INIT(16'hFF80)) 
    ctl_bcc_take1_fl_i_1
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ctl_bcc_take1_fl ),
        .O(ctl_bcc_take1_fl_i_1_n_0));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    ctl_fetch0_fl_i_1
       (.I0(ctl_fetch0_fl_i_2_n_0),
        .I1(\fch/ir0 [11]),
        .I2(ctl_fetch0_fl_i_3_n_0),
        .I3(ctl_fetch0_fl_i_4_n_0),
        .I4(ctl_fetch0_fl_i_5_n_0),
        .I5(ctl_fetch0_fl_i_6_n_0),
        .O(ctl_fetch0));
  LUT6 #(
    .INIT(64'hF700FFFFF700F700)) 
    ctl_fetch0_fl_i_10
       (.I0(ctl_fetch0_fl_i_28_n_0),
        .I1(\fch/ir0 [12]),
        .I2(stat[1]),
        .I3(\ccmd[4]_INST_0_i_4_n_0 ),
        .I4(ctl_fetch0_fl_i_29_n_0),
        .I5(\ccmd[0]_INST_0_i_14_n_0 ),
        .O(ctl_fetch0_fl_i_10_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAFEAAAAAA)) 
    ctl_fetch0_fl_i_11
       (.I0(ctl_fetch0_fl_i_30_n_0),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(stat[0]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_11_n_0));
  LUT6 #(
    .INIT(64'h7FF000F00F000000)) 
    ctl_fetch0_fl_i_12
       (.I0(\fch/ir0 [6]),
        .I1(ctl_fetch0_fl_i_31_n_0),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .I5(ctl_fetch0_fl_i_32_n_0),
        .O(ctl_fetch0_fl_i_12_n_0));
  LUT6 #(
    .INIT(64'h7CFF70FF30FF30FF)) 
    ctl_fetch0_fl_i_13
       (.I0(ctl_fetch0_fl_i_33_n_0),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [14]),
        .I4(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I5(\fch/ir0 [9]),
        .O(ctl_fetch0_fl_i_13_n_0));
  LUT6 #(
    .INIT(64'h00300F3F40704070)) 
    ctl_fetch0_fl_i_14
       (.I0(\stat[1]_i_5__0_n_0 ),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [12]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\rgf/sreg/sr [6]),
        .I5(\fch/ir0 [13]),
        .O(ctl_fetch0_fl_i_14_n_0));
  LUT4 #(
    .INIT(16'h0800)) 
    ctl_fetch0_fl_i_15
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [13]),
        .O(ctl_fetch0_fl_i_15_n_0));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFFFEFE)) 
    ctl_fetch0_fl_i_16
       (.I0(ctl_fetch0_fl_i_34_n_0),
        .I1(stat[2]),
        .I2(stat[1]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [14]),
        .I5(\rgf/sreg/sr [5]),
        .O(ctl_fetch0_fl_i_16_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch0_fl_i_17
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [9]),
        .O(ctl_fetch0_fl_i_17_n_0));
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    ctl_fetch0_fl_i_18
       (.I0(stat[0]),
        .I1(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [11]),
        .I4(\bdatw[12]_INST_0_i_23_n_0 ),
        .I5(ctl_fetch0_fl_i_35_n_0),
        .O(ctl_fetch0_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'h000077D577D577D5)) 
    ctl_fetch0_fl_i_19
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [10]),
        .I4(stat[0]),
        .I5(ctl_fetch0_fl_i_36_n_0),
        .O(ctl_fetch0_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBABAAAA)) 
    ctl_fetch0_fl_i_2
       (.I0(ctl_fetch0_fl_i_7_n_0),
        .I1(ctl_fetch0_fl_i_8_n_0),
        .I2(ctl_fetch0_fl_i_9_n_0),
        .I3(ctl_fetch0_fl_i_10_n_0),
        .I4(\bcmd[2]_INST_0_i_8_n_0 ),
        .I5(ctl_fetch0_fl_i_11_n_0),
        .O(ctl_fetch0_fl_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    ctl_fetch0_fl_i_20
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(stat[2]),
        .I4(\fch/ir0 [15]),
        .O(ctl_fetch0_fl_i_20_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    ctl_fetch0_fl_i_21
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .O(ctl_fetch0_fl_i_21_n_0));
  LUT3 #(
    .INIT(8'h63)) 
    ctl_fetch0_fl_i_22
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [4]),
        .O(ctl_fetch0_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFF1FFFFF15155555)) 
    ctl_fetch0_fl_i_23
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [11]),
        .I2(ctl_fetch0_fl_i_27_n_0),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .I5(stat[1]),
        .O(ctl_fetch0_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'h00000000BAAABBAB)) 
    ctl_fetch0_fl_i_24
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\rgf/sreg/sr [5]),
        .I4(ctl_fetch0_fl_i_37_n_0),
        .I5(ctl_fetch0_fl_i_38_n_0),
        .O(ctl_fetch0_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'hAC00AC00AC000C00)) 
    ctl_fetch0_fl_i_25
       (.I0(ctl_fetch0_fl_i_39_n_0),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [13]),
        .I4(stat[0]),
        .I5(ctl_fetch0_fl_i_40_n_0),
        .O(ctl_fetch0_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hCDCDFDCDFDFDFDFD)) 
    ctl_fetch0_fl_i_26
       (.I0(ctl_fetch0_fl_i_41_n_0),
        .I1(ctl_fetch0_fl_i_42_n_0),
        .I2(\fch/ir0 [9]),
        .I3(stat[0]),
        .I4(\fch/ir0 [7]),
        .I5(\bcmd[1]_INST_0_i_6_n_0 ),
        .O(ctl_fetch0_fl_i_26_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_27
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_27_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch0_fl_i_28
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_28_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch0_fl_i_29
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00F2)) 
    ctl_fetch0_fl_i_3
       (.I0(ctl_fetch0_fl_i_12_n_0),
        .I1(ctl_fetch0_fl_i_13_n_0),
        .I2(\ccmd[0]_INST_0_i_20_n_0 ),
        .I3(ctl_fetch0_fl_i_14_n_0),
        .I4(ctl_fetch0_fl_i_15_n_0),
        .I5(ctl_fetch0_fl_i_16_n_0),
        .O(ctl_fetch0_fl_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFC4F4C4C4C4C4)) 
    ctl_fetch0_fl_i_30
       (.I0(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I1(stat[1]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(ctl_fetch0_fl_i_43_n_0),
        .I5(ctl_fetch0_fl_i_44_n_0),
        .O(ctl_fetch0_fl_i_30_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch0_fl_i_31
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [5]),
        .O(ctl_fetch0_fl_i_31_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00E0E0)) 
    ctl_fetch0_fl_i_32
       (.I0(\rgf/sreg/sr [11]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [7]),
        .O(ctl_fetch0_fl_i_32_n_0));
  LUT3 #(
    .INIT(8'hA9)) 
    ctl_fetch0_fl_i_33
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .O(ctl_fetch0_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'hAAAA0220AAAAAAAA)) 
    ctl_fetch0_fl_i_34
       (.I0(stat[0]),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [5]),
        .I4(ctl_fetch0_fl_i_45_n_0),
        .I5(ctl_fetch0_fl_i_46_n_0),
        .O(ctl_fetch0_fl_i_34_n_0));
  LUT4 #(
    .INIT(16'h0001)) 
    ctl_fetch0_fl_i_35
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [4]),
        .O(ctl_fetch0_fl_i_35_n_0));
  LUT3 #(
    .INIT(8'hD2)) 
    ctl_fetch0_fl_i_36
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [6]),
        .O(ctl_fetch0_fl_i_36_n_0));
  LUT6 #(
    .INIT(64'h8888AAAAAAAA8088)) 
    ctl_fetch0_fl_i_37
       (.I0(\stat[0]_i_8__0_n_0 ),
        .I1(\fch/ir0 [0]),
        .I2(fch_irq_req),
        .I3(irq),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [3]),
        .O(ctl_fetch0_fl_i_37_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF0CFF44FF)) 
    ctl_fetch0_fl_i_38
       (.I0(\rgf/sreg/sr [4]),
        .I1(\fch/ir0 [12]),
        .I2(\stat[1]_i_5__0_n_0 ),
        .I3(\bbus_o[5]_INST_0_i_8_n_0 ),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [13]),
        .O(ctl_fetch0_fl_i_38_n_0));
  LUT6 #(
    .INIT(64'hEEEEEEEEE000E0E0)) 
    ctl_fetch0_fl_i_39
       (.I0(ctl_fetch0_fl_i_47_n_0),
        .I1(\fch/ir0 [8]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(stat[0]),
        .I4(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(ctl_fetch0_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF008000FF)) 
    ctl_fetch0_fl_i_4
       (.I0(stat[0]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [3]),
        .I4(ctl_fetch0_fl_i_17_n_0),
        .I5(brdy),
        .O(ctl_fetch0_fl_i_4_n_0));
  LUT3 #(
    .INIT(8'hBF)) 
    ctl_fetch0_fl_i_40
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [10]),
        .O(ctl_fetch0_fl_i_40_n_0));
  LUT6 #(
    .INIT(64'h000000000C9E0000)) 
    ctl_fetch0_fl_i_41
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [3]),
        .I3(stat[1]),
        .I4(\bcmd[3]_INST_0_i_8_n_0 ),
        .I5(ctl_fetch0_fl_i_48_n_0),
        .O(ctl_fetch0_fl_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFFFFFE)) 
    ctl_fetch0_fl_i_42
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [9]),
        .I5(ctl_fetch0_fl_i_49_n_0),
        .O(ctl_fetch0_fl_i_42_n_0));
  LUT5 #(
    .INIT(32'hFEFFFFFF)) 
    ctl_fetch0_fl_i_43
       (.I0(\fch/ir0 [15]),
        .I1(stat[1]),
        .I2(stat[2]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [14]),
        .O(ctl_fetch0_fl_i_43_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    ctl_fetch0_fl_i_44
       (.I0(\fch/ir0 [15]),
        .I1(stat[0]),
        .I2(stat[2]),
        .O(ctl_fetch0_fl_i_44_n_0));
  LUT6 #(
    .INIT(64'h04F4FFFF04F400FF)) 
    ctl_fetch0_fl_i_45
       (.I0(\rgf/sreg/sr [10]),
        .I1(ctl_fetch0_fl_i_50_n_0),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [6]),
        .O(ctl_fetch0_fl_i_45_n_0));
  LUT6 #(
    .INIT(64'h2FFF2FF0FFFFFFFF)) 
    ctl_fetch0_fl_i_46
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [7]),
        .I4(\rgf/sreg/sr [11]),
        .I5(\fch/ir0 [8]),
        .O(ctl_fetch0_fl_i_46_n_0));
  LUT6 #(
    .INIT(64'h00D0000000000000)) 
    ctl_fetch0_fl_i_47
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\rgf/sreg/sr [10]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [7]),
        .I5(stat[0]),
        .O(ctl_fetch0_fl_i_47_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    ctl_fetch0_fl_i_48
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [5]),
        .I2(ctl_fetch0_fl_i_51_n_0),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [2]),
        .O(ctl_fetch0_fl_i_48_n_0));
  LUT5 #(
    .INIT(32'hAAAAAAA8)) 
    ctl_fetch0_fl_i_49
       (.I0(stat[2]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [9]),
        .O(ctl_fetch0_fl_i_49_n_0));
  LUT6 #(
    .INIT(64'h00000000BAAA0000)) 
    ctl_fetch0_fl_i_5
       (.I0(ctl_fetch0_fl_i_18_n_0),
        .I1(stat[1]),
        .I2(\fch/ir0 [0]),
        .I3(\ccmd[1]_INST_0_i_5_n_0 ),
        .I4(\bcmd[1]_INST_0_i_3_n_0 ),
        .I5(\ccmd[1]_INST_0_i_7_n_0 ),
        .O(ctl_fetch0_fl_i_5_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    ctl_fetch0_fl_i_50
       (.I0(div_crdy0),
        .I1(crdy),
        .I2(\fch/ir0 [7]),
        .O(ctl_fetch0_fl_i_50_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch0_fl_i_51
       (.I0(stat[2]),
        .I1(stat[1]),
        .O(ctl_fetch0_fl_i_51_n_0));
  LUT6 #(
    .INIT(64'h0000000022022232)) 
    ctl_fetch0_fl_i_6
       (.I0(ctl_fetch0_fl_i_19_n_0),
        .I1(ctl_fetch0_fl_i_20_n_0),
        .I2(\ccmd[0]_INST_0_i_13_n_0 ),
        .I3(ctl_fetch0_fl_i_21_n_0),
        .I4(ctl_fetch0_fl_i_22_n_0),
        .I5(ctl_fetch0_fl_i_23_n_0),
        .O(ctl_fetch0_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'h00000000EEEEEEE0)) 
    ctl_fetch0_fl_i_7
       (.I0(ctl_fetch0_fl_i_24_n_0),
        .I1(ctl_fetch0_fl_i_25_n_0),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir0 [14]),
        .I4(\ccmd[0]_INST_0_i_20_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(ctl_fetch0_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000000055DFDFDF)) 
    ctl_fetch0_fl_i_8
       (.I0(stat[0]),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [1]),
        .I4(stat[1]),
        .I5(ctl_fetch0_fl_i_26_n_0),
        .O(ctl_fetch0_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hF7F7FFF7F5F5FFF7)) 
    ctl_fetch0_fl_i_9
       (.I0(ctl_fetch0_fl_i_27_n_0),
        .I1(\rgf/sreg/sr [11]),
        .I2(\fch/ir0 [7]),
        .I3(\rgf/sreg/sr [8]),
        .I4(stat[0]),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(ctl_fetch0_fl_i_9_n_0));
  LUT6 #(
    .INIT(64'h00000000FEAAFEFE)) 
    ctl_fetch1_fl_i_1
       (.I0(ctl_fetch1_fl_reg_i_2_n_0),
        .I1(ctl_fetch1_fl_i_3_n_0),
        .I2(ctl_fetch1_fl_i_4_n_0),
        .I3(ctl_fetch1_fl_i_5_n_0),
        .I4(ctl_fetch1_fl_i_6_n_0),
        .I5(ctl_fetch1_fl_i_7_n_0),
        .O(ctl_fetch1));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFFBFFBB)) 
    ctl_fetch1_fl_i_10
       (.I0(ctl_fetch1_fl_i_26_n_0),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [1]),
        .O(ctl_fetch1_fl_i_10_n_0));
  LUT5 #(
    .INIT(32'h11111511)) 
    ctl_fetch1_fl_i_11
       (.I0(\bcmd[1]_INST_0_i_25_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [0]),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .O(ctl_fetch1_fl_i_11_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAA2A)) 
    ctl_fetch1_fl_i_12
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(ctl_fetch1_fl_i_16_n_0),
        .I2(ctl_fetch1_fl_i_27_n_0),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\fch/ir1 [15]),
        .O(ctl_fetch1_fl_i_12_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch1_fl_i_13
       (.I0(div_crdy1),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(ctl_fetch1_fl_i_13_n_0));
  LUT6 #(
    .INIT(64'h0000555500005100)) 
    ctl_fetch1_fl_i_14
       (.I0(ctl_fetch1_fl_i_28_n_0),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\rgf/sreg/sr [11]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [9]),
        .O(ctl_fetch1_fl_i_14_n_0));
  LUT6 #(
    .INIT(64'h7777777707775555)) 
    ctl_fetch1_fl_i_15
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\rgf/sreg/sr [11]),
        .I3(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(ctl_fetch1_fl_i_15_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_16
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .O(ctl_fetch1_fl_i_16_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFC5000000)) 
    ctl_fetch1_fl_i_17
       (.I0(ctl_fetch1_fl_i_29_n_0),
        .I1(ctl_fetch1_fl_i_30_n_0),
        .I2(ctl_fetch1_fl_i_31_n_0),
        .I3(ctl_fetch1_fl_i_32_n_0),
        .I4(ctl_fetch1_fl_i_33_n_0),
        .I5(ctl_fetch1_fl_i_34_n_0),
        .O(ctl_fetch1_fl_i_17_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_18
       (.I0(\fch/ir1 [6]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .O(ctl_fetch1_fl_i_18_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF55000075)) 
    ctl_fetch1_fl_i_19
       (.I0(\fch/ir1 [0]),
        .I1(fch_irq_req),
        .I2(irq),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [3]),
        .I5(ctl_fetch1_fl_i_35_n_0),
        .O(ctl_fetch1_fl_i_19_n_0));
  LUT6 #(
    .INIT(64'hFBFBBBFBFBFFBBFB)) 
    ctl_fetch1_fl_i_20
       (.I0(\stat[2]_i_5__0_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [14]),
        .I5(\rgf/sreg/sr [5]),
        .O(ctl_fetch1_fl_i_20_n_0));
  LUT6 #(
    .INIT(64'hAC00AC00AC000C00)) 
    ctl_fetch1_fl_i_21
       (.I0(ctl_fetch1_fl_i_36_n_0),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\badr[15]_INST_0_i_120_n_0 ),
        .O(ctl_fetch1_fl_i_21_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_22
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .O(ctl_fetch1_fl_i_22_n_0));
  LUT6 #(
    .INIT(64'hFEFEFEFEFEFFFEFE)) 
    ctl_fetch1_fl_i_23
       (.I0(ctl_fetch1_fl_i_37_n_0),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\rgf/sreg/sr [5]),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [12]),
        .O(ctl_fetch1_fl_i_23_n_0));
  LUT6 #(
    .INIT(64'h0045004500000045)) 
    ctl_fetch1_fl_i_24
       (.I0(ctl_fetch1_fl_i_38_n_0),
        .I1(\badr[15]_INST_0_i_120_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I3(ctl_fetch1_fl_i_39_n_0),
        .I4(\bdatw[31]_INST_0_i_151_n_0 ),
        .I5(ctl_fetch1_fl_i_40_n_0),
        .O(ctl_fetch1_fl_i_24_n_0));
  LUT6 #(
    .INIT(64'h003050300F3F5030)) 
    ctl_fetch1_fl_i_25
       (.I0(\stat[1]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [13]),
        .I5(\rgf/sreg/sr [6]),
        .O(ctl_fetch1_fl_i_25_n_0));
  LUT6 #(
    .INIT(64'hAFFFFFFCAFFFAFFC)) 
    ctl_fetch1_fl_i_26
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [7]),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(ctl_fetch1_fl_i_26_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_fetch1_fl_i_27
       (.I0(\fch/ir1 [10]),
        .I1(div_crdy1),
        .O(ctl_fetch1_fl_i_27_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_fetch1_fl_i_28
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [10]),
        .O(ctl_fetch1_fl_i_28_n_0));
  LUT6 #(
    .INIT(64'hA700A700FFFFA700)) 
    ctl_fetch1_fl_i_29
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [9]),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(ctl_fetch1_fl_i_41_n_0),
        .O(ctl_fetch1_fl_i_29_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4440000)) 
    ctl_fetch1_fl_i_3
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [1]),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(ctl_fetch1_fl_i_10_n_0),
        .O(ctl_fetch1_fl_i_3_n_0));
  LUT3 #(
    .INIT(8'hB4)) 
    ctl_fetch1_fl_i_30
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .O(ctl_fetch1_fl_i_30_n_0));
  LUT4 #(
    .INIT(16'h8000)) 
    ctl_fetch1_fl_i_31
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .O(ctl_fetch1_fl_i_31_n_0));
  LUT5 #(
    .INIT(32'h00000080)) 
    ctl_fetch1_fl_i_32
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat_reg_n_0_[2] ),
        .I4(\fch/ir1 [15]),
        .O(ctl_fetch1_fl_i_32_n_0));
  LUT6 #(
    .INIT(64'h5400FCCC0000CCCC)) 
    ctl_fetch1_fl_i_33
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [7]),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\rgf_selc1_wb[1]_i_31_n_0 ),
        .O(ctl_fetch1_fl_i_33_n_0));
  LUT6 #(
    .INIT(64'h00000000000001CD)) 
    ctl_fetch1_fl_i_34
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(ctl_fetch1_fl_i_42_n_0),
        .I5(\bcmd[3]_INST_0_i_4_n_0 ),
        .O(ctl_fetch1_fl_i_34_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFFFFF)) 
    ctl_fetch1_fl_i_35
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [10]),
        .I2(\bdatw[31]_INST_0_i_173_n_0 ),
        .I3(\fch/ir1 [2]),
        .I4(ctl_fetch1_fl_i_43_n_0),
        .I5(\bcmd[3]_INST_0_i_22_n_0 ),
        .O(ctl_fetch1_fl_i_35_n_0));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEEE0000)) 
    ctl_fetch1_fl_i_36
       (.I0(ctl_fetch1_fl_i_44_n_0),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(div_crdy1),
        .O(ctl_fetch1_fl_i_36_n_0));
  LUT6 #(
    .INIT(64'h8A8AAAAA8A8A8AAA)) 
    ctl_fetch1_fl_i_37
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(ctl_fetch1_fl_i_45_n_0),
        .I2(ctl_fetch1_fl_i_46_n_0),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [6]),
        .O(ctl_fetch1_fl_i_37_n_0));
  LUT6 #(
    .INIT(64'hFF3F5F5F7F3F5F5F)) 
    ctl_fetch1_fl_i_38
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(ctl_fetch1_fl_i_47_n_0),
        .O(ctl_fetch1_fl_i_38_n_0));
  LUT6 #(
    .INIT(64'h0000000001F1FFFF)) 
    ctl_fetch1_fl_i_39
       (.I0(\rgf/sreg/sr [11]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [8]),
        .I5(ctl_fetch1_fl_i_28_n_0),
        .O(ctl_fetch1_fl_i_39_n_0));
  LUT6 #(
    .INIT(64'h8BB8888BBBBBBBBB)) 
    ctl_fetch1_fl_i_4
       (.I0(\bcmd[1]_INST_0_i_11_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [3]),
        .I5(ctl_fetch1_fl_i_11_n_0),
        .O(ctl_fetch1_fl_i_4_n_0));
  LUT3 #(
    .INIT(8'hC9)) 
    ctl_fetch1_fl_i_40
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [5]),
        .O(ctl_fetch1_fl_i_40_n_0));
  LUT3 #(
    .INIT(8'h65)) 
    ctl_fetch1_fl_i_41
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .O(ctl_fetch1_fl_i_41_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    ctl_fetch1_fl_i_42
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [2]),
        .I4(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(ctl_fetch1_fl_i_42_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    ctl_fetch1_fl_i_43
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .O(ctl_fetch1_fl_i_43_n_0));
  LUT6 #(
    .INIT(64'h00D0000000000000)) 
    ctl_fetch1_fl_i_44
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\rgf/sreg/sr [10]),
        .I2(div_crdy1),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(ctl_fetch1_fl_i_44_n_0));
  LUT6 #(
    .INIT(64'hF0400040F040F040)) 
    ctl_fetch1_fl_i_45
       (.I0(\rgf/sreg/sr [10]),
        .I1(ctl_fetch1_fl_i_48_n_0),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\bdatw[31]_INST_0_i_139_n_0 ),
        .I5(\fch/ir1 [10]),
        .O(ctl_fetch1_fl_i_45_n_0));
  LUT6 #(
    .INIT(64'h7F776E66FFFFFFFF)) 
    ctl_fetch1_fl_i_46
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\rgf/sreg/sr [11]),
        .I5(\fch/ir1 [8]),
        .O(ctl_fetch1_fl_i_46_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch1_fl_i_47
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [5]),
        .O(ctl_fetch1_fl_i_47_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    ctl_fetch1_fl_i_48
       (.I0(div_crdy1),
        .I1(\fch/ir1 [7]),
        .O(ctl_fetch1_fl_i_48_n_0));
  LUT6 #(
    .INIT(64'hEAEEEEEEFFEEEEEE)) 
    ctl_fetch1_fl_i_5
       (.I0(ctl_fetch1_fl_i_12_n_0),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(div_crdy1),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [12]),
        .O(ctl_fetch1_fl_i_5_n_0));
  LUT6 #(
    .INIT(64'hAABFAAAABFBFBFBF)) 
    ctl_fetch1_fl_i_6
       (.I0(ctl_fetch1_fl_i_13_n_0),
        .I1(\bcmd[1]_INST_0_i_15_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(ctl_fetch1_fl_i_14_n_0),
        .I4(ctl_fetch1_fl_i_15_n_0),
        .I5(ctl_fetch1_fl_i_16_n_0),
        .O(ctl_fetch1_fl_i_6_n_0));
  LUT6 #(
    .INIT(64'h000000008AAA8888)) 
    ctl_fetch1_fl_i_7
       (.I0(ctl_fetch1_fl_i_17_n_0),
        .I1(\fch/ir1 [3]),
        .I2(ctl_fetch1_fl_i_18_n_0),
        .I3(\fch/ir1 [8]),
        .I4(\bcmd[3]_INST_0_i_13_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(ctl_fetch1_fl_i_7_n_0));
  LUT6 #(
    .INIT(64'hF2F200F2F2F2F2F2)) 
    ctl_fetch1_fl_i_8
       (.I0(ctl_fetch1_fl_i_19_n_0),
        .I1(ctl_fetch1_fl_i_20_n_0),
        .I2(ctl_fetch1_fl_i_21_n_0),
        .I3(\fch/ir1 [12]),
        .I4(\rgf/sreg/sr [7]),
        .I5(ctl_fetch1_fl_i_22_n_0),
        .O(ctl_fetch1_fl_i_8_n_0));
  LUT6 #(
    .INIT(64'hFFABFFABFAAAFFAB)) 
    ctl_fetch1_fl_i_9
       (.I0(ctl_fetch1_fl_i_23_n_0),
        .I1(ctl_fetch1_fl_i_24_n_0),
        .I2(\rgf_selc1_wb[1]_i_38_n_0 ),
        .I3(ctl_fetch1_fl_i_25_n_0),
        .I4(\rgf/sreg/sr [7]),
        .I5(\fch/ir1 [14]),
        .O(ctl_fetch1_fl_i_9_n_0));
  MUXF7 ctl_fetch1_fl_reg_i_2
       (.I0(ctl_fetch1_fl_i_8_n_0),
        .I1(ctl_fetch1_fl_i_9_n_0),
        .O(ctl_fetch1_fl_reg_i_2_n_0),
        .S(\fch/ir1 [11]));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_ext_fl_i_1
       (.I0(\nir_id[24]_i_6_n_0 ),
        .O(\fch/ctl_fetch_ext ));
  LUT1 #(
    .INIT(2'h1)) 
    ctl_fetch_lng_fl_i_1
       (.I0(fch_heir_nir_i_3_n_0),
        .O(\fch/ctl_fetch_lng ));
  LUT3 #(
    .INIT(8'hB8)) 
    dctl_long_f_i_1
       (.I0(\rgf/sreg/sr [8]),
        .I1(div_crdy0),
        .I2(\alu0/div/dctl/dctl_long_f ),
        .O(\alu0/div/dctl_long ));
  LUT3 #(
    .INIT(8'hB8)) 
    dctl_long_f_i_1__0
       (.I0(\rgf/sreg/sr [8]),
        .I1(div_crdy1),
        .I2(\alu1/div/dctl/dctl_long_f ),
        .O(\alu1/div/dctl_long ));
  LUT6 #(
    .INIT(64'h8000FFFF80000000)) 
    dctl_sign_f_i_1
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I4(div_crdy0),
        .I5(\alu0/div/dctl/dctl_sign_f ),
        .O(\alu0/div/dctl/dctl_sign ));
  LUT6 #(
    .INIT(64'hBABABBBABABBBABA)) 
    dctl_sign_f_i_10
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(dctl_sign_f_i_13_n_0),
        .I2(dctl_sign_f_i_14_n_0),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [14]),
        .O(dctl_sign_f_i_10_n_0));
  LUT3 #(
    .INIT(8'hE7)) 
    dctl_sign_f_i_11
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [3]),
        .O(dctl_sign_f_i_11_n_0));
  LUT6 #(
    .INIT(64'h0001020003080200)) 
    dctl_sign_f_i_12
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [5]),
        .I2(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [3]),
        .O(dctl_sign_f_i_12_n_0));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    dctl_sign_f_i_13
       (.I0(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [3]),
        .I4(\bdatw[31]_INST_0_i_173_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .O(dctl_sign_f_i_13_n_0));
  LUT6 #(
    .INIT(64'hFEEEEEEEFFFFFFFF)) 
    dctl_sign_f_i_14
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [15]),
        .O(dctl_sign_f_i_14_n_0));
  LUT6 #(
    .INIT(64'h8000FFFF80000000)) 
    dctl_sign_f_i_1__0
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(acmd1[0]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(div_crdy1),
        .I5(\alu1/div/dctl/dctl_sign_f ),
        .O(\alu1/div/dctl/dctl_sign ));
  LUT6 #(
    .INIT(64'h1010101155555555)) 
    dctl_sign_f_i_2
       (.I0(\niss_dsp_a1[32]_INST_0_i_9_n_0 ),
        .I1(\bcmd[2]_INST_0_i_1_n_0 ),
        .I2(dctl_sign_f_i_3_n_0),
        .I3(dctl_sign_f_i_4_n_0),
        .I4(dctl_sign_f_i_5_n_0),
        .I5(dctl_sign_f_i_6_n_0),
        .O(dctl_sign_f_i_2_n_0));
  LUT6 #(
    .INIT(64'hCCCDCCCDCCCDCFCD)) 
    dctl_sign_f_i_3
       (.I0(dctl_sign_f_i_7_n_0),
        .I1(dctl_sign_f_i_8_n_0),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [6]),
        .I4(dctl_sign_f_i_9_n_0),
        .I5(\fch/ir1 [7]),
        .O(dctl_sign_f_i_3_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    dctl_sign_f_i_4
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .O(dctl_sign_f_i_4_n_0));
  LUT6 #(
    .INIT(64'hBF53BF73AAFABFFB)) 
    dctl_sign_f_i_5
       (.I0(\fch/ir1 [6]),
        .I1(div_crdy1),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [11]),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(\fch/ir1 [7]),
        .O(dctl_sign_f_i_5_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAA8AAAAAAAA)) 
    dctl_sign_f_i_6
       (.I0(dctl_sign_f_i_10_n_0),
        .I1(\rgf_selc1_rn_wb[1]_i_19_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_14_n_0 ),
        .I4(dctl_sign_f_i_11_n_0),
        .I5(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .O(dctl_sign_f_i_6_n_0));
  LUT6 #(
    .INIT(64'hFF00FF00FBBBFFFF)) 
    dctl_sign_f_i_7
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(div_crdy1),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [11]),
        .O(dctl_sign_f_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFB0000000)) 
    dctl_sign_f_i_8
       (.I0(div_crdy1),
        .I1(\fch/ir1 [10]),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_24_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(dctl_sign_f_i_12_n_0),
        .O(dctl_sign_f_i_8_n_0));
  LUT4 #(
    .INIT(16'hFBBB)) 
    dctl_sign_f_i_9
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(div_crdy1),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [8]),
        .O(dctl_sign_f_i_9_n_0));
  LUT6 #(
    .INIT(64'h4F4F5F5F404F5050)) 
    \dctl_stat[0]_i_1 
       (.I0(\alu0/div/dctl_stat [0]),
        .I1(\dctl_stat[1]_i_3_n_0 ),
        .I2(\alu0/div/dctl_stat [1]),
        .I3(\alu0/div/dctl_stat [2]),
        .I4(\alu0/div/dctl_stat [3]),
        .I5(\dctl_stat[0]_i_2_n_0 ),
        .O(\alu0/div/dctl/fsm/dctl_next [0]));
  LUT5 #(
    .INIT(32'h45FF4500)) 
    \dctl_stat[0]_i_1__0 
       (.I0(\alu1/div/dctl_stat [0]),
        .I1(\dctl_stat[1]_i_3__0_n_0 ),
        .I2(\alu1/div/dctl_stat [3]),
        .I3(\alu1/div/dctl_stat [1]),
        .I4(\dctl_stat[0]_i_2__0_n_0 ),
        .O(\alu1/div/dctl/fsm/dctl_next [0]));
  LUT6 #(
    .INIT(64'h007F007F0000007F)) 
    \dctl_stat[0]_i_2 
       (.I0(\alu0/div/den2 ),
        .I1(\alu0/div/dctl/dctl_sign ),
        .I2(\alu0/div/dctl_stat [0]),
        .I3(\dctl_stat[0]_i_3_n_0 ),
        .I4(\dctl_stat[2]_i_2_n_0 ),
        .I5(\alu0/div/dctl_stat [2]),
        .O(\dctl_stat[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h222222EF22EF22EF)) 
    \dctl_stat[0]_i_2__0 
       (.I0(\alu1/div/dctl_stat [3]),
        .I1(\alu1/div/dctl_stat [2]),
        .I2(\dctl_stat[2]_i_2__0_n_0 ),
        .I3(\dctl_stat[0]_i_3__0_n_0 ),
        .I4(\alu1/div/dctl_stat [0]),
        .I5(\alu1/div/dctl/fsm/chg_rem_sgn0 ),
        .O(\dctl_stat[0]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h00FFD700)) 
    \dctl_stat[0]_i_3 
       (.I0(\alu0/div/chg_rem_sgn ),
        .I1(\alu0/div/chg_quo_sgn ),
        .I2(\alu0/div/fdiv_rem_msb_f ),
        .I3(\alu0/div/dctl_stat [3]),
        .I4(\alu0/div/dctl_stat [0]),
        .O(\dctl_stat[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00FFD700)) 
    \dctl_stat[0]_i_3__0 
       (.I0(\alu1/div/chg_rem_sgn ),
        .I1(\alu1/div/chg_quo_sgn ),
        .I2(\alu1/div/fdiv_rem_msb_f ),
        .I3(\alu1/div/dctl_stat [3]),
        .I4(\alu1/div/dctl_stat [0]),
        .O(\dctl_stat[0]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h0F300B38)) 
    \dctl_stat[1]_i_1 
       (.I0(\dctl_stat[1]_i_2_n_0 ),
        .I1(\alu0/div/dctl_stat [3]),
        .I2(\alu0/div/dctl_stat [0]),
        .I3(\alu0/div/dctl_stat [1]),
        .I4(\dctl_stat[1]_i_3_n_0 ),
        .O(\alu0/div/dctl/fsm/dctl_next [1]));
  LUT5 #(
    .INIT(32'h0F300B38)) 
    \dctl_stat[1]_i_1__0 
       (.I0(\dctl_stat[1]_i_2__0_n_0 ),
        .I1(\alu1/div/dctl_stat [3]),
        .I2(\alu1/div/dctl_stat [0]),
        .I3(\alu1/div/dctl_stat [1]),
        .I4(\dctl_stat[1]_i_3__0_n_0 ),
        .O(\alu1/div/dctl/fsm/dctl_next [1]));
  LUT5 #(
    .INIT(32'h0C080800)) 
    \dctl_stat[1]_i_2 
       (.I0(\alu0/div/fdiv_rem_msb_f ),
        .I1(\alu0/div/dctl_stat [2]),
        .I2(\alu0/div/dctl_stat [1]),
        .I3(\alu0/div/chg_quo_sgn ),
        .I4(\alu0/div/chg_rem_sgn ),
        .O(\dctl_stat[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h0C080800)) 
    \dctl_stat[1]_i_2__0 
       (.I0(\alu1/div/fdiv_rem_msb_f ),
        .I1(\alu1/div/dctl_stat [2]),
        .I2(\alu1/div/dctl_stat [1]),
        .I3(\alu1/div/chg_quo_sgn ),
        .I4(\alu1/div/chg_rem_sgn ),
        .O(\dctl_stat[1]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \dctl_stat[1]_i_3 
       (.I0(\alu0/div/chg_rem_sgn ),
        .I1(\alu0/div/chg_quo_sgn ),
        .I2(\alu0/div/dctl_stat [2]),
        .O(\dctl_stat[1]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \dctl_stat[1]_i_3__0 
       (.I0(\alu1/div/chg_rem_sgn ),
        .I1(\alu1/div/chg_quo_sgn ),
        .I2(\alu1/div/dctl_stat [2]),
        .O(\dctl_stat[1]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFC1)) 
    \dctl_stat[2]_i_1 
       (.I0(\dctl_stat[2]_i_2_n_0 ),
        .I1(\alu0/div/dctl_stat [0]),
        .I2(\alu0/div/dctl_stat [1]),
        .I3(\alu0/div/dctl_stat [2]),
        .I4(\alu0/div/dctl_stat [3]),
        .O(\alu0/div/dctl/fsm/dctl_next [2]));
  LUT5 #(
    .INIT(32'h0000FFC1)) 
    \dctl_stat[2]_i_1__0 
       (.I0(\dctl_stat[2]_i_2__0_n_0 ),
        .I1(\alu1/div/dctl_stat [0]),
        .I2(\alu1/div/dctl_stat [1]),
        .I3(\alu1/div/dctl_stat [2]),
        .I4(\alu1/div/dctl_stat [3]),
        .O(\alu1/div/dctl/fsm/dctl_next [2]));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \dctl_stat[2]_i_2 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\dctl_stat[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \dctl_stat[2]_i_2__0 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(acmd1[4]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .O(\dctl_stat[2]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4FFF4F4)) 
    \dctl_stat[3]_i_1 
       (.I0(\dctl_stat[3]_i_2_n_0 ),
        .I1(\alu0/div/dctl/fsm/set_sgn ),
        .I2(\dctl_stat[3]_i_4_n_0 ),
        .I3(\alu0/div/dctl_stat [0]),
        .I4(\alu0/div/dctl_stat [3]),
        .I5(\dctl_stat[3]_i_5_n_0 ),
        .O(\alu0/div/dctl/fsm/dctl_next [3]));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4FFF4F4)) 
    \dctl_stat[3]_i_1__0 
       (.I0(\dctl_stat[3]_i_2__0_n_0 ),
        .I1(\alu1/div/dctl/fsm/set_sgn ),
        .I2(\dctl_stat[3]_i_4__0_n_0 ),
        .I3(\alu1/div/dctl_stat [0]),
        .I4(\alu1/div/dctl_stat [3]),
        .I5(\dctl_stat[3]_i_5__0_n_0 ),
        .O(\alu1/div/dctl/fsm/dctl_next [3]));
  LUT3 #(
    .INIT(8'h4F)) 
    \dctl_stat[3]_i_2 
       (.I0(\alu0/div/den2 ),
        .I1(chg_quo_sgn_i_2_n_0),
        .I2(\alu0/div/dctl/dctl_sign ),
        .O(\dctl_stat[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \dctl_stat[3]_i_2__0 
       (.I0(\alu1/div/den2 ),
        .I1(chg_quo_sgn_i_2__0_n_0),
        .I2(\alu1/div/dctl/dctl_sign ),
        .O(\dctl_stat[3]_i_2__0_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \dctl_stat[3]_i_3 
       (.I0(\alu0/div/dctl_stat [1]),
        .I1(\alu0/div/dctl_stat [2]),
        .I2(\alu0/div/dctl_stat [0]),
        .I3(\alu0/div/dctl_stat [3]),
        .O(\alu0/div/dctl/fsm/set_sgn ));
  LUT4 #(
    .INIT(16'h4000)) 
    \dctl_stat[3]_i_3__0 
       (.I0(\alu1/div/dctl_stat [1]),
        .I1(\alu1/div/dctl_stat [2]),
        .I2(\alu1/div/dctl_stat [0]),
        .I3(\alu1/div/dctl_stat [3]),
        .O(\alu1/div/dctl/fsm/set_sgn ));
  LUT6 #(
    .INIT(64'h00000000F5000003)) 
    \dctl_stat[3]_i_4 
       (.I0(\alu0/div/dctl_long ),
        .I1(\dctl_stat[2]_i_2_n_0 ),
        .I2(\alu0/div/dctl_stat [2]),
        .I3(\alu0/div/dctl_stat [1]),
        .I4(\alu0/div/dctl_stat [0]),
        .I5(\alu0/div/dctl_stat [3]),
        .O(\dctl_stat[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F5000003)) 
    \dctl_stat[3]_i_4__0 
       (.I0(\alu1/div/dctl_long ),
        .I1(\dctl_stat[2]_i_2__0_n_0 ),
        .I2(\alu1/div/dctl_stat [2]),
        .I3(\alu1/div/dctl_stat [1]),
        .I4(\alu1/div/dctl_stat [0]),
        .I5(\alu1/div/dctl_stat [3]),
        .O(\dctl_stat[3]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hF00AFF3AFF3AFFFA)) 
    \dctl_stat[3]_i_5 
       (.I0(chg_quo_sgn_i_2_n_0),
        .I1(\alu0/div/fdiv_rem_msb_f ),
        .I2(\alu0/div/dctl_stat [2]),
        .I3(\alu0/div/dctl_stat [1]),
        .I4(\alu0/div/chg_quo_sgn ),
        .I5(\alu0/div/chg_rem_sgn ),
        .O(\dctl_stat[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF00AFF3AFF3AFFFA)) 
    \dctl_stat[3]_i_5__0 
       (.I0(chg_quo_sgn_i_2__0_n_0),
        .I1(\alu1/div/fdiv_rem_msb_f ),
        .I2(\alu1/div/dctl_stat [2]),
        .I3(\alu1/div/dctl_stat [1]),
        .I4(\alu1/div/chg_quo_sgn ),
        .I5(\alu1/div/chg_rem_sgn ),
        .O(\dctl_stat[3]_i_5__0_n_0 ));
  LUT3 #(
    .INIT(8'hC8)) 
    div_crdy_i_1
       (.I0(div_crdy_i_2_n_0),
        .I1(\dctl_stat[2]_i_2_n_0 ),
        .I2(div_crdy0),
        .O(div_crdy_i_1_n_0));
  LUT3 #(
    .INIT(8'hC8)) 
    div_crdy_i_1__0
       (.I0(div_crdy_i_2__0_n_0),
        .I1(\dctl_stat[2]_i_2__0_n_0 ),
        .I2(div_crdy1),
        .O(div_crdy_i_1__0_n_0));
  LUT5 #(
    .INIT(32'hFFFF5700)) 
    div_crdy_i_2
       (.I0(\alu0/div/dctl/dctl_sign ),
        .I1(\alu0/div/chg_rem_sgn ),
        .I2(\alu0/div/chg_quo_sgn ),
        .I3(div_crdy_i_3_n_0),
        .I4(div_crdy_i_4_n_0),
        .O(div_crdy_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFF5700)) 
    div_crdy_i_2__0
       (.I0(\alu1/div/dctl/dctl_sign ),
        .I1(\alu1/div/chg_rem_sgn ),
        .I2(\alu1/div/chg_quo_sgn ),
        .I3(div_crdy_i_3__0_n_0),
        .I4(div_crdy_i_4__0_n_0),
        .O(div_crdy_i_2__0_n_0));
  LUT5 #(
    .INIT(32'h08000808)) 
    div_crdy_i_3
       (.I0(\alu0/div/dctl_stat [1]),
        .I1(\alu0/div/dctl_stat [0]),
        .I2(\alu0/div/dctl_stat [3]),
        .I3(\alu0/div/dctl_stat [2]),
        .I4(\alu0/div/dctl_long ),
        .O(div_crdy_i_3_n_0));
  LUT5 #(
    .INIT(32'h08000808)) 
    div_crdy_i_3__0
       (.I0(\alu1/div/dctl_stat [1]),
        .I1(\alu1/div/dctl_stat [0]),
        .I2(\alu1/div/dctl_stat [3]),
        .I3(\alu1/div/dctl_stat [2]),
        .I4(\alu1/div/dctl_long ),
        .O(div_crdy_i_3__0_n_0));
  LUT6 #(
    .INIT(64'h000000F000700000)) 
    div_crdy_i_4
       (.I0(\alu0/div/fdiv_rem_msb_f ),
        .I1(\alu0/div/chg_quo_sgn ),
        .I2(\alu0/div/dctl_stat [3]),
        .I3(\alu0/div/dctl_stat [0]),
        .I4(\alu0/div/dctl_stat [2]),
        .I5(\alu0/div/dctl_stat [1]),
        .O(div_crdy_i_4_n_0));
  LUT6 #(
    .INIT(64'h000000F000700000)) 
    div_crdy_i_4__0
       (.I0(\alu1/div/fdiv_rem_msb_f ),
        .I1(\alu1/div/chg_quo_sgn ),
        .I2(\alu1/div/dctl_stat [3]),
        .I3(\alu1/div/dctl_stat [0]),
        .I4(\alu1/div/dctl_stat [2]),
        .I5(\alu1/div/dctl_stat [1]),
        .O(div_crdy_i_4__0_n_0));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [11]),
        .O(\dso[11]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [11]),
        .O(\dso[11]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [10]),
        .O(\dso[11]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [10]),
        .O(\dso[11]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [9]),
        .O(\dso[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [9]),
        .O(\dso[11]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [8]),
        .O(\dso[11]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[11]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [8]),
        .O(\dso[11]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_2 
       (.I0(\alu0/div/p_0_out [11]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_2__0 
       (.I0(\alu1/div/p_0_out [11]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_3 
       (.I0(\alu0/div/p_0_out [10]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_3__0 
       (.I0(\alu1/div/p_0_out [10]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_4 
       (.I0(\alu0/div/p_0_out [9]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_4__0 
       (.I0(\alu1/div/p_0_out [9]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_5 
       (.I0(\alu0/div/p_0_out [8]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_5__0 
       (.I0(\alu1/div/p_0_out [8]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[11]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_6 
       (.I0(\alu0/div/p_0_out [11]),
        .I1(\dso[11]_i_10_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [11]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[11]),
        .O(\dso[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_6__0 
       (.I0(\alu1/div/p_0_out [11]),
        .I1(\dso[11]_i_10__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [11]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[11]),
        .O(\dso[11]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_7 
       (.I0(\alu0/div/p_0_out [10]),
        .I1(\dso[11]_i_11_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [10]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[10]),
        .O(\dso[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_7__0 
       (.I0(\alu1/div/p_0_out [10]),
        .I1(\dso[11]_i_11__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [10]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[10]),
        .O(\dso[11]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_8 
       (.I0(\alu0/div/p_0_out [9]),
        .I1(\dso[11]_i_12_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [9]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[9]),
        .O(\dso[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_8__0 
       (.I0(\alu1/div/p_0_out [9]),
        .I1(\dso[11]_i_12__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [9]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[9]),
        .O(\dso[11]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_9 
       (.I0(\alu0/div/p_0_out [8]),
        .I1(\dso[11]_i_13_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [8]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[8]),
        .O(\dso[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_9__0 
       (.I0(\alu1/div/p_0_out [8]),
        .I1(\dso[11]_i_13__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [8]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[8]),
        .O(\dso[11]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [15]),
        .O(\dso[15]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [15]),
        .O(\dso[15]_i_10__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \dso[15]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/dctl/dctl_long_f ),
        .I3(div_crdy0),
        .I4(\rgf/sreg/sr [8]),
        .O(\dso[15]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \dso[15]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/dctl/dctl_long_f ),
        .I3(div_crdy1),
        .I4(\rgf/sreg/sr [8]),
        .O(\dso[15]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [14]),
        .O(\dso[15]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [14]),
        .O(\dso[15]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [13]),
        .O(\dso[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [13]),
        .O(\dso[15]_i_13__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_14 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [12]),
        .O(\dso[15]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[15]_i_14__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [12]),
        .O(\dso[15]_i_14__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_2 
       (.I0(\alu0/div/p_0_out [15]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_2__0 
       (.I0(\alu1/div/p_0_out [15]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_3 
       (.I0(\alu0/div/p_0_out [14]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_3__0 
       (.I0(\alu1/div/p_0_out [14]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_4 
       (.I0(\alu0/div/p_0_out [13]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_4__0 
       (.I0(\alu1/div/p_0_out [13]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_5 
       (.I0(\alu0/div/p_0_out [12]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_5__0 
       (.I0(\alu1/div/p_0_out [12]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_6 
       (.I0(\alu0/div/p_0_out [15]),
        .I1(\dso[15]_i_10_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [15]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[15]),
        .O(\dso[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_6__0 
       (.I0(\alu1/div/p_0_out [15]),
        .I1(\dso[15]_i_10__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [15]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[15]),
        .O(\dso[15]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_7 
       (.I0(\alu0/div/p_0_out [14]),
        .I1(\dso[15]_i_12_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [14]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[14]),
        .O(\dso[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_7__0 
       (.I0(\alu1/div/p_0_out [14]),
        .I1(\dso[15]_i_12__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [14]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[14]),
        .O(\dso[15]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_8 
       (.I0(\alu0/div/p_0_out [13]),
        .I1(\dso[15]_i_13_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [13]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[13]),
        .O(\dso[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_8__0 
       (.I0(\alu1/div/p_0_out [13]),
        .I1(\dso[15]_i_13__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [13]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[13]),
        .O(\dso[15]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_9 
       (.I0(\alu0/div/p_0_out [12]),
        .I1(\dso[15]_i_14_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [12]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[12]),
        .O(\dso[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_9__0 
       (.I0(\alu1/div/p_0_out [12]),
        .I1(\dso[15]_i_14__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [12]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[12]),
        .O(\dso[15]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [19]),
        .O(\dso[19]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [19]),
        .O(\dso[19]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [18]),
        .O(\dso[19]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [18]),
        .O(\dso[19]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [17]),
        .O(\dso[19]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [17]),
        .O(\dso[19]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [16]),
        .O(\dso[19]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[19]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [16]),
        .O(\dso[19]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_2 
       (.I0(\alu0/div/p_0_out [19]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_2__0 
       (.I0(\alu1/div/p_0_out [19]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_3 
       (.I0(\alu0/div/p_0_out [18]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_3__0 
       (.I0(\alu1/div/p_0_out [18]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_4 
       (.I0(\alu0/div/p_0_out [17]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_4__0 
       (.I0(\alu1/div/p_0_out [17]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_5 
       (.I0(\alu0/div/p_0_out [16]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[19]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_5__0 
       (.I0(\alu1/div/p_0_out [16]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[19]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_6 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [19]),
        .I3(\dso[19]_i_10_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[19]),
        .O(\dso[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_6__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [19]),
        .I3(\dso[19]_i_10__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[19]),
        .O(\dso[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_7 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [18]),
        .I3(\dso[19]_i_11_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[18]),
        .O(\dso[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_7__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [18]),
        .I3(\dso[19]_i_11__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[18]),
        .O(\dso[19]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_8 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [17]),
        .I3(\dso[19]_i_12_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[17]),
        .O(\dso[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_8__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [17]),
        .I3(\dso[19]_i_12__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[17]),
        .O(\dso[19]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_9 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [16]),
        .I3(\dso[19]_i_13_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[16]),
        .O(\dso[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[19]_i_9__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [16]),
        .I3(\dso[19]_i_13__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[16]),
        .O(\dso[19]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [23]),
        .O(\dso[23]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [23]),
        .O(\dso[23]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [22]),
        .O(\dso[23]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [22]),
        .O(\dso[23]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [21]),
        .O(\dso[23]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [21]),
        .O(\dso[23]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [20]),
        .O(\dso[23]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[23]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [20]),
        .O(\dso[23]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_2 
       (.I0(\alu0/div/p_0_out [23]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_2__0 
       (.I0(\alu1/div/p_0_out [23]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_3 
       (.I0(\alu0/div/p_0_out [22]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_3__0 
       (.I0(\alu1/div/p_0_out [22]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_4 
       (.I0(\alu0/div/p_0_out [21]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_4__0 
       (.I0(\alu1/div/p_0_out [21]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_5 
       (.I0(\alu0/div/p_0_out [20]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[23]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_5__0 
       (.I0(\alu1/div/p_0_out [20]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[23]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_6 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [23]),
        .I3(\dso[23]_i_10_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[23]),
        .O(\dso[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_6__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [23]),
        .I3(\dso[23]_i_10__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[23]),
        .O(\dso[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_7 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [22]),
        .I3(\dso[23]_i_11_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[22]),
        .O(\dso[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_7__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [22]),
        .I3(\dso[23]_i_11__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[22]),
        .O(\dso[23]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_8 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [21]),
        .I3(\dso[23]_i_12_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[21]),
        .O(\dso[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_8__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [21]),
        .I3(\dso[23]_i_12__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[21]),
        .O(\dso[23]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_9 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [20]),
        .I3(\dso[23]_i_13_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[20]),
        .O(\dso[23]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[23]_i_9__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [20]),
        .I3(\dso[23]_i_13__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[20]),
        .O(\dso[23]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [27]),
        .O(\dso[27]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [27]),
        .O(\dso[27]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [26]),
        .O(\dso[27]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [26]),
        .O(\dso[27]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [25]),
        .O(\dso[27]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [25]),
        .O(\dso[27]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [24]),
        .O(\dso[27]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[27]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [24]),
        .O(\dso[27]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_2 
       (.I0(\alu0/div/p_0_out [27]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_2__0 
       (.I0(\alu1/div/p_0_out [27]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_3 
       (.I0(\alu0/div/p_0_out [26]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_3__0 
       (.I0(\alu1/div/p_0_out [26]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_4 
       (.I0(\alu0/div/p_0_out [25]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_4__0 
       (.I0(\alu1/div/p_0_out [25]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_5 
       (.I0(\alu0/div/p_0_out [24]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[27]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_5__0 
       (.I0(\alu1/div/p_0_out [24]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[27]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_6 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [27]),
        .I3(\dso[27]_i_10_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[27]),
        .O(\dso[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_6__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [27]),
        .I3(\dso[27]_i_10__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[27]),
        .O(\dso[27]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_7 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [26]),
        .I3(\dso[27]_i_11_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[26]),
        .O(\dso[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_7__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [26]),
        .I3(\dso[27]_i_11__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[26]),
        .O(\dso[27]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_8 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [25]),
        .I3(\dso[27]_i_12_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[25]),
        .O(\dso[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_8__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [25]),
        .I3(\dso[27]_i_12__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[25]),
        .O(\dso[27]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_9 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [24]),
        .I3(\dso[27]_i_13_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[24]),
        .O(\dso[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[27]_i_9__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [24]),
        .I3(\dso[27]_i_13__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[24]),
        .O(\dso[27]_i_9__0_n_0 ));
  LUT3 #(
    .INIT(8'hF1)) 
    \dso[31]_i_1 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\dso[31]_i_5_n_0 ),
        .O(\dso[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_10 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [30]),
        .I3(\dso[31]_i_18_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[30]),
        .O(\dso[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_10__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [30]),
        .I3(\dso[31]_i_18__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[30]),
        .O(\dso[31]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_11 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [29]),
        .I3(\dso[31]_i_19_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[29]),
        .O(\dso[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_11__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [29]),
        .I3(\dso[31]_i_19__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[29]),
        .O(\dso[31]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_12 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [28]),
        .I3(\dso[31]_i_20_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[28]),
        .O(\dso[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_12__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [28]),
        .I3(\dso[31]_i_20__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[28]),
        .O(\dso[31]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF7070F0FF707F)) 
    \dso[31]_i_13 
       (.I0(\alu0/div/dctl/dctl_sign ),
        .I1(\alu0/div/den2 ),
        .I2(\alu0/div/dctl_stat [0]),
        .I3(\alu0/div/chg_quo_sgn ),
        .I4(\alu0/div/dctl_stat [1]),
        .I5(\alu0/div/fdiv_rem_msb_f ),
        .O(\dso[31]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \dso[31]_i_13__0 
       (.I0(\alu1/div/chg_quo_sgn ),
        .I1(\alu1/div/dctl_stat [1]),
        .I2(\alu1/div/fdiv_rem_msb_f ),
        .O(\dso[31]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000F0002200F0FF)) 
    \dso[31]_i_14 
       (.I0(\alu0/div/dctl/dctl_sign ),
        .I1(\alu0/div/den2 ),
        .I2(\dso[31]_i_21_n_0 ),
        .I3(\alu0/div/dctl_stat [2]),
        .I4(\alu0/div/dctl_stat [0]),
        .I5(chg_quo_sgn_i_2_n_0),
        .O(\dso[31]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000F0002200F0FF)) 
    \dso[31]_i_14__0 
       (.I0(\alu1/div/dctl/dctl_sign ),
        .I1(\alu1/div/den2 ),
        .I2(\dso[31]_i_21__0_n_0 ),
        .I3(\alu1/div/dctl_stat [2]),
        .I4(\alu1/div/dctl_stat [0]),
        .I5(chg_quo_sgn_i_2__0_n_0),
        .O(\dso[31]_i_14__0_n_0 ));
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \dso[31]_i_15 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .I2(\alu0/div/dctl/dctl_long_f ),
        .I3(div_crdy0),
        .I4(\rgf/sreg/sr [8]),
        .O(\dso[31]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hEEEFFFEF)) 
    \dso[31]_i_15__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\alu1/div/dctl/dctl_long_f ),
        .I3(div_crdy1),
        .I4(\rgf/sreg/sr [8]),
        .O(\dso[31]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h331100113F110FFF)) 
    \dso[31]_i_16 
       (.I0(\alu0/div/rem [31]),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/quo__0 [31]),
        .I3(\dso[31]_i_3_n_0 ),
        .I4(\alu0/div/dso_0 [31]),
        .I5(\dso[31]_i_4_n_0 ),
        .O(\alu0/div/p_0_out [31]));
  LUT6 #(
    .INIT(64'h331100113F110FFF)) 
    \dso[31]_i_16__0 
       (.I0(\alu1/div/rem [31]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo__0 [31]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .I4(\alu1/div/dso_0 [31]),
        .I5(\dso[31]_i_4__0_n_0 ),
        .O(\alu1/div/p_0_out [31]));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_17 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [31]),
        .O(\dso[31]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_17__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [31]),
        .O(\dso[31]_i_17__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_18 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [30]),
        .O(\dso[31]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_18__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [30]),
        .O(\dso[31]_i_18__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_19 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [29]),
        .O(\dso[31]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_19__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [29]),
        .O(\dso[31]_i_19__0_n_0 ));
  LUT3 #(
    .INIT(8'hF1)) 
    \dso[31]_i_1__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .I2(\dso[31]_i_5__0_n_0 ),
        .O(\dso[31]_i_1__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_20 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [28]),
        .O(\dso[31]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[31]_i_20__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [28]),
        .O(\dso[31]_i_20__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_21 
       (.I0(\alu0/div/chg_quo_sgn ),
        .I1(\alu0/div/fdiv_rem_msb_f ),
        .O(\dso[31]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_21__0 
       (.I0(\alu1/div/chg_quo_sgn ),
        .I1(\alu1/div/fdiv_rem_msb_f ),
        .O(\dso[31]_i_21__0_n_0 ));
  LUT4 #(
    .INIT(16'h0028)) 
    \dso[31]_i_3 
       (.I0(\alu0/div/dctl_stat [3]),
        .I1(\alu0/div/dctl_stat [2]),
        .I2(\alu0/div/dctl_stat [1]),
        .I3(\dso[31]_i_13_n_0 ),
        .O(\dso[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0002000288080008)) 
    \dso[31]_i_3__0 
       (.I0(\alu1/div/dctl_stat [3]),
        .I1(\alu1/div/dctl_stat [2]),
        .I2(\dso[31]_i_13__0_n_0 ),
        .I3(\alu1/div/dctl_stat [0]),
        .I4(\alu1/div/dctl/fsm/chg_rem_sgn0 ),
        .I5(\alu1/div/dctl_stat [1]),
        .O(\dso[31]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hFB00FFFFFBFFFFFF)) 
    \dso[31]_i_4 
       (.I0(\alu0/div/dctl_stat [2]),
        .I1(\alu0/div/chg_quo_sgn ),
        .I2(\alu0/div/dctl_stat [0]),
        .I3(\alu0/div/dctl_stat [1]),
        .I4(\alu0/div/dctl_stat [3]),
        .I5(\dso[31]_i_14_n_0 ),
        .O(\dso[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFB00FFFFFBFFFFFF)) 
    \dso[31]_i_4__0 
       (.I0(\alu1/div/dctl_stat [2]),
        .I1(\alu1/div/chg_quo_sgn ),
        .I2(\alu1/div/dctl_stat [0]),
        .I3(\alu1/div/dctl_stat [1]),
        .I4(\alu1/div/dctl_stat [3]),
        .I5(\dso[31]_i_14__0_n_0 ),
        .O(\dso[31]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_5 
       (.I0(div_crdy0),
        .I1(\dctl_stat[2]_i_2_n_0 ),
        .O(\dso[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_5__0 
       (.I0(div_crdy1),
        .I1(\dctl_stat[2]_i_2__0_n_0 ),
        .O(\dso[31]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_6 
       (.I0(\alu0/div/p_0_out [30]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[31]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_6__0 
       (.I0(\alu1/div/p_0_out [30]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[31]_i_6__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_7 
       (.I0(\alu0/div/p_0_out [29]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[31]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_7__0 
       (.I0(\alu1/div/p_0_out [29]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[31]_i_7__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_8 
       (.I0(\alu0/div/p_0_out [28]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[31]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_8__0 
       (.I0(\alu1/div/p_0_out [28]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[31]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_9 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/p_0_out [31]),
        .I3(\dso[31]_i_17_n_0 ),
        .I4(\dso[31]_i_15_n_0 ),
        .I5(b0bus_0[31]),
        .O(\dso[31]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h88880FF000000FF0)) 
    \dso[31]_i_9__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/p_0_out [31]),
        .I3(\dso[31]_i_17__0_n_0 ),
        .I4(\dso[31]_i_15__0_n_0 ),
        .I5(b1bus_0[31]),
        .O(\dso[31]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [3]),
        .O(\dso[3]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [3]),
        .O(\dso[3]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [2]),
        .O(\dso[3]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [2]),
        .O(\dso[3]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [1]),
        .O(\dso[3]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[3]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [1]),
        .O(\dso[3]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'hFC77)) 
    \dso[3]_i_13 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [0]),
        .I3(\dso[31]_i_3_n_0 ),
        .O(\dso[3]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFC77)) 
    \dso[3]_i_13__0 
       (.I0(\dso[31]_i_4__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [0]),
        .I3(\dso[31]_i_3__0_n_0 ),
        .O(\dso[3]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_2 
       (.I0(\alu0/div/p_0_out [3]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_2__0 
       (.I0(\alu1/div/p_0_out [3]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_3 
       (.I0(\alu0/div/p_0_out [2]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_3__0 
       (.I0(\alu1/div/p_0_out [2]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_4 
       (.I0(\alu0/div/p_0_out [1]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_4__0 
       (.I0(\alu1/div/p_0_out [1]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_5 
       (.I0(\alu0/div/p_0_out [0]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_5__0 
       (.I0(\alu1/div/p_0_out [0]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[3]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_6 
       (.I0(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I1(\alu1/div/p_0_out [3]),
        .I2(\dso[3]_i_10__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\alu1/div/add_out [3]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_6__0 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\alu0/div/p_0_out [3]),
        .I2(\dso[3]_i_10_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\alu0/div/add_out [3]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[3]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_7 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(\alu1/div/p_0_out [2]),
        .I2(\dso[3]_i_11__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\alu1/div/add_out [2]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_7__0 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\alu0/div/p_0_out [2]),
        .I2(\dso[3]_i_11_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\alu0/div/add_out [2]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[3]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_8 
       (.I0(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I1(\alu1/div/p_0_out [1]),
        .I2(\dso[3]_i_12__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\alu1/div/add_out [1]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_8__0 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\alu0/div/p_0_out [1]),
        .I2(\dso[3]_i_12_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\alu0/div/add_out [1]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[3]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h0606F606F6F6F606)) 
    \dso[3]_i_9 
       (.I0(\alu0/div/p_0_out [0]),
        .I1(\dso[3]_i_13_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [0]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\dso[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[3]_i_9__0 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(\alu1/div/p_0_out [0]),
        .I2(\dso[3]_i_13__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\alu1/div/add_out [0]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[3]_i_9__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [7]),
        .O(\dso[7]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [7]),
        .O(\dso[7]_i_10__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_11 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [6]),
        .O(\dso[7]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_11__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [6]),
        .O(\dso[7]_i_11__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_12 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [5]),
        .O(\dso[7]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_12__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [5]),
        .O(\dso[7]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_13 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\dso[31]_i_4_n_0 ),
        .I3(\alu0/div/rem [4]),
        .O(\dso[7]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \dso[7]_i_13__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\dso[31]_i_4__0_n_0 ),
        .I3(\alu1/div/rem [4]),
        .O(\dso[7]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_2 
       (.I0(\alu0/div/p_0_out [7]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_2__0 
       (.I0(\alu1/div/p_0_out [7]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_3 
       (.I0(\alu0/div/p_0_out [6]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_3__0 
       (.I0(\alu1/div/p_0_out [6]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_4 
       (.I0(\alu0/div/p_0_out [5]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_4__0 
       (.I0(\alu1/div/p_0_out [5]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_5 
       (.I0(\alu0/div/p_0_out [4]),
        .I1(\dso[31]_i_15_n_0 ),
        .O(\dso[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_5__0 
       (.I0(\alu1/div/p_0_out [4]),
        .I1(\dso[31]_i_15__0_n_0 ),
        .O(\dso[7]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_6 
       (.I0(\alu0/div/p_0_out [7]),
        .I1(\dso[7]_i_10_n_0 ),
        .I2(\dso[31]_i_15_n_0 ),
        .I3(\alu0/div/add_out [7]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(b0bus_0[7]),
        .O(\dso[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_6__0 
       (.I0(\alu1/div/p_0_out [7]),
        .I1(\dso[7]_i_10__0_n_0 ),
        .I2(\dso[31]_i_15__0_n_0 ),
        .I3(\alu1/div/add_out [7]),
        .I4(\dso[15]_i_11__0_n_0 ),
        .I5(b1bus_0[7]),
        .O(\dso[7]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_7 
       (.I0(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .I1(\alu1/div/p_0_out [6]),
        .I2(\dso[7]_i_11__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\alu1/div/add_out [6]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_7__0 
       (.I0(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I1(\alu0/div/p_0_out [6]),
        .I2(\dso[7]_i_11_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\alu0/div/add_out [6]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[7]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_8 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\alu1/div/p_0_out [5]),
        .I2(\dso[7]_i_12__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\alu1/div/add_out [5]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_8__0 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\alu0/div/p_0_out [5]),
        .I2(\dso[7]_i_12_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\alu0/div/add_out [5]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[7]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_9 
       (.I0(\bdatw[12]_INST_0_i_4_n_0 ),
        .I1(\alu1/div/p_0_out [4]),
        .I2(\dso[7]_i_13__0_n_0 ),
        .I3(\dso[31]_i_15__0_n_0 ),
        .I4(\alu1/div/add_out [4]),
        .I5(\dso[15]_i_11__0_n_0 ),
        .O(\dso[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h553C553CFF3C003C)) 
    \dso[7]_i_9__0 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\alu0/div/p_0_out [4]),
        .I2(\dso[7]_i_13_n_0 ),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\alu0/div/add_out [4]),
        .I5(\dso[15]_i_11_n_0 ),
        .O(\dso[7]_i_9__0_n_0 ));
  CARRY4 \dso_reg[11]_i_1 
       (.CI(\dso_reg[7]_i_1_n_0 ),
        .CO({\dso_reg[11]_i_1_n_0 ,\dso_reg[11]_i_1_n_1 ,\dso_reg[11]_i_1_n_2 ,\dso_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[11]_i_2_n_0 ,\dso[11]_i_3_n_0 ,\dso[11]_i_4_n_0 ,\dso[11]_i_5_n_0 }),
        .O({\dso_reg[11]_i_1_n_4 ,\dso_reg[11]_i_1_n_5 ,\dso_reg[11]_i_1_n_6 ,\dso_reg[11]_i_1_n_7 }),
        .S({\dso[11]_i_6_n_0 ,\dso[11]_i_7_n_0 ,\dso[11]_i_8_n_0 ,\dso[11]_i_9_n_0 }));
  CARRY4 \dso_reg[11]_i_1__0 
       (.CI(\dso_reg[7]_i_1__0_n_0 ),
        .CO({\dso_reg[11]_i_1__0_n_0 ,\dso_reg[11]_i_1__0_n_1 ,\dso_reg[11]_i_1__0_n_2 ,\dso_reg[11]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[11]_i_2__0_n_0 ,\dso[11]_i_3__0_n_0 ,\dso[11]_i_4__0_n_0 ,\dso[11]_i_5__0_n_0 }),
        .O({\dso_reg[11]_i_1__0_n_4 ,\dso_reg[11]_i_1__0_n_5 ,\dso_reg[11]_i_1__0_n_6 ,\dso_reg[11]_i_1__0_n_7 }),
        .S({\dso[11]_i_6__0_n_0 ,\dso[11]_i_7__0_n_0 ,\dso[11]_i_8__0_n_0 ,\dso[11]_i_9__0_n_0 }));
  CARRY4 \dso_reg[15]_i_1 
       (.CI(\dso_reg[11]_i_1_n_0 ),
        .CO({\dso_reg[15]_i_1_n_0 ,\dso_reg[15]_i_1_n_1 ,\dso_reg[15]_i_1_n_2 ,\dso_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[15]_i_2_n_0 ,\dso[15]_i_3_n_0 ,\dso[15]_i_4_n_0 ,\dso[15]_i_5_n_0 }),
        .O({\dso_reg[15]_i_1_n_4 ,\dso_reg[15]_i_1_n_5 ,\dso_reg[15]_i_1_n_6 ,\dso_reg[15]_i_1_n_7 }),
        .S({\dso[15]_i_6_n_0 ,\dso[15]_i_7_n_0 ,\dso[15]_i_8_n_0 ,\dso[15]_i_9_n_0 }));
  CARRY4 \dso_reg[15]_i_1__0 
       (.CI(\dso_reg[11]_i_1__0_n_0 ),
        .CO({\dso_reg[15]_i_1__0_n_0 ,\dso_reg[15]_i_1__0_n_1 ,\dso_reg[15]_i_1__0_n_2 ,\dso_reg[15]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[15]_i_2__0_n_0 ,\dso[15]_i_3__0_n_0 ,\dso[15]_i_4__0_n_0 ,\dso[15]_i_5__0_n_0 }),
        .O({\dso_reg[15]_i_1__0_n_4 ,\dso_reg[15]_i_1__0_n_5 ,\dso_reg[15]_i_1__0_n_6 ,\dso_reg[15]_i_1__0_n_7 }),
        .S({\dso[15]_i_6__0_n_0 ,\dso[15]_i_7__0_n_0 ,\dso[15]_i_8__0_n_0 ,\dso[15]_i_9__0_n_0 }));
  CARRY4 \dso_reg[19]_i_1 
       (.CI(\dso_reg[15]_i_1_n_0 ),
        .CO({\dso_reg[19]_i_1_n_0 ,\dso_reg[19]_i_1_n_1 ,\dso_reg[19]_i_1_n_2 ,\dso_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[19]_i_2_n_0 ,\dso[19]_i_3_n_0 ,\dso[19]_i_4_n_0 ,\dso[19]_i_5_n_0 }),
        .O({\dso_reg[19]_i_1_n_4 ,\dso_reg[19]_i_1_n_5 ,\dso_reg[19]_i_1_n_6 ,\dso_reg[19]_i_1_n_7 }),
        .S({\dso[19]_i_6_n_0 ,\dso[19]_i_7_n_0 ,\dso[19]_i_8_n_0 ,\dso[19]_i_9_n_0 }));
  CARRY4 \dso_reg[19]_i_1__0 
       (.CI(\dso_reg[15]_i_1__0_n_0 ),
        .CO({\dso_reg[19]_i_1__0_n_0 ,\dso_reg[19]_i_1__0_n_1 ,\dso_reg[19]_i_1__0_n_2 ,\dso_reg[19]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[19]_i_2__0_n_0 ,\dso[19]_i_3__0_n_0 ,\dso[19]_i_4__0_n_0 ,\dso[19]_i_5__0_n_0 }),
        .O({\dso_reg[19]_i_1__0_n_4 ,\dso_reg[19]_i_1__0_n_5 ,\dso_reg[19]_i_1__0_n_6 ,\dso_reg[19]_i_1__0_n_7 }),
        .S({\dso[19]_i_6__0_n_0 ,\dso[19]_i_7__0_n_0 ,\dso[19]_i_8__0_n_0 ,\dso[19]_i_9__0_n_0 }));
  CARRY4 \dso_reg[23]_i_1 
       (.CI(\dso_reg[19]_i_1_n_0 ),
        .CO({\dso_reg[23]_i_1_n_0 ,\dso_reg[23]_i_1_n_1 ,\dso_reg[23]_i_1_n_2 ,\dso_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[23]_i_2_n_0 ,\dso[23]_i_3_n_0 ,\dso[23]_i_4_n_0 ,\dso[23]_i_5_n_0 }),
        .O({\dso_reg[23]_i_1_n_4 ,\dso_reg[23]_i_1_n_5 ,\dso_reg[23]_i_1_n_6 ,\dso_reg[23]_i_1_n_7 }),
        .S({\dso[23]_i_6_n_0 ,\dso[23]_i_7_n_0 ,\dso[23]_i_8_n_0 ,\dso[23]_i_9_n_0 }));
  CARRY4 \dso_reg[23]_i_1__0 
       (.CI(\dso_reg[19]_i_1__0_n_0 ),
        .CO({\dso_reg[23]_i_1__0_n_0 ,\dso_reg[23]_i_1__0_n_1 ,\dso_reg[23]_i_1__0_n_2 ,\dso_reg[23]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[23]_i_2__0_n_0 ,\dso[23]_i_3__0_n_0 ,\dso[23]_i_4__0_n_0 ,\dso[23]_i_5__0_n_0 }),
        .O({\dso_reg[23]_i_1__0_n_4 ,\dso_reg[23]_i_1__0_n_5 ,\dso_reg[23]_i_1__0_n_6 ,\dso_reg[23]_i_1__0_n_7 }),
        .S({\dso[23]_i_6__0_n_0 ,\dso[23]_i_7__0_n_0 ,\dso[23]_i_8__0_n_0 ,\dso[23]_i_9__0_n_0 }));
  CARRY4 \dso_reg[27]_i_1 
       (.CI(\dso_reg[23]_i_1_n_0 ),
        .CO({\dso_reg[27]_i_1_n_0 ,\dso_reg[27]_i_1_n_1 ,\dso_reg[27]_i_1_n_2 ,\dso_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[27]_i_2_n_0 ,\dso[27]_i_3_n_0 ,\dso[27]_i_4_n_0 ,\dso[27]_i_5_n_0 }),
        .O({\dso_reg[27]_i_1_n_4 ,\dso_reg[27]_i_1_n_5 ,\dso_reg[27]_i_1_n_6 ,\dso_reg[27]_i_1_n_7 }),
        .S({\dso[27]_i_6_n_0 ,\dso[27]_i_7_n_0 ,\dso[27]_i_8_n_0 ,\dso[27]_i_9_n_0 }));
  CARRY4 \dso_reg[27]_i_1__0 
       (.CI(\dso_reg[23]_i_1__0_n_0 ),
        .CO({\dso_reg[27]_i_1__0_n_0 ,\dso_reg[27]_i_1__0_n_1 ,\dso_reg[27]_i_1__0_n_2 ,\dso_reg[27]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[27]_i_2__0_n_0 ,\dso[27]_i_3__0_n_0 ,\dso[27]_i_4__0_n_0 ,\dso[27]_i_5__0_n_0 }),
        .O({\dso_reg[27]_i_1__0_n_4 ,\dso_reg[27]_i_1__0_n_5 ,\dso_reg[27]_i_1__0_n_6 ,\dso_reg[27]_i_1__0_n_7 }),
        .S({\dso[27]_i_6__0_n_0 ,\dso[27]_i_7__0_n_0 ,\dso[27]_i_8__0_n_0 ,\dso[27]_i_9__0_n_0 }));
  CARRY4 \dso_reg[31]_i_2 
       (.CI(\dso_reg[27]_i_1_n_0 ),
        .CO({\dso_reg[31]_i_2_n_1 ,\dso_reg[31]_i_2_n_2 ,\dso_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\dso[31]_i_6_n_0 ,\dso[31]_i_7_n_0 ,\dso[31]_i_8_n_0 }),
        .O({\dso_reg[31]_i_2_n_4 ,\dso_reg[31]_i_2_n_5 ,\dso_reg[31]_i_2_n_6 ,\dso_reg[31]_i_2_n_7 }),
        .S({\dso[31]_i_9_n_0 ,\dso[31]_i_10_n_0 ,\dso[31]_i_11_n_0 ,\dso[31]_i_12_n_0 }));
  CARRY4 \dso_reg[31]_i_2__0 
       (.CI(\dso_reg[27]_i_1__0_n_0 ),
        .CO({\dso_reg[31]_i_2__0_n_1 ,\dso_reg[31]_i_2__0_n_2 ,\dso_reg[31]_i_2__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\dso[31]_i_6__0_n_0 ,\dso[31]_i_7__0_n_0 ,\dso[31]_i_8__0_n_0 }),
        .O({\dso_reg[31]_i_2__0_n_4 ,\dso_reg[31]_i_2__0_n_5 ,\dso_reg[31]_i_2__0_n_6 ,\dso_reg[31]_i_2__0_n_7 }),
        .S({\dso[31]_i_9__0_n_0 ,\dso[31]_i_10__0_n_0 ,\dso[31]_i_11__0_n_0 ,\dso[31]_i_12__0_n_0 }));
  CARRY4 \dso_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\dso_reg[3]_i_1_n_0 ,\dso_reg[3]_i_1_n_1 ,\dso_reg[3]_i_1_n_2 ,\dso_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[3]_i_2_n_0 ,\dso[3]_i_3_n_0 ,\dso[3]_i_4_n_0 ,\dso[3]_i_5_n_0 }),
        .O({\dso_reg[3]_i_1_n_4 ,\dso_reg[3]_i_1_n_5 ,\dso_reg[3]_i_1_n_6 ,\dso_reg[3]_i_1_n_7 }),
        .S({\dso[3]_i_6__0_n_0 ,\dso[3]_i_7__0_n_0 ,\dso[3]_i_8__0_n_0 ,\dso[3]_i_9_n_0 }));
  CARRY4 \dso_reg[3]_i_1__0 
       (.CI(\<const0> ),
        .CO({\dso_reg[3]_i_1__0_n_0 ,\dso_reg[3]_i_1__0_n_1 ,\dso_reg[3]_i_1__0_n_2 ,\dso_reg[3]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[3]_i_2__0_n_0 ,\dso[3]_i_3__0_n_0 ,\dso[3]_i_4__0_n_0 ,\dso[3]_i_5__0_n_0 }),
        .O({\dso_reg[3]_i_1__0_n_4 ,\dso_reg[3]_i_1__0_n_5 ,\dso_reg[3]_i_1__0_n_6 ,\dso_reg[3]_i_1__0_n_7 }),
        .S({\dso[3]_i_6_n_0 ,\dso[3]_i_7_n_0 ,\dso[3]_i_8_n_0 ,\dso[3]_i_9__0_n_0 }));
  CARRY4 \dso_reg[7]_i_1 
       (.CI(\dso_reg[3]_i_1_n_0 ),
        .CO({\dso_reg[7]_i_1_n_0 ,\dso_reg[7]_i_1_n_1 ,\dso_reg[7]_i_1_n_2 ,\dso_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[7]_i_2_n_0 ,\dso[7]_i_3_n_0 ,\dso[7]_i_4_n_0 ,\dso[7]_i_5_n_0 }),
        .O({\dso_reg[7]_i_1_n_4 ,\dso_reg[7]_i_1_n_5 ,\dso_reg[7]_i_1_n_6 ,\dso_reg[7]_i_1_n_7 }),
        .S({\dso[7]_i_6_n_0 ,\dso[7]_i_7__0_n_0 ,\dso[7]_i_8__0_n_0 ,\dso[7]_i_9__0_n_0 }));
  CARRY4 \dso_reg[7]_i_1__0 
       (.CI(\dso_reg[3]_i_1__0_n_0 ),
        .CO({\dso_reg[7]_i_1__0_n_0 ,\dso_reg[7]_i_1__0_n_1 ,\dso_reg[7]_i_1__0_n_2 ,\dso_reg[7]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[7]_i_2__0_n_0 ,\dso[7]_i_3__0_n_0 ,\dso[7]_i_4__0_n_0 ,\dso[7]_i_5__0_n_0 }),
        .O({\dso_reg[7]_i_1__0_n_4 ,\dso_reg[7]_i_1__0_n_5 ,\dso_reg[7]_i_1__0_n_6 ,\dso_reg[7]_i_1__0_n_7 }),
        .S({\dso[7]_i_6__0_n_0 ,\dso[7]_i_7_n_0 ,\dso[7]_i_8_n_0 ,\dso[7]_i_9_n_0 }));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(\fch/eir [1]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[0]),
        .O(\eir_fl[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(\fch/eir [2]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[1]),
        .O(\eir_fl[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \eir_fl[31]_i_1 
       (.I0(fch_term),
        .I1(rst_n),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .O(\eir_fl[31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(\fch/eir [3]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[2]),
        .O(\eir_fl[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(\fch/eir [4]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[3]),
        .O(\eir_fl[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(\fch/eir [5]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[4]),
        .O(\eir_fl[5]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_1 
       (.I0(\fch/eir [6]),
        .I1(\fch_irq_lev[1]_i_2_n_0 ),
        .I2(irq_vec[5]),
        .O(\eir_fl[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8A8AAA0A8080A000)) 
    eir_inferred_i_1
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[31] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [31]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_34_n_0),
        .O(\fch/eir [31]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_10
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[22] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [22]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_43_n_0),
        .O(\fch/eir [22]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_11
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[21] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [21]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_44_n_0),
        .O(\fch/eir [21]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_12
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[20] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [20]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_45_n_0),
        .O(\fch/eir [20]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_13
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[19] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [19]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_46_n_0),
        .O(\fch/eir [19]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_14
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[18] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [18]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_47_n_0),
        .O(\fch/eir [18]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_15
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[17] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [17]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_48_n_0),
        .O(\fch/eir [17]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_16
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[16] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [16]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_49_n_0),
        .O(\fch/eir [16]));
  LUT6 #(
    .INIT(64'h00000000FF8F0000)) 
    eir_inferred_i_17
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [15]),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(eir_inferred_i_50_n_0),
        .I4(\fch/rst_n_fl ),
        .I5(eir_inferred_i_51_n_0),
        .O(\fch/eir [15]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_18
       (.I0(eir_inferred_i_52_n_0),
        .I1(eir_inferred_i_53_n_0),
        .I2(\fch/rst_n_fl ),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(eir_inferred_i_54_n_0),
        .O(\fch/eir [14]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_19
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [13]),
        .I2(eir_inferred_i_55_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_56_n_0),
        .O(\fch/eir [13]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_2
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[30] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [30]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_35_n_0),
        .O(\fch/eir [30]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_20
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [12]),
        .I2(eir_inferred_i_57_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_58_n_0),
        .O(\fch/eir [12]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_21
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [11]),
        .I2(eir_inferred_i_59_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_60_n_0),
        .O(\fch/eir [11]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_22
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [10]),
        .I2(eir_inferred_i_61_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_62_n_0),
        .O(\fch/eir [10]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_23
       (.I0(eir_inferred_i_63_n_0),
        .I1(eir_inferred_i_64_n_0),
        .I2(\fch/rst_n_fl ),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(eir_inferred_i_65_n_0),
        .O(\fch/eir [9]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_24
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [8]),
        .I2(eir_inferred_i_66_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_67_n_0),
        .O(\fch/eir [8]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_25
       (.I0(eir_inferred_i_68_n_0),
        .I1(eir_inferred_i_69_n_0),
        .I2(\fch/rst_n_fl ),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(eir_inferred_i_70_n_0),
        .O(\fch/eir [7]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_26
       (.I0(eir_inferred_i_71_n_0),
        .I1(eir_inferred_i_72_n_0),
        .I2(\fch/rst_n_fl ),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(eir_inferred_i_73_n_0),
        .O(\fch/eir [6]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_27
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [5]),
        .I2(eir_inferred_i_74_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_75_n_0),
        .O(\fch/eir [5]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_28
       (.I0(eir_inferred_i_76_n_0),
        .I1(eir_inferred_i_77_n_0),
        .I2(\fch/rst_n_fl ),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(eir_inferred_i_78_n_0),
        .O(\fch/eir [4]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_29
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [3]),
        .I2(eir_inferred_i_79_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_80_n_0),
        .O(\fch/eir [3]));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_3
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[29] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [29]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_36_n_0),
        .O(\fch/eir [29]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_30
       (.I0(eir_inferred_i_81_n_0),
        .I1(eir_inferred_i_82_n_0),
        .I2(\fch/rst_n_fl ),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(eir_inferred_i_83_n_0),
        .O(\fch/eir [2]));
  LUT5 #(
    .INIT(32'hE0E0E000)) 
    eir_inferred_i_31
       (.I0(eir_inferred_i_84_n_0),
        .I1(eir_inferred_i_85_n_0),
        .I2(\fch/rst_n_fl ),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(eir_inferred_i_86_n_0),
        .O(\fch/eir [1]));
  LUT6 #(
    .INIT(64'hF800FF00F8000000)) 
    eir_inferred_i_32
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/data0 [0]),
        .I2(eir_inferred_i_87_n_0),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/ctl_fetch_ext_fl ),
        .I5(eir_inferred_i_88_n_0),
        .O(\fch/eir [0]));
  LUT3 #(
    .INIT(8'h01)) 
    eir_inferred_i_33
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/fch_leir_lir ),
        .I2(\fch/fch_leir_hir ),
        .O(eir_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_34
       (.I0(\fch/data0 [15]),
        .I1(fdat[31]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/eir_fl_reg_n_0_[31] ),
        .O(eir_inferred_i_34_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_35
       (.I0(\fch/data0 [14]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[30]),
        .I3(\fch/eir_fl_reg_n_0_[30] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_35_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_36
       (.I0(\fch/data0 [13]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[29]),
        .I3(\fch/eir_fl_reg_n_0_[29] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_37
       (.I0(\fch/data0 [12]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[28]),
        .I3(\fch/eir_fl_reg_n_0_[28] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_38
       (.I0(\fch/data0 [11]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[27]),
        .I3(\fch/eir_fl_reg_n_0_[27] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_39
       (.I0(\fch/data0 [10]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[26]),
        .I3(\fch/eir_fl_reg_n_0_[26] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_4
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[28] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [28]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_37_n_0),
        .O(\fch/eir [28]));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_40
       (.I0(\fch/data0 [9]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[25]),
        .I3(\fch/eir_fl_reg_n_0_[25] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_41
       (.I0(\fch/data0 [8]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[24]),
        .I3(\fch/eir_fl_reg_n_0_[24] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_42
       (.I0(\fch/data0 [7]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[23]),
        .I3(\fch/eir_fl_reg_n_0_[23] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_42_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_43
       (.I0(\fch/data0 [6]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[22]),
        .I3(\fch/eir_fl_reg_n_0_[22] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_43_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_44
       (.I0(\fch/data0 [5]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[21]),
        .I3(\fch/eir_fl_reg_n_0_[21] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_44_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_45
       (.I0(\fch/data0 [4]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[20]),
        .I3(\fch/eir_fl_reg_n_0_[20] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_45_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_46
       (.I0(\fch/data0 [3]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[19]),
        .I3(\fch/eir_fl_reg_n_0_[19] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_47
       (.I0(\fch/data0 [2]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[18]),
        .I3(\fch/eir_fl_reg_n_0_[18] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_47_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_48
       (.I0(\fch/data0 [1]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[17]),
        .I3(\fch/eir_fl_reg_n_0_[17] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_48_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF474700FF)) 
    eir_inferred_i_49
       (.I0(\fch/data0 [0]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[16]),
        .I3(\fch/eir_fl_reg_n_0_[16] ),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_5
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[27] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [27]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_38_n_0),
        .O(\fch/eir [27]));
  LUT6 #(
    .INIT(64'h3033300030223022)) 
    eir_inferred_i_50
       (.I0(\fch/data0 [31]),
        .I1(\fch/fch_leir_nir ),
        .I2(fdat[31]),
        .I3(\fch/fch_leir_hir ),
        .I4(fdat[15]),
        .I5(\fch/fch_leir_lir ),
        .O(eir_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'h00000000474700FF)) 
    eir_inferred_i_51
       (.I0(fdat[31]),
        .I1(\fch/fch_heir_nir ),
        .I2(fdat[15]),
        .I3(\fch/data0 [31]),
        .I4(eir_inferred_i_89_n_0),
        .I5(\fch/ctl_fetch_ext_fl ),
        .O(eir_inferred_i_51_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_52
       (.I0(\fch/fch_leir_lir ),
        .I1(\fch/fch_leir_hir ),
        .I2(\fch/data0 [30]),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(\fch/data0 [14]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_52_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_53
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/fch_leir_lir ),
        .I2(fdat[14]),
        .I3(\fch/fch_leir_hir ),
        .I4(fdat[30]),
        .O(eir_inferred_i_53_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_54
       (.I0(fdat[30]),
        .I1(fdat[14]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [30]),
        .O(eir_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_55
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[29]),
        .I2(\fch/fch_leir_hir ),
        .I3(fdat[13]),
        .I4(\fch/fch_leir_lir ),
        .I5(\fch/data0 [29]),
        .O(eir_inferred_i_55_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_56
       (.I0(fdat[29]),
        .I1(fdat[13]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [29]),
        .O(eir_inferred_i_56_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_57
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[28]),
        .I2(\fch/fch_leir_hir ),
        .I3(fdat[12]),
        .I4(\fch/fch_leir_lir ),
        .I5(\fch/data0 [28]),
        .O(eir_inferred_i_57_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_58
       (.I0(fdat[28]),
        .I1(fdat[12]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [28]),
        .O(eir_inferred_i_58_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_59
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[27]),
        .I2(\fch/fch_leir_hir ),
        .I3(fdat[11]),
        .I4(\fch/fch_leir_lir ),
        .I5(\fch/data0 [27]),
        .O(eir_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_6
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[26] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [26]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_39_n_0),
        .O(\fch/eir [26]));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_60
       (.I0(fdat[27]),
        .I1(fdat[11]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [27]),
        .O(eir_inferred_i_60_n_0));
  LUT6 #(
    .INIT(64'h4545454040404540)) 
    eir_inferred_i_61
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[26]),
        .I2(\fch/fch_leir_hir ),
        .I3(\fch/data0 [26]),
        .I4(\fch/fch_leir_lir ),
        .I5(fdat[10]),
        .O(eir_inferred_i_61_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_62
       (.I0(fdat[26]),
        .I1(fdat[10]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [26]),
        .O(eir_inferred_i_62_n_0));
  LUT6 #(
    .INIT(64'hD5D5D5DFD5D5D5D5)) 
    eir_inferred_i_63
       (.I0(\fch/ctl_fetch_ext_fl ),
        .I1(\fch/data0 [9]),
        .I2(\fch/fch_leir_nir ),
        .I3(\fch/fch_leir_lir ),
        .I4(\fch/fch_leir_hir ),
        .I5(\fch/data0 [25]),
        .O(eir_inferred_i_63_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_64
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/fch_leir_lir ),
        .I2(fdat[9]),
        .I3(\fch/fch_leir_hir ),
        .I4(fdat[25]),
        .O(eir_inferred_i_64_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_65
       (.I0(fdat[25]),
        .I1(fdat[9]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [25]),
        .O(eir_inferred_i_65_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_66
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[24]),
        .I2(\fch/fch_leir_hir ),
        .I3(fdat[8]),
        .I4(\fch/fch_leir_lir ),
        .I5(\fch/data0 [24]),
        .O(eir_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_67
       (.I0(fdat[24]),
        .I1(fdat[8]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [24]),
        .O(eir_inferred_i_67_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_68
       (.I0(\fch/fch_leir_lir ),
        .I1(\fch/fch_leir_hir ),
        .I2(\fch/data0 [23]),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(\fch/data0 [7]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_68_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_69
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/fch_leir_lir ),
        .I2(fdat[7]),
        .I3(\fch/fch_leir_hir ),
        .I4(fdat[23]),
        .O(eir_inferred_i_69_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_7
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[25] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [25]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_40_n_0),
        .O(\fch/eir [25]));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_70
       (.I0(fdat[23]),
        .I1(fdat[7]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [23]),
        .O(eir_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'hD5D5D5DFD5D5D5D5)) 
    eir_inferred_i_71
       (.I0(\fch/ctl_fetch_ext_fl ),
        .I1(\fch/data0 [6]),
        .I2(\fch/fch_leir_nir ),
        .I3(\fch/fch_leir_lir ),
        .I4(\fch/fch_leir_hir ),
        .I5(\fch/data0 [22]),
        .O(eir_inferred_i_71_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_72
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/fch_leir_lir ),
        .I2(fdat[6]),
        .I3(\fch/fch_leir_hir ),
        .I4(fdat[22]),
        .O(eir_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_73
       (.I0(fdat[22]),
        .I1(fdat[6]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [22]),
        .O(eir_inferred_i_73_n_0));
  LUT6 #(
    .INIT(64'h4540454545404040)) 
    eir_inferred_i_74
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[21]),
        .I2(\fch/fch_leir_hir ),
        .I3(fdat[5]),
        .I4(\fch/fch_leir_lir ),
        .I5(\fch/data0 [21]),
        .O(eir_inferred_i_74_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_75
       (.I0(fdat[21]),
        .I1(fdat[5]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [21]),
        .O(eir_inferred_i_75_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_76
       (.I0(\fch/fch_leir_lir ),
        .I1(\fch/fch_leir_hir ),
        .I2(\fch/data0 [20]),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(\fch/data0 [4]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_76_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_77
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/fch_leir_lir ),
        .I2(fdat[4]),
        .I3(\fch/fch_leir_hir ),
        .I4(fdat[20]),
        .O(eir_inferred_i_77_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_78
       (.I0(fdat[20]),
        .I1(fdat[4]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [20]),
        .O(eir_inferred_i_78_n_0));
  LUT6 #(
    .INIT(64'h4545454040404540)) 
    eir_inferred_i_79
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[19]),
        .I2(\fch/fch_leir_hir ),
        .I3(\fch/data0 [19]),
        .I4(\fch/fch_leir_lir ),
        .I5(fdat[3]),
        .O(eir_inferred_i_79_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_8
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[24] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [24]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_41_n_0),
        .O(\fch/eir [24]));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_80
       (.I0(fdat[19]),
        .I1(fdat[3]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [19]),
        .O(eir_inferred_i_80_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_81
       (.I0(\fch/fch_leir_lir ),
        .I1(\fch/fch_leir_hir ),
        .I2(\fch/data0 [18]),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(\fch/data0 [2]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_81_n_0));
  LUT5 #(
    .INIT(32'h0000F808)) 
    eir_inferred_i_82
       (.I0(\fch/fch_leir_lir ),
        .I1(fdat[2]),
        .I2(\fch/fch_leir_hir ),
        .I3(fdat[18]),
        .I4(\fch/fch_leir_nir ),
        .O(eir_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_83
       (.I0(fdat[18]),
        .I1(fdat[2]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [18]),
        .O(eir_inferred_i_83_n_0));
  LUT6 #(
    .INIT(64'hFFFF00FF10FF10FF)) 
    eir_inferred_i_84
       (.I0(\fch/fch_leir_lir ),
        .I1(\fch/fch_leir_hir ),
        .I2(\fch/data0 [17]),
        .I3(\fch/ctl_fetch_ext_fl ),
        .I4(\fch/data0 [1]),
        .I5(\fch/fch_leir_nir ),
        .O(eir_inferred_i_84_n_0));
  LUT5 #(
    .INIT(32'h55400040)) 
    eir_inferred_i_85
       (.I0(\fch/fch_leir_nir ),
        .I1(\fch/fch_leir_lir ),
        .I2(fdat[1]),
        .I3(\fch/fch_leir_hir ),
        .I4(fdat[17]),
        .O(eir_inferred_i_85_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_86
       (.I0(fdat[17]),
        .I1(fdat[1]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [17]),
        .O(eir_inferred_i_86_n_0));
  LUT6 #(
    .INIT(64'h4545454040404540)) 
    eir_inferred_i_87
       (.I0(\fch/fch_leir_nir ),
        .I1(fdat[16]),
        .I2(\fch/fch_leir_hir ),
        .I3(\fch/data0 [16]),
        .I4(\fch/fch_leir_lir ),
        .I5(fdat[0]),
        .O(eir_inferred_i_87_n_0));
  LUT6 #(
    .INIT(64'hAFAFCFFFA0A0C000)) 
    eir_inferred_i_88
       (.I0(fdat[16]),
        .I1(fdat[0]),
        .I2(\fch/ctl_fetch_lng_fl ),
        .I3(\fch/fch_heir_hir ),
        .I4(\fch/fch_heir_nir ),
        .I5(\fch/data0 [16]),
        .O(eir_inferred_i_88_n_0));
  LUT3 #(
    .INIT(8'hA8)) 
    eir_inferred_i_89
       (.I0(\fch/ctl_fetch_lng_fl ),
        .I1(\fch/fch_heir_hir ),
        .I2(\fch/fch_heir_nir ),
        .O(eir_inferred_i_89_n_0));
  LUT6 #(
    .INIT(64'h8080A000AAAAAAAA)) 
    eir_inferred_i_9
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/eir_fl_reg_n_0_[23] ),
        .I2(\fch/ctl_fetch_ext_fl ),
        .I3(\fch/data0 [23]),
        .I4(eir_inferred_i_33_n_0),
        .I5(eir_inferred_i_42_n_0),
        .O(\fch/eir [23]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[10]_INST_0 
       (.I0(\fch/p_2_in [10]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [10]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[12]_INST_0_i_1_n_6 ),
        .O(\^fadr [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[11]_INST_0 
       (.I0(\fch/p_2_in [11]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [11]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[12]_INST_0_i_1_n_5 ),
        .O(\^fadr [11]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[11]_INST_0_i_1 
       (.CI(\fadr[7]_INST_0_i_1_n_0 ),
        .CO({\fadr[11]_INST_0_i_1_n_0 ,\fadr[11]_INST_0_i_1_n_1 ,\fadr[11]_INST_0_i_1_n_2 ,\fadr[11]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in [11:8]),
        .S(\rgf/pcnt/pc [11:8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[12]_INST_0 
       (.I0(\fch/p_2_in [12]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [12]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[12]_INST_0_i_1_n_4 ),
        .O(\^fadr [12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[12]_INST_0_i_1 
       (.CI(\fadr[8]_INST_0_i_1_n_0 ),
        .CO({\fadr[12]_INST_0_i_1_n_0 ,\fadr[12]_INST_0_i_1_n_1 ,\fadr[12]_INST_0_i_1_n_2 ,\fadr[12]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fadr[12]_INST_0_i_1_n_4 ,\fadr[12]_INST_0_i_1_n_5 ,\fadr[12]_INST_0_i_1_n_6 ,\fadr[12]_INST_0_i_1_n_7 }),
        .S(\rgf/pcnt/pc [12:9]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[13]_INST_0 
       (.I0(\fch/p_2_in [13]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [13]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[15]_INST_0_i_4_n_7 ),
        .O(\^fadr [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[14]_INST_0 
       (.I0(\fch/p_2_in [14]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [14]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[15]_INST_0_i_4_n_6 ),
        .O(\^fadr [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[15]_INST_0 
       (.I0(\fch/p_2_in [15]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [15]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[15]_INST_0_i_4_n_5 ),
        .O(\^fadr [15]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[15]_INST_0_i_1 
       (.CI(\fadr[11]_INST_0_i_1_n_0 ),
        .CO({\fadr[15]_INST_0_i_1_n_1 ,\fadr[15]_INST_0_i_1_n_2 ,\fadr[15]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in [15:12]),
        .S(\rgf/pcnt/pc [15:12]));
  LUT2 #(
    .INIT(4'h8)) 
    \fadr[15]_INST_0_i_10 
       (.I0(\fadr[15]_INST_0_i_6_n_0 ),
        .I1(fch_heir_nir_i_3_n_0),
        .O(\fadr[15]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0100010101000000)) 
    \fadr[15]_INST_0_i_11 
       (.I0(\fadr[15]_INST_0_i_8_n_0 ),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [2]),
        .I3(\fch/fch_issu1 ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/fch_issu1_fl ),
        .O(\fadr[15]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \fadr[15]_INST_0_i_12 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [3]),
        .O(\fadr[15]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \fadr[15]_INST_0_i_13 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [12]),
        .I4(\fadr[15]_INST_0_i_17_n_0 ),
        .O(\fadr[15]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \fadr[15]_INST_0_i_14 
       (.I0(\nir_id[24]_i_6_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [10]),
        .O(\fadr[15]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h1555)) 
    \fadr[15]_INST_0_i_15 
       (.I0(\fch/ctl_bcc_take1_fl ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .O(\fadr[15]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFD555FFFFFFFF)) 
    \fadr[15]_INST_0_i_16 
       (.I0(\fadr[15]_INST_0_i_15_n_0 ),
        .I1(stat[1]),
        .I2(stat[2]),
        .I3(stat[0]),
        .I4(\fch/ctl_bcc_take0_fl ),
        .I5(fch_term),
        .O(\fadr[15]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \fadr[15]_INST_0_i_17 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [1]),
        .O(\fadr[15]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    \fadr[15]_INST_0_i_2 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fadr[15]_INST_0_i_6_n_0 ),
        .I4(\fadr[15]_INST_0_i_7_n_0 ),
        .I5(\fadr[15]_INST_0_i_8_n_0 ),
        .O(\fadr[15]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h5155FFFF)) 
    \fadr[15]_INST_0_i_3 
       (.I0(\fadr[15]_INST_0_i_9_n_0 ),
        .I1(\fch/stat [1]),
        .I2(\fadr[15]_INST_0_i_10_n_0 ),
        .I3(\fadr[15]_INST_0_i_11_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\fadr[15]_INST_0_i_3_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[15]_INST_0_i_4 
       (.CI(\fadr[12]_INST_0_i_1_n_0 ),
        .CO({\fadr[15]_INST_0_i_4_n_2 ,\fadr[15]_INST_0_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fadr[15]_INST_0_i_4_n_5 ,\fadr[15]_INST_0_i_4_n_6 ,\fadr[15]_INST_0_i_4_n_7 }),
        .S({\<const0> ,\rgf/pcnt/pc [15:13]}));
  LUT6 #(
    .INIT(64'hAAAAA8AAAAAAAAAA)) 
    \fadr[15]_INST_0_i_5 
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [15]),
        .I3(\fadr[15]_INST_0_i_12_n_0 ),
        .I4(\fadr[15]_INST_0_i_13_n_0 ),
        .I5(\fadr[15]_INST_0_i_14_n_0 ),
        .O(\fadr[15]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \fadr[15]_INST_0_i_6 
       (.I0(\nir_id[24]_i_6_n_0 ),
        .I1(fch_term),
        .O(\fadr[15]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fadr[15]_INST_0_i_7 
       (.I0(\fch/stat [2]),
        .I1(fch_heir_nir_i_3_n_0),
        .O(\fadr[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFD55500000000)) 
    \fadr[15]_INST_0_i_8 
       (.I0(\fadr[15]_INST_0_i_15_n_0 ),
        .I1(stat[1]),
        .I2(stat[2]),
        .I3(stat[0]),
        .I4(\fch/ctl_bcc_take0_fl ),
        .I5(fch_term),
        .O(\fadr[15]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \fadr[15]_INST_0_i_9 
       (.I0(\fadr[15]_INST_0_i_16_n_0 ),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [1]),
        .I3(\fch/stat [2]),
        .O(\fadr[15]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[1]_INST_0 
       (.I0(\fch/p_2_in [1]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [1]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[4]_INST_0_i_1_n_7 ),
        .O(\^fadr [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[2]_INST_0 
       (.I0(\fch/p_2_in [2]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [2]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[4]_INST_0_i_1_n_6 ),
        .O(\^fadr [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[3]_INST_0 
       (.I0(\fch/p_2_in [3]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [3]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[4]_INST_0_i_1_n_5 ),
        .O(\^fadr [3]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[3]_INST_0_i_1 
       (.CI(\<const0> ),
        .CO({\fadr[3]_INST_0_i_1_n_0 ,\fadr[3]_INST_0_i_1_n_1 ,\fadr[3]_INST_0_i_1_n_2 ,\fadr[3]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/pcnt/pc [1],\<const0> }),
        .O({\fch/p_2_in [3:1],\fch/p_2_in0_in [0]}),
        .S({\rgf/pcnt/pc [3:2],\fadr[3]_INST_0_i_2_n_0 ,\rgf/pcnt/pc [0]}));
  LUT1 #(
    .INIT(2'h1)) 
    \fadr[3]_INST_0_i_2 
       (.I0(\rgf/pcnt/pc [1]),
        .O(\fadr[3]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[4]_INST_0 
       (.I0(\fch/p_2_in [4]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [4]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[4]_INST_0_i_1_n_4 ),
        .O(\^fadr [4]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[4]_INST_0_i_1 
       (.CI(\<const0> ),
        .CO({\fadr[4]_INST_0_i_1_n_0 ,\fadr[4]_INST_0_i_1_n_1 ,\fadr[4]_INST_0_i_1_n_2 ,\fadr[4]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\rgf/pcnt/pc [2],\<const0> }),
        .O({\fadr[4]_INST_0_i_1_n_4 ,\fadr[4]_INST_0_i_1_n_5 ,\fadr[4]_INST_0_i_1_n_6 ,\fadr[4]_INST_0_i_1_n_7 }),
        .S({\rgf/pcnt/pc [4:3],\fadr[4]_INST_0_i_2_n_0 ,\rgf/pcnt/pc [1]}));
  LUT1 #(
    .INIT(2'h1)) 
    \fadr[4]_INST_0_i_2 
       (.I0(\rgf/pcnt/pc [2]),
        .O(\fadr[4]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[5]_INST_0 
       (.I0(\fch/p_2_in [5]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [5]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[8]_INST_0_i_1_n_7 ),
        .O(\^fadr [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[6]_INST_0 
       (.I0(\fch/p_2_in [6]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [6]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[8]_INST_0_i_1_n_6 ),
        .O(\^fadr [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[7]_INST_0 
       (.I0(\fch/p_2_in [7]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [7]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[8]_INST_0_i_1_n_5 ),
        .O(\^fadr [7]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[7]_INST_0_i_1 
       (.CI(\fadr[3]_INST_0_i_1_n_0 ),
        .CO({\fadr[7]_INST_0_i_1_n_0 ,\fadr[7]_INST_0_i_1_n_1 ,\fadr[7]_INST_0_i_1_n_2 ,\fadr[7]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in [7:4]),
        .S(\rgf/pcnt/pc [7:4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[8]_INST_0 
       (.I0(\fch/p_2_in [8]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [8]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[8]_INST_0_i_1_n_4 ),
        .O(\^fadr [8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \fadr[8]_INST_0_i_1 
       (.CI(\fadr[4]_INST_0_i_1_n_0 ),
        .CO({\fadr[8]_INST_0_i_1_n_0 ,\fadr[8]_INST_0_i_1_n_1 ,\fadr[8]_INST_0_i_1_n_2 ,\fadr[8]_INST_0_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\fadr[8]_INST_0_i_1_n_4 ,\fadr[8]_INST_0_i_1_n_5 ,\fadr[8]_INST_0_i_1_n_6 ,\fadr[8]_INST_0_i_1_n_7 }),
        .S(\rgf/pcnt/pc [8:5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \fadr[9]_INST_0 
       (.I0(\fch/p_2_in [9]),
        .I1(\fadr[15]_INST_0_i_2_n_0 ),
        .I2(\rgf/pcnt/pc [9]),
        .I3(\fadr[15]_INST_0_i_3_n_0 ),
        .I4(\fadr[12]_INST_0_i_1_n_7 ),
        .O(\^fadr [9]));
  FDRE \fch/ctl_bcc_take0_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take0_fl_i_2_n_0),
        .Q(\fch/ctl_bcc_take0_fl ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/ctl_bcc_take1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_bcc_take1_fl_i_1_n_0),
        .Q(\fch/ctl_bcc_take1_fl ),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/ctl_fetch0_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch0),
        .Q(\fch/ctl_fetch0_fl ),
        .R(\<const0> ));
  FDRE \fch/ctl_fetch1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch1),
        .Q(\fch/ctl_fetch1_fl ),
        .R(\<const0> ));
  FDRE \fch/ctl_fetch_ext_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ctl_fetch_ext ),
        .Q(\fch/ctl_fetch_ext_fl ),
        .R(\<const0> ));
  FDRE \fch/ctl_fetch_lng_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ctl_fetch_lng ),
        .Q(\fch/ctl_fetch_lng_fl ),
        .R(\<const0> ));
  FDRE \fch/eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [0]),
        .Q(\fch/data0 [16]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [10]),
        .Q(\fch/data0 [26]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [11]),
        .Q(\fch/data0 [27]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [12]),
        .Q(\fch/data0 [28]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [13]),
        .Q(\fch/data0 [29]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [14]),
        .Q(\fch/data0 [30]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [15]),
        .Q(\fch/data0 [31]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [16]),
        .Q(\fch/eir_fl_reg_n_0_[16] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [17]),
        .Q(\fch/eir_fl_reg_n_0_[17] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [18]),
        .Q(\fch/eir_fl_reg_n_0_[18] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [19]),
        .Q(\fch/eir_fl_reg_n_0_[19] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[1]_i_1_n_0 ),
        .Q(\fch/data0 [17]),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/eir_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [20]),
        .Q(\fch/eir_fl_reg_n_0_[20] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [21]),
        .Q(\fch/eir_fl_reg_n_0_[21] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [22]),
        .Q(\fch/eir_fl_reg_n_0_[22] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [23]),
        .Q(\fch/eir_fl_reg_n_0_[23] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [24]),
        .Q(\fch/eir_fl_reg_n_0_[24] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [25]),
        .Q(\fch/eir_fl_reg_n_0_[25] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [26]),
        .Q(\fch/eir_fl_reg_n_0_[26] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [27]),
        .Q(\fch/eir_fl_reg_n_0_[27] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [28]),
        .Q(\fch/eir_fl_reg_n_0_[28] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [29]),
        .Q(\fch/eir_fl_reg_n_0_[29] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[2]_i_1_n_0 ),
        .Q(\fch/data0 [18]),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/eir_fl_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [30]),
        .Q(\fch/eir_fl_reg_n_0_[30] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [31]),
        .Q(\fch/eir_fl_reg_n_0_[31] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[3]_i_1_n_0 ),
        .Q(\fch/data0 [19]),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[4]_i_1_n_0 ),
        .Q(\fch/data0 [20]),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[5]_i_1_n_0 ),
        .Q(\fch/data0 [21]),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[6]_i_1_n_0 ),
        .Q(\fch/data0 [22]),
        .R(ctl_bcc_take0_fl_i_1_n_0));
  FDRE \fch/eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [7]),
        .Q(\fch/data0 [23]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [8]),
        .Q(\fch/data0 [24]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/eir [9]),
        .Q(\fch/data0 [25]),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \fch/fadr_1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\^fadr [1]),
        .Q(\fch/fadr_1_fl ),
        .R(\<const0> ));
  FDRE \fch/fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[0]_i_1_n_0 ),
        .Q(fch_irq_lev[0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[1]_i_1_n_0 ),
        .Q(fch_irq_lev[1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/fch_irq_req_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(\fch/fch_irq_req_fl ),
        .R(\<const0> ));
  FDRE \fch/fch_issu1_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fch_issu1_ir ),
        .Q(\fch/fch_issu1_fl ),
        .R(\<const0> ));
  FDRE \fch/fch_term_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(\fch/fch_term_fl ),
        .R(\<const0> ));
  FDRE \fch/fctl/fch_heir_hir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_heir_hir_t ),
        .Q(\fch/fch_heir_hir ),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/fctl/fch_heir_nir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_heir_nir_t ),
        .Q(\fch/fch_heir_nir ),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/fctl/fch_leir_hir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_leir_hir_t ),
        .Q(\fch/fch_leir_hir ),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/fctl/fch_leir_lir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_leir_lir_t ),
        .Q(\fch/fch_leir_lir ),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/fctl/fch_leir_nir_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/fch_leir_nir_t ),
        .Q(\fch/fch_leir_nir ),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/fctl/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/stat_nx [0]),
        .Q(\fch/stat [0]),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/fctl/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/stat_nx [1]),
        .Q(\fch/stat [1]),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/fctl/stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/fctl/stat_nx [2]),
        .Q(\fch/stat [2]),
        .R(\stat[2]_i_1_n_0 ));
  FDRE \fch/ir0_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [0]),
        .Q(\fch/ir0_fl [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [10]),
        .Q(\fch/ir0_fl [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [11]),
        .Q(\fch/ir0_fl [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [12]),
        .Q(\fch/ir0_fl [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [13]),
        .Q(\fch/ir0_fl [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [14]),
        .Q(\fch/ir0_fl [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [15]),
        .Q(\fch/ir0_fl [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [1]),
        .Q(\fch/ir0_fl [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [2]),
        .Q(\fch/ir0_fl [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [3]),
        .Q(\fch/ir0_fl [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [4]),
        .Q(\fch/ir0_fl [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [5]),
        .Q(\fch/ir0_fl [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [6]),
        .Q(\fch/ir0_fl [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [7]),
        .Q(\fch/ir0_fl [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [8]),
        .Q(\fch/ir0_fl [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir0 [9]),
        .Q(\fch/ir0_fl [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ir0_id_fl[20]_i_1_n_0 ),
        .Q(\fch/ir0_id_fl [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir0_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\ir0_id_fl[21]_i_1_n_0 ),
        .Q(\fch/ir0_id_fl [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [0]),
        .Q(\fch/ir1_fl [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [10]),
        .Q(\fch/ir1_fl [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [11]),
        .Q(\fch/ir1_fl [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [12]),
        .Q(\fch/ir1_fl [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [13]),
        .Q(\fch/ir1_fl [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [14]),
        .Q(\fch/ir1_fl [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [15]),
        .Q(\fch/ir1_fl [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [1]),
        .Q(\fch/ir1_fl [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [2]),
        .Q(\fch/ir1_fl [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [3]),
        .Q(\fch/ir1_fl [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [4]),
        .Q(\fch/ir1_fl [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [5]),
        .Q(\fch/ir1_fl [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [6]),
        .Q(\fch/ir1_fl [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [7]),
        .Q(\fch/ir1_fl [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [8]),
        .Q(\fch/ir1_fl [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch/ir1 [9]),
        .Q(\fch/ir1_fl [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_id_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_wrbufn1),
        .Q(\fch/ir1_id_fl [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/ir1_id_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_memacc1),
        .Q(\fch/ir1_id_fl [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[12] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [12]),
        .Q(\fch/nir_id [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[13] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [13]),
        .Q(\fch/nir_id [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[14] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [14]),
        .Q(\fch/nir_id [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[15] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [15]),
        .Q(\fch/nir_id [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[16] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [16]),
        .Q(\fch/nir_id [16]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[17] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [17]),
        .Q(\fch/nir_id [17]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[18] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [18]),
        .Q(\fch/nir_id [18]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[19] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [19]),
        .Q(\fch/nir_id [19]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[20] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\nir_id[20]_i_1_n_0 ),
        .Q(\fch/nir_id [20]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[21] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [21]),
        .Q(\fch/nir_id [21]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_id_reg[24] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(\fch/lir_id_0 [24]),
        .Q(\fch/nir_id [24]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[0] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[0]),
        .Q(\fch/data0 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[10] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[10]),
        .Q(\fch/data0 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[11] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[11]),
        .Q(\fch/data0 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[12] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[12]),
        .Q(\fch/data0 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[13] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[13]),
        .Q(\fch/data0 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[14] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[14]),
        .Q(\fch/data0 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[15] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[15]),
        .Q(\fch/data0 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[1] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[1]),
        .Q(\fch/data0 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[2] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[2]),
        .Q(\fch/data0 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[3] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[3]),
        .Q(\fch/data0 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[4] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[4]),
        .Q(\fch/data0 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[5] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[5]),
        .Q(\fch/data0 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[6] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[6]),
        .Q(\fch/data0 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[7] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[7]),
        .Q(\fch/data0 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[8] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[8]),
        .Q(\fch/data0 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/nir_reg[9] 
       (.C(clk),
        .CE(\fch/fctl/fch_nir_lir ),
        .D(fdat[9]),
        .Q(\fch/data0 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[0]),
        .Q(fch_pc0[0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[10]),
        .Q(fch_pc0[10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[11]),
        .Q(fch_pc0[11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[12]),
        .Q(fch_pc0[12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[13]),
        .Q(fch_pc0[13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[14]),
        .Q(fch_pc0[14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[15]),
        .Q(fch_pc0[15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[1]),
        .Q(fch_pc0[1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[2]),
        .Q(fch_pc0[2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[3]),
        .Q(fch_pc0[3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[4]),
        .Q(fch_pc0[4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[5]),
        .Q(fch_pc0[5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[6]),
        .Q(fch_pc0[6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[7]),
        .Q(fch_pc0[7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[8]),
        .Q(fch_pc0[8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc0_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(fch_pc[9]),
        .Q(fch_pc0[9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[0] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[3]_i_1_n_7 ),
        .Q(fch_pc1[0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[10] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[11]_i_1_n_5 ),
        .Q(fch_pc1[10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[11] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[11]_i_1_n_4 ),
        .Q(fch_pc1[11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[12] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_i_1_n_7 ),
        .Q(fch_pc1[12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[13] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_i_1_n_6 ),
        .Q(fch_pc1[13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[14] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_i_1_n_5 ),
        .Q(fch_pc1[14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[15] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[15]_i_1_n_4 ),
        .Q(fch_pc1[15]),
        .R(\alu1/div/p_0_in__0 ));
  FDSE \fch/pc1_reg[1] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[3]_i_1_n_6 ),
        .Q(fch_pc1[1]),
        .S(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[2] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[3]_i_1_n_5 ),
        .Q(fch_pc1[2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[3] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[3]_i_1_n_4 ),
        .Q(fch_pc1[3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[4] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[7]_i_1_n_7 ),
        .Q(fch_pc1[4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[5] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[7]_i_1_n_6 ),
        .Q(fch_pc1[5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[6] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[7]_i_1_n_5 ),
        .Q(fch_pc1[6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[7] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[7]_i_1_n_4 ),
        .Q(fch_pc1[7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[8] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[11]_i_1_n_7 ),
        .Q(fch_pc1[8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/pc1_reg[9] 
       (.C(clk),
        .CE(fch_term),
        .D(\pc1_reg[11]_i_1_n_6 ),
        .Q(fch_pc1[9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \fch/rst_n_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(\fch/rst_n_fl ),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0228000000000000)) 
    fch_heir_hir_i_1
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\fch/fch_issu1_ir ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(\fadr[15]_INST_0_i_6_n_0 ),
        .I5(\fadr[15]_INST_0_i_7_n_0 ),
        .O(\fch/fctl/fch_heir_hir_t ));
  LUT6 #(
    .INIT(64'h0000000088822282)) 
    fch_heir_nir_i_1
       (.I0(fch_heir_nir_i_2_n_0),
        .I1(\fch/stat [1]),
        .I2(\fch/fch_issu1_fl ),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/fch_issu1 ),
        .I5(fch_heir_nir_i_3_n_0),
        .O(\fch/fctl/fch_heir_nir_t ));
  LUT3 #(
    .INIT(8'h08)) 
    fch_heir_nir_i_2
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\nir_id[24]_i_6_n_0 ),
        .I2(\nir_id[24]_i_4_n_0 ),
        .O(fch_heir_nir_i_2_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_heir_nir_i_3
       (.I0(ctl_fetch_lng0),
        .I1(ctl_fetch_lng1),
        .O(fch_heir_nir_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    fch_heir_nir_i_4
       (.I0(fch_heir_nir_i_6_n_0),
        .I1(\ccmd[1]_INST_0_i_16_n_0 ),
        .I2(fch_heir_nir_i_7_n_0),
        .I3(\fch/ir0 [7]),
        .I4(\rgf/sreg/sr [9]),
        .I5(\fch/ir0 [15]),
        .O(ctl_fetch_lng0));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    fch_heir_nir_i_5
       (.I0(\rgf/sreg/sr [9]),
        .I1(\fch/ir1 [7]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\ctl1/stat_reg_n_0_[2] ),
        .I4(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I5(fch_heir_nir_i_8_n_0),
        .O(ctl_fetch_lng1));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    fch_heir_nir_i_6
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [10]),
        .O(fch_heir_nir_i_6_n_0));
  LUT4 #(
    .INIT(16'h0100)) 
    fch_heir_nir_i_7
       (.I0(stat[1]),
        .I1(stat[2]),
        .I2(stat[0]),
        .I3(\fch/ir0 [11]),
        .O(fch_heir_nir_i_7_n_0));
  LUT6 #(
    .INIT(64'hFDFFFFFFFFFFFFFF)) 
    fch_heir_nir_i_8
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [15]),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I4(\bdatw[31]_INST_0_i_151_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_23_n_0 ),
        .O(fch_heir_nir_i_8_n_0));
  LUT4 #(
    .INIT(16'hFB08)) 
    \fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(fch_irq_req),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .I3(fch_irq_lev[0]),
        .O(\fch_irq_lev[0]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hFB08)) 
    \fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(fch_irq_req),
        .I2(\fch_irq_lev[1]_i_2_n_0 ),
        .I3(fch_irq_lev[1]),
        .O(\fch_irq_lev[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h7FFF00007FFF7FFF)) 
    \fch_irq_lev[1]_i_2 
       (.I0(\rgf_selc0_wb[1]_i_12_n_0 ),
        .I1(\fch/ir0 [0]),
        .I2(\fch_irq_lev[1]_i_3_n_0 ),
        .I3(\fch_irq_lev[1]_i_4_n_0 ),
        .I4(\fch_irq_lev[1]_i_5_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\fch_irq_lev[1]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fch_irq_lev[1]_i_3 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [6]),
        .O(\fch_irq_lev[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \fch_irq_lev[1]_i_4 
       (.I0(\fch_irq_lev[1]_i_6_n_0 ),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [2]),
        .I3(brdy),
        .I4(fch_irq_req),
        .I5(\stat[2]_i_4_n_0 ),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF7FF)) 
    \fch_irq_lev[1]_i_5 
       (.I0(\niss_dsp_a1[32]_INST_0_i_24_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\fch_irq_lev[1]_i_7_n_0 ),
        .I3(\fch_irq_lev[1]_i_8_n_0 ),
        .I4(\fch/ir1 [8]),
        .I5(\fch_irq_lev[1]_i_9_n_0 ),
        .O(\fch_irq_lev[1]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fch_irq_lev[1]_i_6 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [7]),
        .O(\fch_irq_lev[1]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \fch_irq_lev[1]_i_7 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [11]),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\ctl1/stat_reg_n_0_[2] ),
        .O(\fch_irq_lev[1]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fch_irq_lev[1]_i_8 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [5]),
        .O(\fch_irq_lev[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \fch_irq_lev[1]_i_9 
       (.I0(\fch/ir1 [6]),
        .I1(fch_irq_req),
        .I2(\bdatw[9]_INST_0_i_10_n_0 ),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [3]),
        .I5(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .O(\fch_irq_lev[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h20F20000)) 
    fch_irq_req_fl_i_1
       (.I0(\rgf/sreg/sr [2]),
        .I1(irq_lev[0]),
        .I2(\rgf/sreg/sr [3]),
        .I3(irq_lev[1]),
        .I4(irq),
        .O(fch_irq_req));
  LUT3 #(
    .INIT(8'hB8)) 
    fch_issu1_fl_i_1
       (.I0(\fch/fch_issu1 ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_issu1_fl ),
        .O(\fch/fch_issu1_ir ));
  LUT6 #(
    .INIT(64'h0A02AA82A080AA82)) 
    fch_issu1_inferred_i_1
       (.I0(fch_issu1_inferred_i_2_n_0),
        .I1(fch_issu1_inferred_i_3_n_0),
        .I2(fch_issu1_inferred_i_4_n_0),
        .I3(fch_issu1_inferred_i_5_n_0),
        .I4(fch_issu1_inferred_i_6_n_0),
        .I5(fch_issu1_inferred_i_7_n_0),
        .O(\fch/fch_issu1 ));
  LUT6 #(
    .INIT(64'hEFFFEFEEEFFFEFFF)) 
    fch_issu1_inferred_i_10
       (.I0(fch_issu1_inferred_i_35_n_0),
        .I1(\rgf/sreg/sr [9]),
        .I2(fch_issu1_inferred_i_36_n_0),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_37_n_0),
        .I5(fch_issu1_inferred_i_38_n_0),
        .O(fch_issu1_inferred_i_10_n_0));
  LUT6 #(
    .INIT(64'h0200002002220000)) 
    fch_issu1_inferred_i_100
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[6]),
        .I3(fdat[9]),
        .I4(fdat[8]),
        .I5(fdat[7]),
        .O(fch_issu1_inferred_i_100_n_0));
  LUT5 #(
    .INIT(32'hF000B030)) 
    fch_issu1_inferred_i_101
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[10]),
        .I3(fdat[6]),
        .I4(fdat[9]),
        .O(fch_issu1_inferred_i_101_n_0));
  LUT6 #(
    .INIT(64'hDFDDFDFFFFFFFDFD)) 
    fch_issu1_inferred_i_102
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[5]),
        .I3(fdat[3]),
        .I4(fdat[4]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_102_n_0));
  LUT6 #(
    .INIT(64'h4B00EB00FFFFFFFF)) 
    fch_issu1_inferred_i_103
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_103_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    fch_issu1_inferred_i_104
       (.I0(fdat[4]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .O(fch_issu1_inferred_i_104_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_105
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .O(fch_issu1_inferred_i_105_n_0));
  LUT6 #(
    .INIT(64'h00000000D755D555)) 
    fch_issu1_inferred_i_106
       (.I0(fdat[31]),
        .I1(fdat[28]),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .I4(fdat[27]),
        .I5(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_106_n_0));
  LUT5 #(
    .INIT(32'hA8AAAAAA)) 
    fch_issu1_inferred_i_107
       (.I0(fch_issu1_inferred_i_157_n_0),
        .I1(fdat[19]),
        .I2(fdat[27]),
        .I3(fdat[28]),
        .I4(fch_issu1_inferred_i_94_n_0),
        .O(fch_issu1_inferred_i_107_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_108
       (.I0(fdat[30]),
        .I1(fdat[29]),
        .O(fch_issu1_inferred_i_108_n_0));
  LUT6 #(
    .INIT(64'h2AAAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_109
       (.I0(fch_issu1_inferred_i_158_n_0),
        .I1(fdat[8]),
        .I2(fdat[0]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .I5(fch_issu1_inferred_i_159_n_0),
        .O(fch_issu1_inferred_i_109_n_0));
  LUT6 #(
    .INIT(64'h00E0FFEFFFEFFFEF)) 
    fch_issu1_inferred_i_11
       (.I0(fch_issu1_inferred_i_39_n_0),
        .I1(fch_issu1_inferred_i_40_n_0),
        .I2(\fch/stat [1]),
        .I3(\fch/stat [0]),
        .I4(fch_issu1_inferred_i_41_n_0),
        .I5(fch_issu1_inferred_i_42_n_0),
        .O(fch_issu1_inferred_i_11_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    fch_issu1_inferred_i_110
       (.I0(fdat[31]),
        .I1(fdat[29]),
        .I2(fdat[30]),
        .O(fch_issu1_inferred_i_110_n_0));
  LUT5 #(
    .INIT(32'hAC00A000)) 
    fch_issu1_inferred_i_111
       (.I0(fch_issu1_inferred_i_160_n_0),
        .I1(fdat[19]),
        .I2(fdat[27]),
        .I3(fdat[28]),
        .I4(fch_issu1_inferred_i_161_n_0),
        .O(fch_issu1_inferred_i_111_n_0));
  LUT6 #(
    .INIT(64'h0888008888888888)) 
    fch_issu1_inferred_i_112
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_162_n_0),
        .I2(fdat[14]),
        .I3(fdat[13]),
        .I4(fdat[11]),
        .I5(fdat[12]),
        .O(fch_issu1_inferred_i_112_n_0));
  LUT6 #(
    .INIT(64'h0000005D00000000)) 
    fch_issu1_inferred_i_113
       (.I0(\nir_id[21]_i_9_n_0 ),
        .I1(fch_issu1_inferred_i_163_n_0),
        .I2(fch_issu1_inferred_i_164_n_0),
        .I3(fch_issu1_inferred_i_165_n_0),
        .I4(fch_issu1_inferred_i_100_n_0),
        .I5(fch_issu1_inferred_i_93_n_0),
        .O(fch_issu1_inferred_i_113_n_0));
  LUT6 #(
    .INIT(64'h0000000003332333)) 
    fch_issu1_inferred_i_114
       (.I0(fdat[11]),
        .I1(\fch/fadr_1_fl ),
        .I2(fdat[12]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_114_n_0));
  LUT5 #(
    .INIT(32'h0000007F)) 
    fch_issu1_inferred_i_115
       (.I0(\nir_id[21]_i_8_n_0 ),
        .I1(\nir_id[21]_i_7_n_0 ),
        .I2(fch_issu1_inferred_i_166_n_0),
        .I3(fdat[14]),
        .I4(fdat[15]),
        .O(fch_issu1_inferred_i_115_n_0));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    fch_issu1_inferred_i_116
       (.I0(fch_issu1_inferred_i_167_n_0),
        .I1(fch_issu1_inferred_i_168_n_0),
        .I2(fch_issu1_inferred_i_169_n_0),
        .I3(fch_issu1_inferred_i_170_n_0),
        .I4(fdat[28]),
        .I5(fdat[29]),
        .O(fch_issu1_inferred_i_116_n_0));
  LUT6 #(
    .INIT(64'h5555555504000000)) 
    fch_issu1_inferred_i_117
       (.I0(fdat[31]),
        .I1(\ir0_id_fl[21]_i_11_n_0 ),
        .I2(fch_issu1_inferred_i_171_n_0),
        .I3(fdat[17]),
        .I4(\ir0_id_fl[21]_i_5_n_0 ),
        .I5(fdat[30]),
        .O(fch_issu1_inferred_i_117_n_0));
  LUT6 #(
    .INIT(64'h0000000020002333)) 
    fch_issu1_inferred_i_118
       (.I0(fch_issu1_inferred_i_172_n_0),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fdat[27]),
        .I4(fdat[20]),
        .I5(fch_issu1_inferred_i_46_n_0),
        .O(fch_issu1_inferred_i_118_n_0));
  LUT6 #(
    .INIT(64'h440F440F0000000F)) 
    fch_issu1_inferred_i_119
       (.I0(fdat[2]),
        .I1(fch_issu1_inferred_i_159_n_0),
        .I2(fdat[5]),
        .I3(fdat[9]),
        .I4(fch_issu1_inferred_i_105_n_0),
        .I5(fdat[8]),
        .O(fch_issu1_inferred_i_119_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    fch_issu1_inferred_i_12
       (.I0(fch_issu1_inferred_i_21_n_0),
        .I1(fch_issu1_inferred_i_33_n_0),
        .I2(fch_issu1_inferred_i_43_n_0),
        .I3(fch_issu1_inferred_i_24_n_0),
        .I4(fch_issu1_inferred_i_44_n_0),
        .I5(fch_issu1_inferred_i_26_n_0),
        .O(fch_issu1_inferred_i_12_n_0));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFFBAAAA)) 
    fch_issu1_inferred_i_120
       (.I0(fch_issu1_inferred_i_115_n_0),
        .I1(fch_issu1_inferred_i_173_n_0),
        .I2(\nir_id[21]_i_6_n_0 ),
        .I3(fdat[10]),
        .I4(fdat[15]),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_120_n_0));
  LUT6 #(
    .INIT(64'hBFBFFFBFFFBFFFBF)) 
    fch_issu1_inferred_i_121
       (.I0(fch_issu1_inferred_i_55_n_0),
        .I1(fdat[29]),
        .I2(fdat[28]),
        .I3(fdat[21]),
        .I4(fdat[27]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_121_n_0));
  LUT6 #(
    .INIT(64'h55550100FFFFFFFF)) 
    fch_issu1_inferred_i_122
       (.I0(fch_issu1_inferred_i_174_n_0),
        .I1(fdat[18]),
        .I2(fch_issu1_inferred_i_99_n_0),
        .I3(fch_issu1_inferred_i_175_n_0),
        .I4(fch_issu1_inferred_i_176_n_0),
        .I5(fch_issu1_inferred_i_48_n_0),
        .O(fch_issu1_inferred_i_122_n_0));
  LUT6 #(
    .INIT(64'h0000000020002333)) 
    fch_issu1_inferred_i_123
       (.I0(fch_issu1_inferred_i_177_n_0),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fdat[27]),
        .I4(fdat[21]),
        .I5(fch_issu1_inferred_i_46_n_0),
        .O(fch_issu1_inferred_i_123_n_0));
  LUT6 #(
    .INIT(64'hAAAAFFBEAAAAAAAA)) 
    fch_issu1_inferred_i_124
       (.I0(fch_issu1_inferred_i_110_n_0),
        .I1(fdat[17]),
        .I2(fdat[19]),
        .I3(fdat[16]),
        .I4(fch_issu1_inferred_i_178_n_0),
        .I5(\ir0_id_fl[20]_i_7_n_0 ),
        .O(fch_issu1_inferred_i_124_n_0));
  LUT6 #(
    .INIT(64'hA008AA08AAA8AAA8)) 
    fch_issu1_inferred_i_125
       (.I0(fdat[26]),
        .I1(fdat[16]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_125_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAA00200000)) 
    fch_issu1_inferred_i_126
       (.I0(fch_issu1_inferred_i_179_n_0),
        .I1(fdat[24]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_126_n_0));
  LUT6 #(
    .INIT(64'h0001555504415555)) 
    fch_issu1_inferred_i_127
       (.I0(fch_issu1_inferred_i_180_n_0),
        .I1(fch_issu1_inferred_i_149_n_0),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fdat[19]),
        .O(fch_issu1_inferred_i_127_n_0));
  LUT6 #(
    .INIT(64'h7777FF77F7777777)) 
    fch_issu1_inferred_i_128
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .I2(fdat[16]),
        .I3(fdat[24]),
        .I4(fdat[26]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_128_n_0));
  LUT6 #(
    .INIT(64'hA2A0AAA8AAA8AAA8)) 
    fch_issu1_inferred_i_129
       (.I0(fdat[26]),
        .I1(fdat[24]),
        .I2(fdat[25]),
        .I3(fdat[18]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_129_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_13
       (.I0(\fch/stat [1]),
        .I1(\fch/stat [0]),
        .O(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'hAAAAFAFAEFEAAAAA)) 
    fch_issu1_inferred_i_130
       (.I0(fch_issu1_inferred_i_181_n_0),
        .I1(fdat[18]),
        .I2(fdat[24]),
        .I3(fdat[23]),
        .I4(fdat[26]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_130_n_0));
  LUT6 #(
    .INIT(64'hAA0A2AAAAA0A2A00)) 
    fch_issu1_inferred_i_131
       (.I0(fdat[26]),
        .I1(fdat[22]),
        .I2(fdat[23]),
        .I3(fdat[24]),
        .I4(fdat[25]),
        .I5(fdat[17]),
        .O(fch_issu1_inferred_i_131_n_0));
  LUT6 #(
    .INIT(64'hFFFFAEAAFAAAFAAA)) 
    fch_issu1_inferred_i_132
       (.I0(fch_issu1_inferred_i_181_n_0),
        .I1(fdat[17]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fch_issu1_inferred_i_182_n_0),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_132_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_133
       (.I0(fdat[20]),
        .I1(fdat[19]),
        .O(fch_issu1_inferred_i_133_n_0));
  LUT6 #(
    .INIT(64'h0000000057755557)) 
    fch_issu1_inferred_i_134
       (.I0(fch_issu1_inferred_i_48_n_0),
        .I1(fdat[22]),
        .I2(fdat[21]),
        .I3(fdat[20]),
        .I4(fdat[23]),
        .I5(fch_issu1_inferred_i_183_n_0),
        .O(fch_issu1_inferred_i_134_n_0));
  LUT6 #(
    .INIT(64'h000000007F000000)) 
    fch_issu1_inferred_i_135
       (.I0(fdat[24]),
        .I1(fdat[26]),
        .I2(fdat[28]),
        .I3(fdat[30]),
        .I4(fdat[29]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_135_n_0));
  LUT6 #(
    .INIT(64'hCFCCEEEEEEEEEEFF)) 
    fch_issu1_inferred_i_136
       (.I0(fdat[15]),
        .I1(fch_issu1_inferred_i_184_n_0),
        .I2(fch_issu1_inferred_i_185_n_0),
        .I3(fdat[12]),
        .I4(fdat[13]),
        .I5(fdat[14]),
        .O(fch_issu1_inferred_i_136_n_0));
  LUT6 #(
    .INIT(64'hFFFFFF7FFFFFFFFF)) 
    fch_issu1_inferred_i_137
       (.I0(fdat[12]),
        .I1(fdat[10]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_137_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_138
       (.I0(fdat[23]),
        .I1(fdat[22]),
        .O(fch_issu1_inferred_i_138_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    fch_issu1_inferred_i_139
       (.I0(fdat[24]),
        .I1(fdat[25]),
        .O(fch_issu1_inferred_i_139_n_0));
  LUT6 #(
    .INIT(64'h3111133131311111)) 
    fch_issu1_inferred_i_14
       (.I0(fdat[31]),
        .I1(fch_issu1_inferred_i_45_n_0),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .I4(fdat[28]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_14_n_0));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    fch_issu1_inferred_i_140
       (.I0(fch_issu1_inferred_i_180_n_0),
        .I1(fdat[24]),
        .I2(fch_issu1_inferred_i_149_n_0),
        .I3(fdat[31]),
        .I4(fdat[19]),
        .I5(fdat[22]),
        .O(fch_issu1_inferred_i_140_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAABBBF)) 
    fch_issu1_inferred_i_141
       (.I0(fdat[31]),
        .I1(fdat[26]),
        .I2(fch_issu1_inferred_i_149_n_0),
        .I3(fdat[23]),
        .I4(fdat[22]),
        .I5(fch_issu1_inferred_i_186_n_0),
        .O(fch_issu1_inferred_i_141_n_0));
  LUT6 #(
    .INIT(64'h0000808088080800)) 
    fch_issu1_inferred_i_142
       (.I0(fdat[26]),
        .I1(fdat[25]),
        .I2(fdat[20]),
        .I3(fdat[23]),
        .I4(fdat[22]),
        .I5(fdat[21]),
        .O(fch_issu1_inferred_i_142_n_0));
  LUT6 #(
    .INIT(64'hF777F7F777777777)) 
    fch_issu1_inferred_i_143
       (.I0(fdat[29]),
        .I1(fdat[30]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fch_issu1_inferred_i_179_n_0),
        .O(fch_issu1_inferred_i_143_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAEFAAAAAA)) 
    fch_issu1_inferred_i_144
       (.I0(\nir_id[13]_i_5_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[8]),
        .I3(fdat[7]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_144_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF380E0000)) 
    fch_issu1_inferred_i_145
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(\nir_id[19]_i_7_n_0 ),
        .I5(fch_issu1_inferred_i_187_n_0),
        .O(fch_issu1_inferred_i_145_n_0));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    fch_issu1_inferred_i_146
       (.I0(\nir_id[20]_i_8_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[3]),
        .I4(fdat[8]),
        .I5(fdat[15]),
        .O(fch_issu1_inferred_i_146_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF19FF0000)) 
    fch_issu1_inferred_i_147
       (.I0(fdat[3]),
        .I1(fdat[1]),
        .I2(fdat[0]),
        .I3(fch_issu1_inferred_i_153_n_0),
        .I4(fch_issu1_inferred_i_152_n_0),
        .I5(fch_issu1_inferred_i_188_n_0),
        .O(fch_issu1_inferred_i_147_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFBD)) 
    fch_issu1_inferred_i_148
       (.I0(fdat[16]),
        .I1(fdat[19]),
        .I2(fdat[17]),
        .I3(fdat[30]),
        .I4(fdat[29]),
        .I5(fdat[28]),
        .O(fch_issu1_inferred_i_148_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_149
       (.I0(fdat[21]),
        .I1(fdat[20]),
        .O(fch_issu1_inferred_i_149_n_0));
  LUT6 #(
    .INIT(64'h0000000000001101)) 
    fch_issu1_inferred_i_15
       (.I0(fch_issu1_inferred_i_46_n_0),
        .I1(fch_issu1_inferred_i_47_n_0),
        .I2(fch_issu1_inferred_i_48_n_0),
        .I3(fch_issu1_inferred_i_49_n_0),
        .I4(fdat[31]),
        .I5(fch_issu1_inferred_i_50_n_0),
        .O(fch_issu1_inferred_i_15_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_150
       (.I0(fdat[23]),
        .I1(fdat[22]),
        .O(fch_issu1_inferred_i_150_n_0));
  LUT6 #(
    .INIT(64'h0000000000000888)) 
    fch_issu1_inferred_i_151
       (.I0(fdat[9]),
        .I1(\nir_id[21]_i_6_n_0 ),
        .I2(fdat[10]),
        .I3(\nir_id[18]_i_7_n_0 ),
        .I4(fdat[8]),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_151_n_0));
  LUT3 #(
    .INIT(8'h01)) 
    fch_issu1_inferred_i_152
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .O(fch_issu1_inferred_i_152_n_0));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    fch_issu1_inferred_i_153
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[9]),
        .I3(fdat[7]),
        .I4(fdat[6]),
        .I5(\nir_id[21]_i_10_n_0 ),
        .O(fch_issu1_inferred_i_153_n_0));
  LUT6 #(
    .INIT(64'h3030000230300000)) 
    fch_issu1_inferred_i_154
       (.I0(fch_issu1_inferred_i_189_n_0),
        .I1(fch_issu1_inferred_i_190_n_0),
        .I2(fdat[28]),
        .I3(fdat[29]),
        .I4(fdat[23]),
        .I5(fch_issu1_inferred_i_149_n_0),
        .O(fch_issu1_inferred_i_154_n_0));
  LUT6 #(
    .INIT(64'h28FFFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_155
       (.I0(fdat[22]),
        .I1(fdat[19]),
        .I2(fdat[21]),
        .I3(fdat[24]),
        .I4(fdat[28]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_155_n_0));
  LUT5 #(
    .INIT(32'hC70FF73F)) 
    fch_issu1_inferred_i_156
       (.I0(fdat[25]),
        .I1(fdat[20]),
        .I2(fdat[22]),
        .I3(fdat[21]),
        .I4(fdat[23]),
        .O(fch_issu1_inferred_i_156_n_0));
  LUT6 #(
    .INIT(64'hFFD0FF00FFFFFF00)) 
    fch_issu1_inferred_i_157
       (.I0(fch_issu1_inferred_i_191_n_0),
        .I1(fdat[16]),
        .I2(fdat[25]),
        .I3(fch_issu1_inferred_i_192_n_0),
        .I4(fdat[26]),
        .I5(fch_issu1_inferred_i_49_n_0),
        .O(fch_issu1_inferred_i_157_n_0));
  LUT6 #(
    .INIT(64'hFF040A62FFFFFFFF)) 
    fch_issu1_inferred_i_158
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[3]),
        .O(fch_issu1_inferred_i_158_n_0));
  LUT5 #(
    .INIT(32'h4B83EBA9)) 
    fch_issu1_inferred_i_159
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .I3(fdat[7]),
        .I4(fdat[3]),
        .O(fch_issu1_inferred_i_159_n_0));
  LUT4 #(
    .INIT(16'h0220)) 
    fch_issu1_inferred_i_16
       (.I0(fdat[30]),
        .I1(fdat[29]),
        .I2(fdat[28]),
        .I3(fdat[27]),
        .O(fch_issu1_inferred_i_16_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAEAAAAAAA)) 
    fch_issu1_inferred_i_160
       (.I0(fch_issu1_inferred_i_193_n_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fdat[16]),
        .I5(fch_issu1_inferred_i_194_n_0),
        .O(fch_issu1_inferred_i_160_n_0));
  LUT5 #(
    .INIT(32'hF000D050)) 
    fch_issu1_inferred_i_161
       (.I0(fdat[24]),
        .I1(fdat[23]),
        .I2(fdat[26]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .O(fch_issu1_inferred_i_161_n_0));
  LUT4 #(
    .INIT(16'h00A2)) 
    fch_issu1_inferred_i_162
       (.I0(fdat[8]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_162_n_0));
  LUT6 #(
    .INIT(64'h7FF777FDF55555FF)) 
    fch_issu1_inferred_i_163
       (.I0(fdat[9]),
        .I1(fdat[3]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_163_n_0));
  LUT6 #(
    .INIT(64'hE2EEE2EEE2CCE2EE)) 
    fch_issu1_inferred_i_164
       (.I0(fdat[4]),
        .I1(fdat[9]),
        .I2(fdat[1]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_164_n_0));
  LUT6 #(
    .INIT(64'hAAAAFEAEEEEEFEAE)) 
    fch_issu1_inferred_i_165
       (.I0(fch_issu1_inferred_i_91_n_0),
        .I1(fdat[4]),
        .I2(fch_issu1_inferred_i_195_n_0),
        .I3(fch_issu1_inferred_i_196_n_0),
        .I4(fdat[11]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_165_n_0));
  LUT5 #(
    .INIT(32'h00000020)) 
    fch_issu1_inferred_i_166
       (.I0(fdat[0]),
        .I1(fdat[3]),
        .I2(fdat[1]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .O(fch_issu1_inferred_i_166_n_0));
  LUT6 #(
    .INIT(64'h55551055FFFFFFFF)) 
    fch_issu1_inferred_i_167
       (.I0(fch_issu1_inferred_i_197_n_0),
        .I1(fch_issu1_inferred_i_99_n_0),
        .I2(fch_issu1_inferred_i_175_n_0),
        .I3(fdat[25]),
        .I4(fch_issu1_inferred_i_198_n_0),
        .I5(fch_issu1_inferred_i_48_n_0),
        .O(fch_issu1_inferred_i_167_n_0));
  LUT6 #(
    .INIT(64'h0200002002220000)) 
    fch_issu1_inferred_i_168
       (.I0(fdat[27]),
        .I1(fdat[26]),
        .I2(fdat[22]),
        .I3(fdat[25]),
        .I4(fdat[24]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_168_n_0));
  LUT6 #(
    .INIT(64'h00FFF7F70000A2A2)) 
    fch_issu1_inferred_i_169
       (.I0(fch_issu1_inferred_i_199_n_0),
        .I1(fdat[23]),
        .I2(fdat[24]),
        .I3(fdat[26]),
        .I4(fdat[27]),
        .I5(fdat[20]),
        .O(fch_issu1_inferred_i_169_n_0));
  LUT5 #(
    .INIT(32'h22AAA2AA)) 
    fch_issu1_inferred_i_17
       (.I0(fdat[31]),
        .I1(fdat[28]),
        .I2(fdat[27]),
        .I3(fdat[29]),
        .I4(fdat[30]),
        .O(fch_issu1_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'h0010101055555555)) 
    fch_issu1_inferred_i_170
       (.I0(fdat[27]),
        .I1(fdat[25]),
        .I2(fdat[24]),
        .I3(fdat[23]),
        .I4(fdat[22]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_170_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFDFF)) 
    fch_issu1_inferred_i_171
       (.I0(fch_issu1_inferred_i_149_n_0),
        .I1(fdat[22]),
        .I2(fdat[19]),
        .I3(fdat[16]),
        .I4(fdat[29]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_171_n_0));
  LUT6 #(
    .INIT(64'h03A300A003A303A3)) 
    fch_issu1_inferred_i_172
       (.I0(fch_issu1_inferred_i_191_n_0),
        .I1(fdat[20]),
        .I2(fdat[25]),
        .I3(fdat[17]),
        .I4(fdat[24]),
        .I5(fch_issu1_inferred_i_150_n_0),
        .O(fch_issu1_inferred_i_172_n_0));
  LUT5 #(
    .INIT(32'h55555155)) 
    fch_issu1_inferred_i_173
       (.I0(\fch/fadr_1_fl ),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .O(fch_issu1_inferred_i_173_n_0));
  LUT5 #(
    .INIT(32'h00FF0010)) 
    fch_issu1_inferred_i_174
       (.I0(fdat[24]),
        .I1(fdat[22]),
        .I2(fdat[23]),
        .I3(fdat[25]),
        .I4(fdat[21]),
        .O(fch_issu1_inferred_i_174_n_0));
  LUT4 #(
    .INIT(16'h9EFF)) 
    fch_issu1_inferred_i_175
       (.I0(fdat[21]),
        .I1(fdat[20]),
        .I2(fdat[19]),
        .I3(fdat[22]),
        .O(fch_issu1_inferred_i_175_n_0));
  LUT6 #(
    .INIT(64'h2F2F2F2F2F0F0F2F)) 
    fch_issu1_inferred_i_176
       (.I0(fch_issu1_inferred_i_200_n_0),
        .I1(fdat[18]),
        .I2(fdat[25]),
        .I3(fdat[20]),
        .I4(fdat[21]),
        .I5(fdat[22]),
        .O(fch_issu1_inferred_i_176_n_0));
  LUT6 #(
    .INIT(64'h202F2020202F202F)) 
    fch_issu1_inferred_i_177
       (.I0(fch_issu1_inferred_i_191_n_0),
        .I1(fdat[18]),
        .I2(fdat[25]),
        .I3(fdat[21]),
        .I4(fdat[24]),
        .I5(fch_issu1_inferred_i_150_n_0),
        .O(fch_issu1_inferred_i_177_n_0));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    fch_issu1_inferred_i_178
       (.I0(fdat[28]),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fdat[27]),
        .I4(fdat[30]),
        .O(fch_issu1_inferred_i_178_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_179
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .O(fch_issu1_inferred_i_179_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF200)) 
    fch_issu1_inferred_i_18
       (.I0(fch_issu1_inferred_i_51_n_0),
        .I1(fch_issu1_inferred_i_52_n_0),
        .I2(fch_issu1_inferred_i_53_n_0),
        .I3(fch_issu1_inferred_i_48_n_0),
        .I4(fch_issu1_inferred_i_54_n_0),
        .I5(fch_issu1_inferred_i_55_n_0),
        .O(fch_issu1_inferred_i_18_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_180
       (.I0(fdat[25]),
        .I1(fdat[26]),
        .O(fch_issu1_inferred_i_180_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_181
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .O(fch_issu1_inferred_i_181_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFA28A)) 
    fch_issu1_inferred_i_182
       (.I0(fdat[22]),
        .I1(fdat[20]),
        .I2(fdat[19]),
        .I3(fdat[21]),
        .I4(fch_issu1_inferred_i_99_n_0),
        .I5(fch_issu1_inferred_i_201_n_0),
        .O(fch_issu1_inferred_i_182_n_0));
  LUT6 #(
    .INIT(64'hABEBBFFFAFEFBFFF)) 
    fch_issu1_inferred_i_183
       (.I0(fdat[31]),
        .I1(fdat[24]),
        .I2(fdat[25]),
        .I3(fdat[26]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_183_n_0));
  LUT6 #(
    .INIT(64'h0000000005775577)) 
    fch_issu1_inferred_i_184
       (.I0(fdat[11]),
        .I1(fdat[15]),
        .I2(fdat[8]),
        .I3(fdat[12]),
        .I4(fdat[10]),
        .I5(\nir_id[13]_i_5_n_0 ),
        .O(fch_issu1_inferred_i_184_n_0));
  LUT6 #(
    .INIT(64'h02200002AAAAAAAA)) 
    fch_issu1_inferred_i_185
       (.I0(fch_issu1_inferred_i_202_n_0),
        .I1(fdat[6]),
        .I2(fdat[5]),
        .I3(fdat[4]),
        .I4(fdat[7]),
        .I5(\nir_id[21]_i_9_n_0 ),
        .O(fch_issu1_inferred_i_185_n_0));
  LUT6 #(
    .INIT(64'h5ADADEDEA5E5FFFF)) 
    fch_issu1_inferred_i_186
       (.I0(fdat[26]),
        .I1(fch_issu1_inferred_i_179_n_0),
        .I2(fdat[24]),
        .I3(fdat[22]),
        .I4(fdat[23]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_186_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF00FF2F)) 
    fch_issu1_inferred_i_187
       (.I0(\nir_id[24]_i_22_n_0 ),
        .I1(fdat[7]),
        .I2(fdat[10]),
        .I3(fdat[15]),
        .I4(fdat[6]),
        .I5(fch_issu1_inferred_i_203_n_0),
        .O(fch_issu1_inferred_i_187_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF550015)) 
    fch_issu1_inferred_i_188
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fch_issu1_inferred_i_204_n_0),
        .I3(\nir_id[13]_i_5_n_0 ),
        .I4(fdat[15]),
        .I5(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_188_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    fch_issu1_inferred_i_189
       (.I0(fdat[18]),
        .I1(fdat[25]),
        .O(fch_issu1_inferred_i_189_n_0));
  LUT6 #(
    .INIT(64'hFFFBFFFBFFFFFFFB)) 
    fch_issu1_inferred_i_19
       (.I0(\fch/fadr_1_fl ),
        .I1(fdat[14]),
        .I2(fdat[15]),
        .I3(fch_issu1_inferred_i_56_n_0),
        .I4(\nir_id[21]_i_9_n_0 ),
        .I5(fch_issu1_inferred_i_57_n_0),
        .O(fch_issu1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEFE)) 
    fch_issu1_inferred_i_190
       (.I0(fdat[22]),
        .I1(fdat[24]),
        .I2(fdat[23]),
        .I3(fdat[25]),
        .I4(fdat[26]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_190_n_0));
  LUT6 #(
    .INIT(64'h88C0C0C0488000C4)) 
    fch_issu1_inferred_i_191
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[22]),
        .I3(fdat[21]),
        .I4(fdat[20]),
        .I5(fdat[19]),
        .O(fch_issu1_inferred_i_191_n_0));
  LUT6 #(
    .INIT(64'h7F55FFFFFFFFFFFF)) 
    fch_issu1_inferred_i_192
       (.I0(fch_issu1_inferred_i_95_n_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fdat[19]),
        .I4(fdat[28]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_192_n_0));
  LUT6 #(
    .INIT(64'h0000AAA2AA0A828A)) 
    fch_issu1_inferred_i_193
       (.I0(fdat[19]),
        .I1(fdat[23]),
        .I2(fdat[24]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[26]),
        .O(fch_issu1_inferred_i_193_n_0));
  LUT5 #(
    .INIT(32'h9715F052)) 
    fch_issu1_inferred_i_194
       (.I0(fdat[22]),
        .I1(fdat[23]),
        .I2(fdat[21]),
        .I3(fdat[19]),
        .I4(fdat[20]),
        .O(fch_issu1_inferred_i_194_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_195
       (.I0(fdat[9]),
        .I1(fdat[6]),
        .O(fch_issu1_inferred_i_195_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_196
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .O(fch_issu1_inferred_i_196_n_0));
  LUT6 #(
    .INIT(64'hB8B8B888B8B8B8B8)) 
    fch_issu1_inferred_i_197
       (.I0(fdat[17]),
        .I1(fdat[25]),
        .I2(fdat[20]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_197_n_0));
  LUT6 #(
    .INIT(64'h40C0C0004000C0C0)) 
    fch_issu1_inferred_i_198
       (.I0(fdat[19]),
        .I1(fdat[24]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[21]),
        .I5(fdat[20]),
        .O(fch_issu1_inferred_i_198_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    fch_issu1_inferred_i_199
       (.I0(fdat[25]),
        .I1(fdat[22]),
        .O(fch_issu1_inferred_i_199_n_0));
  LUT6 #(
    .INIT(64'h0C080C080C000008)) 
    fch_issu1_inferred_i_2
       (.I0(fch_issu1_inferred_i_8_n_0),
        .I1(fch_issu1_inferred_i_9_n_0),
        .I2(fch_issu1_inferred_i_10_n_0),
        .I3(fch_issu1_inferred_i_3_n_0),
        .I4(fch_issu1_inferred_i_11_n_0),
        .I5(fch_issu1_inferred_i_12_n_0),
        .O(fch_issu1_inferred_i_2_n_0));
  LUT6 #(
    .INIT(64'h00002AA2000002AA)) 
    fch_issu1_inferred_i_20
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .I2(fdat[13]),
        .I3(fdat[12]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[11]),
        .O(fch_issu1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'h08888888)) 
    fch_issu1_inferred_i_200
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[21]),
        .I3(fdat[22]),
        .I4(fdat[19]),
        .O(fch_issu1_inferred_i_200_n_0));
  LUT6 #(
    .INIT(64'h08880880FFFFFFFF)) 
    fch_issu1_inferred_i_201
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[22]),
        .I3(fdat[21]),
        .I4(fdat[20]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_201_n_0));
  LUT6 #(
    .INIT(64'h0F0C0800000C0800)) 
    fch_issu1_inferred_i_202
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .I2(fdat[15]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_202_n_0));
  LUT6 #(
    .INIT(64'h4CFFFF55FF445DFF)) 
    fch_issu1_inferred_i_203
       (.I0(fdat[7]),
        .I1(\nir_id[14]_i_9_n_0 ),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_203_n_0));
  LUT2 #(
    .INIT(4'h6)) 
    fch_issu1_inferred_i_204
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(fch_issu1_inferred_i_204_n_0));
  LUT6 #(
    .INIT(64'h0D0D000F0D0D0D0D)) 
    fch_issu1_inferred_i_21
       (.I0(\fch/fadr_1_fl ),
        .I1(\nir_id[16]_i_2_n_0 ),
        .I2(fch_issu1_inferred_i_58_n_0),
        .I3(\fch/nir_id [16]),
        .I4(\fch/stat [0]),
        .I5(\fch/stat [1]),
        .O(fch_issu1_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFFDF)) 
    fch_issu1_inferred_i_22
       (.I0(fdat[14]),
        .I1(fdat[15]),
        .I2(fdat[13]),
        .I3(fch_issu1_inferred_i_45_n_0),
        .I4(fch_issu1_inferred_i_59_n_0),
        .I5(fch_issu1_inferred_i_60_n_0),
        .O(fch_issu1_inferred_i_22_n_0));
  MUXF7 fch_issu1_inferred_i_23
       (.I0(fch_issu1_inferred_i_61_n_0),
        .I1(fch_issu1_inferred_i_62_n_0),
        .O(fch_issu1_inferred_i_23_n_0),
        .S(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'h00000000DD0FDDDD)) 
    fch_issu1_inferred_i_24
       (.I0(\fch/fadr_1_fl ),
        .I1(\nir_id[17]_i_2_n_0 ),
        .I2(\fch/nir_id [17]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fch_issu1_inferred_i_63_n_0),
        .O(fch_issu1_inferred_i_24_n_0));
  MUXF7 fch_issu1_inferred_i_25
       (.I0(fch_issu1_inferred_i_64_n_0),
        .I1(fch_issu1_inferred_i_65_n_0),
        .O(fch_issu1_inferred_i_25_n_0),
        .S(fch_issu1_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'h00000000DD0FDDDD)) 
    fch_issu1_inferred_i_26
       (.I0(\fch/fadr_1_fl ),
        .I1(\nir_id[18]_i_2_n_0 ),
        .I2(\fch/nir_id [18]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fch_issu1_inferred_i_66_n_0),
        .O(fch_issu1_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h0FDD0FDD00000FDD)) 
    fch_issu1_inferred_i_27
       (.I0(\fch/fadr_1_fl ),
        .I1(\nir_id[12]_i_2_n_0 ),
        .I2(\fch/nir_id [12]),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_67_n_0),
        .I5(fch_issu1_inferred_i_68_n_0),
        .O(fch_issu1_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hF2F22222F2F2FF22)) 
    fch_issu1_inferred_i_28
       (.I0(fch_issu1_inferred_i_67_n_0),
        .I1(fch_issu1_inferred_i_69_n_0),
        .I2(\fch/nir_id [14]),
        .I3(\fch/fadr_1_fl ),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(\nir_id[14]_i_2_n_0 ),
        .O(fch_issu1_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h0000FF0FDD0DDD0D)) 
    fch_issu1_inferred_i_29
       (.I0(\fch/fadr_1_fl ),
        .I1(\nir_id[13]_i_2_n_0 ),
        .I2(fch_issu1_inferred_i_67_n_0),
        .I3(fch_issu1_inferred_i_70_n_0),
        .I4(\fch/nir_id [13]),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h0FDD0FDD00000FDD)) 
    fch_issu1_inferred_i_3
       (.I0(\fch/fadr_1_fl ),
        .I1(\nir_id[19]_i_2_n_0 ),
        .I2(\fch/nir_id [19]),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_14_n_0),
        .I5(fch_issu1_inferred_i_15_n_0),
        .O(fch_issu1_inferred_i_3_n_0));
  LUT6 #(
    .INIT(64'h0000000004000004)) 
    fch_issu1_inferred_i_30
       (.I0(fch_issu1_inferred_i_54_n_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fdat[24]),
        .I4(fdat[27]),
        .I5(fch_issu1_inferred_i_45_n_0),
        .O(fch_issu1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h0E0E0E0EFFFFFF00)) 
    fch_issu1_inferred_i_31
       (.I0(fch_issu1_inferred_i_71_n_0),
        .I1(fch_issu1_inferred_i_72_n_0),
        .I2(fch_issu1_inferred_i_73_n_0),
        .I3(fch_issu1_inferred_i_74_n_0),
        .I4(\fch/fadr_1_fl ),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(fch_issu1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFFF01)) 
    fch_issu1_inferred_i_32
       (.I0(fch_issu1_inferred_i_75_n_0),
        .I1(fdat[28]),
        .I2(fch_issu1_inferred_i_76_n_0),
        .I3(fch_issu1_inferred_i_77_n_0),
        .I4(fch_issu1_inferred_i_78_n_0),
        .I5(fch_issu1_inferred_i_79_n_0),
        .O(fch_issu1_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h0700F7FFF7FFF7FF)) 
    fch_issu1_inferred_i_33
       (.I0(fch_issu1_inferred_i_80_n_0),
        .I1(fdat[16]),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(fdat[0]),
        .I5(fch_issu1_inferred_i_41_n_0),
        .O(fch_issu1_inferred_i_33_n_0));
  LUT4 #(
    .INIT(16'hF66F)) 
    fch_issu1_inferred_i_34
       (.I0(fch_issu1_inferred_i_43_n_0),
        .I1(fch_issu1_inferred_i_29_n_0),
        .I2(fch_issu1_inferred_i_44_n_0),
        .I3(fch_issu1_inferred_i_28_n_0),
        .O(fch_issu1_inferred_i_34_n_0));
  LUT6 #(
    .INIT(64'h6006000000000000)) 
    fch_issu1_inferred_i_35
       (.I0(fch_issu1_inferred_i_31_n_0),
        .I1(fch_issu1_inferred_i_29_n_0),
        .I2(fch_issu1_inferred_i_28_n_0),
        .I3(fch_issu1_inferred_i_32_n_0),
        .I4(fch_issu1_inferred_i_7_n_0),
        .I5(fch_issu1_inferred_i_27_n_0),
        .O(fch_issu1_inferred_i_35_n_0));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    fch_issu1_inferred_i_36
       (.I0(fch_issu1_inferred_i_81_n_0),
        .I1(fdat[31]),
        .I2(fdat[25]),
        .I3(fch_issu1_inferred_i_82_n_0),
        .I4(fch_issu1_inferred_i_83_n_0),
        .I5(\fch/nir_id [24]),
        .O(fch_issu1_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF00F2)) 
    fch_issu1_inferred_i_37
       (.I0(\nir_id[21]_i_6_n_0 ),
        .I1(fch_issu1_inferred_i_84_n_0),
        .I2(fch_issu1_inferred_i_85_n_0),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_16_n_0),
        .I5(\fch/fadr_1_fl ),
        .O(fch_issu1_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'hBFBBBBBBAAAAAAAA)) 
    fch_issu1_inferred_i_38
       (.I0(fdat[31]),
        .I1(fch_issu1_inferred_i_86_n_0),
        .I2(fdat[20]),
        .I3(\ir0_id_fl[21]_i_5_n_0 ),
        .I4(fch_issu1_inferred_i_87_n_0),
        .I5(fch_issu1_inferred_i_88_n_0),
        .O(fch_issu1_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDFDFFF)) 
    fch_issu1_inferred_i_39
       (.I0(fch_issu1_inferred_i_89_n_0),
        .I1(fdat[31]),
        .I2(fdat[26]),
        .I3(fch_issu1_inferred_i_90_n_0),
        .I4(fdat[25]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'hB0B00000B0B0FF00)) 
    fch_issu1_inferred_i_4
       (.I0(fch_issu1_inferred_i_16_n_0),
        .I1(fch_issu1_inferred_i_17_n_0),
        .I2(fch_issu1_inferred_i_18_n_0),
        .I3(fch_issu1_inferred_i_19_n_0),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fch_issu1_inferred_i_20_n_0),
        .O(fch_issu1_inferred_i_4_n_0));
  LUT6 #(
    .INIT(64'h8080808090808080)) 
    fch_issu1_inferred_i_40
       (.I0(fdat[25]),
        .I1(fdat[26]),
        .I2(fdat[27]),
        .I3(fdat[24]),
        .I4(fdat[22]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_40_n_0));
  LUT6 #(
    .INIT(64'h0000001500000000)) 
    fch_issu1_inferred_i_41
       (.I0(fch_issu1_inferred_i_91_n_0),
        .I1(\nir_id[19]_i_7_n_0 ),
        .I2(fdat[11]),
        .I3(fch_issu1_inferred_i_92_n_0),
        .I4(\fch/fadr_1_fl ),
        .I5(fch_issu1_inferred_i_93_n_0),
        .O(fch_issu1_inferred_i_41_n_0));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFFFF)) 
    fch_issu1_inferred_i_42
       (.I0(fdat[11]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[6]),
        .O(fch_issu1_inferred_i_42_n_0));
  LUT6 #(
    .INIT(64'h0F440F0F00440000)) 
    fch_issu1_inferred_i_43
       (.I0(fdat[17]),
        .I1(fch_issu1_inferred_i_80_n_0),
        .I2(fdat[1]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fch_issu1_inferred_i_41_n_0),
        .O(fch_issu1_inferred_i_43_n_0));
  LUT6 #(
    .INIT(64'h0F440F0F00440000)) 
    fch_issu1_inferred_i_44
       (.I0(fdat[18]),
        .I1(fch_issu1_inferred_i_80_n_0),
        .I2(fdat[2]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fch_issu1_inferred_i_41_n_0),
        .O(fch_issu1_inferred_i_44_n_0));
  LUT3 #(
    .INIT(8'hBA)) 
    fch_issu1_inferred_i_45
       (.I0(\fch/fadr_1_fl ),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [1]),
        .O(fch_issu1_inferred_i_45_n_0));
  LUT6 #(
    .INIT(64'h3FFF7FFFFFFF7FFF)) 
    fch_issu1_inferred_i_46
       (.I0(fch_issu1_inferred_i_94_n_0),
        .I1(fdat[28]),
        .I2(fdat[29]),
        .I3(fdat[30]),
        .I4(fdat[27]),
        .I5(fch_issu1_inferred_i_95_n_0),
        .O(fch_issu1_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    fch_issu1_inferred_i_47
       (.I0(fdat[27]),
        .I1(fdat[26]),
        .I2(fdat[24]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_47_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_48
       (.I0(fdat[26]),
        .I1(fdat[27]),
        .O(fch_issu1_inferred_i_48_n_0));
  LUT4 #(
    .INIT(16'hEFFF)) 
    fch_issu1_inferred_i_49
       (.I0(fdat[25]),
        .I1(fdat[24]),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .O(fch_issu1_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h6FF6FFFFFFFF6FF6)) 
    fch_issu1_inferred_i_5
       (.I0(fch_issu1_inferred_i_21_n_0),
        .I1(fch_issu1_inferred_i_22_n_0),
        .I2(fch_issu1_inferred_i_23_n_0),
        .I3(fch_issu1_inferred_i_24_n_0),
        .I4(fch_issu1_inferred_i_25_n_0),
        .I5(fch_issu1_inferred_i_26_n_0),
        .O(fch_issu1_inferred_i_5_n_0));
  LUT6 #(
    .INIT(64'h00000000AE000000)) 
    fch_issu1_inferred_i_50
       (.I0(fch_issu1_inferred_i_96_n_0),
        .I1(fdat[20]),
        .I2(fch_issu1_inferred_i_97_n_0),
        .I3(fch_issu1_inferred_i_48_n_0),
        .I4(fdat[25]),
        .I5(fch_issu1_inferred_i_98_n_0),
        .O(fch_issu1_inferred_i_50_n_0));
  LUT6 #(
    .INIT(64'hC6FFFFFF86FFFFFF)) 
    fch_issu1_inferred_i_51
       (.I0(fdat[20]),
        .I1(fdat[21]),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .I4(fdat[24]),
        .I5(fdat[19]),
        .O(fch_issu1_inferred_i_51_n_0));
  LUT6 #(
    .INIT(64'h0000D7F5FFFFFFFF)) 
    fch_issu1_inferred_i_52
       (.I0(fdat[22]),
        .I1(fdat[21]),
        .I2(fdat[20]),
        .I3(fdat[19]),
        .I4(fch_issu1_inferred_i_99_n_0),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_52_n_0));
  LUT4 #(
    .INIT(16'h0004)) 
    fch_issu1_inferred_i_53
       (.I0(fdat[25]),
        .I1(fdat[23]),
        .I2(fdat[22]),
        .I3(fdat[24]),
        .O(fch_issu1_inferred_i_53_n_0));
  LUT4 #(
    .INIT(16'hBFFF)) 
    fch_issu1_inferred_i_54
       (.I0(fdat[31]),
        .I1(fdat[30]),
        .I2(fdat[29]),
        .I3(fdat[28]),
        .O(fch_issu1_inferred_i_54_n_0));
  LUT6 #(
    .INIT(64'h000A06020FFF2FAF)) 
    fch_issu1_inferred_i_55
       (.I0(fdat[24]),
        .I1(fdat[23]),
        .I2(fdat[26]),
        .I3(fdat[22]),
        .I4(fdat[25]),
        .I5(fdat[27]),
        .O(fch_issu1_inferred_i_55_n_0));
  LUT5 #(
    .INIT(32'hBFBFBFFF)) 
    fch_issu1_inferred_i_56
       (.I0(fch_issu1_inferred_i_100_n_0),
        .I1(fdat[13]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .I4(fch_issu1_inferred_i_101_n_0),
        .O(fch_issu1_inferred_i_56_n_0));
  LUT6 #(
    .INIT(64'h5D55DD005D55DDDD)) 
    fch_issu1_inferred_i_57
       (.I0(fch_issu1_inferred_i_102_n_0),
        .I1(fch_issu1_inferred_i_103_n_0),
        .I2(fch_issu1_inferred_i_104_n_0),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fch_issu1_inferred_i_105_n_0),
        .O(fch_issu1_inferred_i_57_n_0));
  LUT6 #(
    .INIT(64'hF2F2F2F2F2F2F200)) 
    fch_issu1_inferred_i_58
       (.I0(fdat[24]),
        .I1(fch_issu1_inferred_i_45_n_0),
        .I2(fch_issu1_inferred_i_106_n_0),
        .I3(fch_issu1_inferred_i_107_n_0),
        .I4(fdat[31]),
        .I5(fch_issu1_inferred_i_108_n_0),
        .O(fch_issu1_inferred_i_58_n_0));
  LUT5 #(
    .INIT(32'hA3FFAFFF)) 
    fch_issu1_inferred_i_59
       (.I0(fch_issu1_inferred_i_109_n_0),
        .I1(fdat[3]),
        .I2(fdat[11]),
        .I3(fdat[12]),
        .I4(fch_issu1_inferred_i_101_n_0),
        .O(fch_issu1_inferred_i_59_n_0));
  LUT6 #(
    .INIT(64'h0990000000000990)) 
    fch_issu1_inferred_i_6
       (.I0(fch_issu1_inferred_i_27_n_0),
        .I1(fch_issu1_inferred_i_22_n_0),
        .I2(fch_issu1_inferred_i_25_n_0),
        .I3(fch_issu1_inferred_i_28_n_0),
        .I4(fch_issu1_inferred_i_23_n_0),
        .I5(fch_issu1_inferred_i_29_n_0),
        .O(fch_issu1_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'hFFF8F0F0F8F8F0F0)) 
    fch_issu1_inferred_i_60
       (.I0(fch_issu1_inferred_i_110_n_0),
        .I1(fch_issu1_inferred_i_111_n_0),
        .I2(fch_issu1_inferred_i_112_n_0),
        .I3(fch_issu1_inferred_i_17_n_0),
        .I4(fch_issu1_inferred_i_13_n_0),
        .I5(fdat[24]),
        .O(fch_issu1_inferred_i_60_n_0));
  LUT6 #(
    .INIT(64'h00000000FFBB000B)) 
    fch_issu1_inferred_i_61
       (.I0(fch_issu1_inferred_i_113_n_0),
        .I1(fdat[14]),
        .I2(\fch/fadr_1_fl ),
        .I3(fdat[15]),
        .I4(fch_issu1_inferred_i_114_n_0),
        .I5(fch_issu1_inferred_i_115_n_0),
        .O(fch_issu1_inferred_i_61_n_0));
  LUT5 #(
    .INIT(32'hD0FFD0D0)) 
    fch_issu1_inferred_i_62
       (.I0(fdat[30]),
        .I1(fch_issu1_inferred_i_116_n_0),
        .I2(fch_issu1_inferred_i_117_n_0),
        .I3(fdat[25]),
        .I4(fch_issu1_inferred_i_17_n_0),
        .O(fch_issu1_inferred_i_62_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00A2)) 
    fch_issu1_inferred_i_63
       (.I0(fdat[25]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fch_issu1_inferred_i_106_n_0),
        .I5(fch_issu1_inferred_i_118_n_0),
        .O(fch_issu1_inferred_i_63_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF2203)) 
    fch_issu1_inferred_i_64
       (.I0(fch_issu1_inferred_i_119_n_0),
        .I1(fch_issu1_inferred_i_56_n_0),
        .I2(fdat[5]),
        .I3(\nir_id[21]_i_9_n_0 ),
        .I4(fch_issu1_inferred_i_92_n_0),
        .I5(fch_issu1_inferred_i_120_n_0),
        .O(fch_issu1_inferred_i_64_n_0));
  LUT6 #(
    .INIT(64'h7500FFFF75007500)) 
    fch_issu1_inferred_i_65
       (.I0(fdat[30]),
        .I1(fch_issu1_inferred_i_121_n_0),
        .I2(fch_issu1_inferred_i_122_n_0),
        .I3(fch_issu1_inferred_i_117_n_0),
        .I4(fdat[26]),
        .I5(fch_issu1_inferred_i_17_n_0),
        .O(fch_issu1_inferred_i_65_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF00A2)) 
    fch_issu1_inferred_i_66
       (.I0(fdat[26]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fch_issu1_inferred_i_106_n_0),
        .I5(fch_issu1_inferred_i_123_n_0),
        .O(fch_issu1_inferred_i_66_n_0));
  LUT6 #(
    .INIT(64'h4155455540554055)) 
    fch_issu1_inferred_i_67
       (.I0(fch_issu1_inferred_i_45_n_0),
        .I1(fdat[28]),
        .I2(fdat[29]),
        .I3(fdat[31]),
        .I4(fdat[27]),
        .I5(fdat[30]),
        .O(fch_issu1_inferred_i_67_n_0));
  LUT6 #(
    .INIT(64'h20AA20AA20AAAAAA)) 
    fch_issu1_inferred_i_68
       (.I0(fch_issu1_inferred_i_124_n_0),
        .I1(fch_issu1_inferred_i_125_n_0),
        .I2(fch_issu1_inferred_i_126_n_0),
        .I3(fdat[30]),
        .I4(fch_issu1_inferred_i_127_n_0),
        .I5(fch_issu1_inferred_i_128_n_0),
        .O(fch_issu1_inferred_i_68_n_0));
  LUT6 #(
    .INIT(64'h20AA20AA20AAAAAA)) 
    fch_issu1_inferred_i_69
       (.I0(fch_issu1_inferred_i_124_n_0),
        .I1(fch_issu1_inferred_i_129_n_0),
        .I2(fch_issu1_inferred_i_126_n_0),
        .I3(fdat[30]),
        .I4(fch_issu1_inferred_i_127_n_0),
        .I5(fch_issu1_inferred_i_130_n_0),
        .O(fch_issu1_inferred_i_69_n_0));
  LUT6 #(
    .INIT(64'h0D0F0D0D0D000D0D)) 
    fch_issu1_inferred_i_7
       (.I0(\fch/fadr_1_fl ),
        .I1(\fch/lir_id_0 [15]),
        .I2(fch_issu1_inferred_i_30_n_0),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(\fch/nir_id [15]),
        .O(fch_issu1_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'h0000080008080808)) 
    fch_issu1_inferred_i_70
       (.I0(fdat[30]),
        .I1(fdat[29]),
        .I2(fdat[31]),
        .I3(fch_issu1_inferred_i_126_n_0),
        .I4(fch_issu1_inferred_i_131_n_0),
        .I5(fch_issu1_inferred_i_132_n_0),
        .O(fch_issu1_inferred_i_70_n_0));
  LUT6 #(
    .INIT(64'hFFFFF7FFFFFFFFFF)) 
    fch_issu1_inferred_i_71
       (.I0(fdat[21]),
        .I1(fdat[25]),
        .I2(fdat[23]),
        .I3(fch_issu1_inferred_i_133_n_0),
        .I4(fdat[31]),
        .I5(fdat[22]),
        .O(fch_issu1_inferred_i_71_n_0));
  LUT3 #(
    .INIT(8'h7F)) 
    fch_issu1_inferred_i_72
       (.I0(fdat[28]),
        .I1(fdat[26]),
        .I2(fdat[24]),
        .O(fch_issu1_inferred_i_72_n_0));
  LUT6 #(
    .INIT(64'h2000233330000330)) 
    fch_issu1_inferred_i_73
       (.I0(fch_issu1_inferred_i_134_n_0),
        .I1(fch_issu1_inferred_i_135_n_0),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .I4(fdat[31]),
        .I5(fdat[28]),
        .O(fch_issu1_inferred_i_73_n_0));
  LUT6 #(
    .INIT(64'hA8AAAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_74
       (.I0(fch_issu1_inferred_i_136_n_0),
        .I1(fch_issu1_inferred_i_137_n_0),
        .I2(fdat[15]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[5]),
        .O(fch_issu1_inferred_i_74_n_0));
  LUT6 #(
    .INIT(64'h0000A80000002800)) 
    fch_issu1_inferred_i_75
       (.I0(\ir0_id_fl[21]_i_7_n_0 ),
        .I1(fdat[19]),
        .I2(fdat[17]),
        .I3(fch_issu1_inferred_i_138_n_0),
        .I4(fdat[27]),
        .I5(fdat[16]),
        .O(fch_issu1_inferred_i_75_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_76
       (.I0(fdat[30]),
        .I1(fdat[29]),
        .O(fch_issu1_inferred_i_76_n_0));
  LUT6 #(
    .INIT(64'hFFFF0FFF00FF07FF)) 
    fch_issu1_inferred_i_77
       (.I0(fdat[26]),
        .I1(fch_issu1_inferred_i_139_n_0),
        .I2(fdat[27]),
        .I3(fch_issu1_inferred_i_13_n_0),
        .I4(fch_issu1_inferred_i_108_n_0),
        .I5(fdat[31]),
        .O(fch_issu1_inferred_i_77_n_0));
  LUT6 #(
    .INIT(64'h0000000022207775)) 
    fch_issu1_inferred_i_78
       (.I0(fdat[28]),
        .I1(fch_issu1_inferred_i_140_n_0),
        .I2(fch_issu1_inferred_i_141_n_0),
        .I3(fch_issu1_inferred_i_142_n_0),
        .I4(fdat[31]),
        .I5(fch_issu1_inferred_i_143_n_0),
        .O(fch_issu1_inferred_i_78_n_0));
  LUT6 #(
    .INIT(64'h00000000FBFFFBAA)) 
    fch_issu1_inferred_i_79
       (.I0(fch_issu1_inferred_i_144_n_0),
        .I1(fch_issu1_inferred_i_145_n_0),
        .I2(fch_issu1_inferred_i_146_n_0),
        .I3(fdat[12]),
        .I4(fdat[15]),
        .I5(fch_issu1_inferred_i_147_n_0),
        .O(fch_issu1_inferred_i_79_n_0));
  LUT5 #(
    .INIT(32'hF99FFFFF)) 
    fch_issu1_inferred_i_8
       (.I0(fch_issu1_inferred_i_24_n_0),
        .I1(fch_issu1_inferred_i_31_n_0),
        .I2(fch_issu1_inferred_i_26_n_0),
        .I3(fch_issu1_inferred_i_32_n_0),
        .I4(fch_issu1_inferred_i_21_n_0),
        .O(fch_issu1_inferred_i_8_n_0));
  LUT6 #(
    .INIT(64'h000076AA00000000)) 
    fch_issu1_inferred_i_80
       (.I0(fdat[27]),
        .I1(fdat[25]),
        .I2(fch_issu1_inferred_i_90_n_0),
        .I3(fdat[26]),
        .I4(fdat[31]),
        .I5(fch_issu1_inferred_i_89_n_0),
        .O(fch_issu1_inferred_i_80_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    fch_issu1_inferred_i_81
       (.I0(fdat[26]),
        .I1(fdat[27]),
        .O(fch_issu1_inferred_i_81_n_0));
  LUT6 #(
    .INIT(64'h5554555555555555)) 
    fch_issu1_inferred_i_82
       (.I0(fch_issu1_inferred_i_89_n_0),
        .I1(fch_issu1_inferred_i_148_n_0),
        .I2(fdat[24]),
        .I3(fdat[18]),
        .I4(fch_issu1_inferred_i_149_n_0),
        .I5(fch_issu1_inferred_i_138_n_0),
        .O(fch_issu1_inferred_i_82_n_0));
  LUT6 #(
    .INIT(64'h0000110100004000)) 
    fch_issu1_inferred_i_83
       (.I0(fch_issu1_inferred_i_54_n_0),
        .I1(fdat[27]),
        .I2(fdat[26]),
        .I3(fch_issu1_inferred_i_150_n_0),
        .I4(fdat[24]),
        .I5(fdat[25]),
        .O(fch_issu1_inferred_i_83_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFF00)) 
    fch_issu1_inferred_i_84
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[10]),
        .I4(fdat[11]),
        .I5(fdat[9]),
        .O(fch_issu1_inferred_i_84_n_0));
  LUT6 #(
    .INIT(64'hBAAEAAAAAAAAAAAA)) 
    fch_issu1_inferred_i_85
       (.I0(fch_issu1_inferred_i_151_n_0),
        .I1(fdat[0]),
        .I2(fdat[3]),
        .I3(fdat[1]),
        .I4(fch_issu1_inferred_i_152_n_0),
        .I5(fch_issu1_inferred_i_153_n_0),
        .O(fch_issu1_inferred_i_85_n_0));
  LUT6 #(
    .INIT(64'hAAAAABEAAAAAAAAA)) 
    fch_issu1_inferred_i_86
       (.I0(fch_issu1_inferred_i_154_n_0),
        .I1(fdat[26]),
        .I2(fdat[25]),
        .I3(fch_issu1_inferred_i_138_n_0),
        .I4(fch_issu1_inferred_i_155_n_0),
        .I5(fch_issu1_inferred_i_156_n_0),
        .O(fch_issu1_inferred_i_86_n_0));
  LUT3 #(
    .INIT(8'h41)) 
    fch_issu1_inferred_i_87
       (.I0(fdat[17]),
        .I1(fdat[16]),
        .I2(fdat[19]),
        .O(fch_issu1_inferred_i_87_n_0));
  LUT4 #(
    .INIT(16'hF001)) 
    fch_issu1_inferred_i_88
       (.I0(fdat[28]),
        .I1(fdat[27]),
        .I2(fdat[30]),
        .I3(fdat[29]),
        .O(fch_issu1_inferred_i_88_n_0));
  LUT3 #(
    .INIT(8'h80)) 
    fch_issu1_inferred_i_89
       (.I0(fdat[28]),
        .I1(fdat[29]),
        .I2(fdat[30]),
        .O(fch_issu1_inferred_i_89_n_0));
  LUT5 #(
    .INIT(32'hFFFF6FF6)) 
    fch_issu1_inferred_i_9
       (.I0(fch_issu1_inferred_i_7_n_0),
        .I1(fch_issu1_inferred_i_11_n_0),
        .I2(fch_issu1_inferred_i_27_n_0),
        .I3(fch_issu1_inferred_i_33_n_0),
        .I4(fch_issu1_inferred_i_34_n_0),
        .O(fch_issu1_inferred_i_9_n_0));
  LUT3 #(
    .INIT(8'h8F)) 
    fch_issu1_inferred_i_90
       (.I0(fdat[22]),
        .I1(fdat[23]),
        .I2(fdat[24]),
        .O(fch_issu1_inferred_i_90_n_0));
  LUT6 #(
    .INIT(64'h0000150055555555)) 
    fch_issu1_inferred_i_91
       (.I0(fdat[11]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(fch_issu1_inferred_i_91_n_0));
  LUT2 #(
    .INIT(4'hB)) 
    fch_issu1_inferred_i_92
       (.I0(fdat[15]),
        .I1(fdat[14]),
        .O(fch_issu1_inferred_i_92_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_issu1_inferred_i_93
       (.I0(fdat[13]),
        .I1(fdat[12]),
        .O(fch_issu1_inferred_i_93_n_0));
  LUT5 #(
    .INIT(32'h319977BF)) 
    fch_issu1_inferred_i_94
       (.I0(fdat[26]),
        .I1(fdat[25]),
        .I2(fdat[23]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .O(fch_issu1_inferred_i_94_n_0));
  LUT5 #(
    .INIT(32'hDDDFFFDF)) 
    fch_issu1_inferred_i_95
       (.I0(fdat[25]),
        .I1(fdat[26]),
        .I2(fdat[23]),
        .I3(fdat[24]),
        .I4(fdat[22]),
        .O(fch_issu1_inferred_i_95_n_0));
  LUT6 #(
    .INIT(64'h503FFFFFFFFFFFFF)) 
    fch_issu1_inferred_i_96
       (.I0(fdat[19]),
        .I1(fdat[20]),
        .I2(fdat[21]),
        .I3(fdat[22]),
        .I4(fdat[24]),
        .I5(fdat[23]),
        .O(fch_issu1_inferred_i_96_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    fch_issu1_inferred_i_97
       (.I0(fdat[21]),
        .I1(fdat[22]),
        .O(fch_issu1_inferred_i_97_n_0));
  LUT6 #(
    .INIT(64'h0400400000004404)) 
    fch_issu1_inferred_i_98
       (.I0(fdat[23]),
        .I1(fdat[24]),
        .I2(fdat[19]),
        .I3(fdat[22]),
        .I4(fdat[21]),
        .I5(fdat[20]),
        .O(fch_issu1_inferred_i_98_n_0));
  LUT5 #(
    .INIT(32'hFF0EFFFF)) 
    fch_issu1_inferred_i_99
       (.I0(fdat[21]),
        .I1(fdat[20]),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .I4(fdat[24]),
        .O(fch_issu1_inferred_i_99_n_0));
  LUT6 #(
    .INIT(64'h8B888B8B8B8B8B8B)) 
    fch_leir_hir_i_1
       (.I0(fch_leir_hir_i_2_n_0),
        .I1(\fadr[15]_INST_0_i_5_n_0 ),
        .I2(\rgf/pcnt/pc [1]),
        .I3(\fch/stat [2]),
        .I4(\fch/stat [0]),
        .I5(\fch/stat [1]),
        .O(\fch/fctl/fch_leir_hir_t ));
  LUT5 #(
    .INIT(32'h0000091C)) 
    fch_leir_hir_i_2
       (.I0(\fch/stat [2]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fch_issu1_ir ),
        .I4(fch_leir_nir_i_2_n_0),
        .O(fch_leir_hir_i_2_n_0));
  LUT5 #(
    .INIT(32'h0000AA2A)) 
    fch_leir_lir_i_1
       (.I0(\rgf/pcnt/pc [1]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [2]),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\fch/fctl/fch_leir_lir_t ));
  LUT6 #(
    .INIT(64'h0002020000020002)) 
    fch_leir_nir_i_1
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\fch/stat [0]),
        .I2(fch_leir_nir_i_2_n_0),
        .I3(\fch/stat [1]),
        .I4(\fch/stat [2]),
        .I5(\fch/fch_issu1_ir ),
        .O(\fch/fctl/fch_leir_nir_t ));
  LUT2 #(
    .INIT(4'hE)) 
    fch_leir_nir_i_2
       (.I0(fch_term),
        .I1(\nir_id[24]_i_6_n_0 ),
        .O(fch_leir_nir_i_2_n_0));
  LUT2 #(
    .INIT(4'h8)) 
    fch_term_fl_i_1
       (.I0(ctl_fetch0),
        .I1(ctl_fetch1),
        .O(fch_term));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [0]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[0]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[0]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[0]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[0]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[0]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[0]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[0]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[0]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[0]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[0]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[0]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[0]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[0]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[0]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[0]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[0]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[0]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[0]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[0]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[0]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[0]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[0]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[0]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[0]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[0]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [0]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c0bus_0 [0]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[0]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[0]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[0]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[0]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[0]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[0]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[0]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/rgf_c0bus_0 [0]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[0]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [10]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[10]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[10]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[10]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[10]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[10]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[10]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[10]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[10]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[10]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[10]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[10]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[10]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[10]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[10]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[10]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[10]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[10]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[10]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[10]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[10]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[10]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[10]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[10]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[10]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[10]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [10]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c0bus_0 [10]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[10]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[10]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[10]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[10]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[10]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[10]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[10]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/rgf_c0bus_0 [10]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[10]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [11]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[11]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[11]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[11]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[11]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[11]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[11]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[11]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[11]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[11]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[11]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[11]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[11]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[11]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[11]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[11]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[11]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[11]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[11]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[11]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[11]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[11]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[11]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[11]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[11]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[11]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [11]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c0bus_0 [11]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[11]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[11]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[11]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[11]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[11]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[11]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[11]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/rgf_c0bus_0 [11]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[11]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [12]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[12]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[12]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[12]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[12]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[12]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[12]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[12]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[12]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[12]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[12]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[12]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[12]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[12]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[12]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[12]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[12]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[12]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[12]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[12]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[12]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[12]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[12]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[12]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[12]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[12]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [12]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c0bus_0 [12]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[12]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[12]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[12]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[12]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[12]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[12]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[12]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/rgf_c0bus_0 [12]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[12]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [13]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[13]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[13]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[13]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[13]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[13]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[13]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[13]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[13]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[13]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[13]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[13]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[13]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[13]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[13]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[13]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[13]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[13]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[13]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[13]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[13]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[13]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[13]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[13]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[13]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[13]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [13]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c0bus_0 [13]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[13]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[13]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[13]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[13]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[13]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[13]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[13]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/rgf_c0bus_0 [13]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[13]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [14]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[14]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[14]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[14]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[14]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[14]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[14]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[14]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[14]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[14]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[14]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[14]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[14]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[14]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[14]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[14]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[14]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[14]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[14]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[14]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[14]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[14]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[14]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[14]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[14]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[14]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [14]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c0bus_0 [14]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[14]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[14]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[14]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[14]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[14]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[14]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[14]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/rgf_c0bus_0 [14]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[14]_i_1__9_n_0 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1 
       (.I0(\rgf/bank02/grn07/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [7]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__0 
       (.I0(\rgf/bank02/grn06/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [6]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__1 
       (.I0(\rgf/bank02/grn05/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [5]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__1_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__10 
       (.I0(\rgf/bank13/grn21/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__10_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__11 
       (.I0(\rgf/bank02/grn27/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [7]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__11_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__12 
       (.I0(\rgf/bank02/grn26/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [6]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__12_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__13 
       (.I0(\rgf/bank02/grn25/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [5]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__13_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__14 
       (.I0(\rgf/bank02/grn24/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [4]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__14_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__15 
       (.I0(\rgf/bank02/grn22/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [2]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__15_n_0 ));
  LUT5 #(
    .INIT(32'hAEAEAEAA)) 
    \grn[15]_i_1__16 
       (.I0(\rgf/bank02/grn21/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__16_n_0 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__17 
       (.I0(\rgf/bank13/grn07/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [7]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__17_n_0 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__18 
       (.I0(\rgf/bank13/grn02/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [2]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__18_n_0 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__19 
       (.I0(\rgf/bank13/grn01/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__19_n_0 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__2 
       (.I0(\rgf/bank02/grn04/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [4]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__2_n_0 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__20 
       (.I0(\rgf/bank13/grn06/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [6]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__20_n_0 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__21 
       (.I0(\rgf/bank13/grn04/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [4]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__21_n_0 ));
  LUT5 #(
    .INIT(32'hEAAAEAEA)) 
    \grn[15]_i_1__22 
       (.I0(\rgf/bank13/grn05/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [5]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hF1F0F0F0F1F0F1F0)) 
    \grn[15]_i_1__23 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hF0F1F0F1F0F1F0F0)) 
    \grn[15]_i_1__24 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn23/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hF1F0F1F0F1F0F0F0)) 
    \grn[15]_i_1__25 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank13/grn23/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hF0F1F0F0F0F1F0F1)) 
    \grn[15]_i_1__26 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_3_n_0 ),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hF1F0F0F0F1F0F1F0)) 
    \grn[15]_i_1__27 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_4__2_n_0 ),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hF0F1F0F1F0F1F0F0)) 
    \grn[15]_i_1__28 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_4__2_n_0 ),
        .I2(\rgf/bank02/grn20/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hF1F0F1F0F1F0F0F0)) 
    \grn[15]_i_1__29 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_4__2_n_0 ),
        .I2(\rgf/bank13/grn20/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__29_n_0 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__3 
       (.I0(\rgf/bank02/grn02/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [2]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hF0F1F0F0F0F1F0F1)) 
    \grn[15]_i_1__30 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\grn[15]_i_4__2_n_0 ),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__30_n_0 ));
  LUT5 #(
    .INIT(32'hAEAAAEAE)) 
    \grn[15]_i_1__4 
       (.I0(\rgf/bank02/grn01/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__5 
       (.I0(\rgf/bank13/grn27/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [7]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__5_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__6 
       (.I0(\rgf/bank13/grn26/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [6]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__7 
       (.I0(\rgf/bank13/grn25/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [5]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__7_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__8 
       (.I0(\rgf/bank13/grn24/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [4]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__8_n_0 ));
  LUT5 #(
    .INIT(32'hEAEAEAAA)) 
    \grn[15]_i_1__9 
       (.I0(\rgf/bank13/grn22/grn1__0 ),
        .I1(\rgf/c0bus_sel_0 [2]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [15]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__0 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[15]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[15]_i_2__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__10 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[15]_i_2__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__11 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[15]_i_2__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__12 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[15]_i_2__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__13 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[15]_i_2__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__14 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[15]_i_2__14_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__15 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[15]_i_2__15_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__16 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[15]_i_2__16_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__17 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[15]_i_2__17_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__18 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[15]_i_2__18_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__19 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[15]_i_2__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__2 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[15]_i_2__2_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__20 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[15]_i_2__20_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__21 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[15]_i_2__21_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__22 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[15]_i_2__22_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__23 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[15]_i_2__23_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__24 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[15]_i_2__24_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__25 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[15]_i_2__25_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__26 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[15]_i_2__26_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__27 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[15]_i_2__27_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__28 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[15]_i_2__28_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__29 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[15]_i_2__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__3 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[15]_i_2__3_n_0 ));
  LUT5 #(
    .INIT(32'hB8B8FF00)) 
    \grn[15]_i_2__30 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [15]),
        .I3(\rgf/c0bus_bk2 ),
        .I4(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[15]_i_2__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__4 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[15]_i_2__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__5 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[15]_i_2__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__6 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[15]_i_2__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__7 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[15]_i_2__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__8 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[15]_i_2__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[15]_i_2__9 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/rgf_c0bus_0 [15]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[15]_i_2__9_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .O(\grn[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__0 
       (.I0(\rgf/bank_sel [0]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn01/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__1 
       (.I0(\rgf/bank_sel [0]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn02/grn1__0 ));
  LUT6 #(
    .INIT(64'h00000000000000E0)) 
    \grn[15]_i_3__10 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn23/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__11 
       (.I0(\grn[15]_i_4__6_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn22/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__12 
       (.I0(\grn[15]_i_4__6_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn21/grn1__0 ));
  LUT6 #(
    .INIT(64'h00000000000000E0)) 
    \grn[15]_i_3__13 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\tr[31]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn20/grn1__0 ));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    \grn[15]_i_3__14 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\tr[31]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn20/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__15 
       (.I0(\rgf/bank_sel [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn21/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__16 
       (.I0(\rgf/bank_sel [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn22/grn1__0 ));
  LUT6 #(
    .INIT(64'h000000000000000E)) 
    \grn[15]_i_3__17 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn23/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__18 
       (.I0(\rgf/bank_sel [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn24/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__19 
       (.I0(\rgf/bank_sel [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn25/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__2 
       (.I0(\rgf/bank_sel [0]),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn04/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__20 
       (.I0(\rgf/bank_sel [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn26/grn1__0 ));
  LUT6 #(
    .INIT(64'h0000000E00000000)) 
    \grn[15]_i_3__21 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\grn[15]_i_7__0_n_0 ),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn27/grn1__0 ));
  LUT6 #(
    .INIT(64'h000000D000000000)) 
    \grn[15]_i_3__22 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\grn[15]_i_7__0_n_0 ),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn07/grn1__0 ));
  LUT6 #(
    .INIT(64'h00000000000000D0)) 
    \grn[15]_i_3__23 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn03/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__24 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn02/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__25 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn01/grn1__0 ));
  LUT6 #(
    .INIT(64'h00000000000000D0)) 
    \grn[15]_i_3__26 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\tr[31]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn00/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__27 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn06/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__28 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn04/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__29 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn05/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__3 
       (.I0(\rgf/bank_sel [0]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn05/grn1__0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_3__30 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_6__0_n_0 ),
        .O(\grn[15]_i_3__30_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__4 
       (.I0(\rgf/bank_sel [0]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn06/grn1__0 ));
  LUT6 #(
    .INIT(64'h0000000D00000000)) 
    \grn[15]_i_3__5 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\grn[15]_i_7__0_n_0 ),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank02/grn07/grn1__0 ));
  LUT6 #(
    .INIT(64'h000000E000000000)) 
    \grn[15]_i_3__6 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\grn[15]_i_7__0_n_0 ),
        .I5(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/bank13/grn27/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__7 
       (.I0(\grn[15]_i_4__6_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn26/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \grn[15]_i_3__8 
       (.I0(\grn[15]_i_4__6_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [1]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn25/grn1__0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \grn[15]_i_3__9 
       (.I0(\grn[15]_i_4__6_n_0 ),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank13/grn24/grn1__0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \grn[15]_i_4 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\grn[15]_i_6__0_n_0 ),
        .I2(\grn[15]_i_3_n_0 ),
        .O(\rgf/c0bus_sel_0 [7]));
  LUT3 #(
    .INIT(8'h04)) 
    \grn[15]_i_4__0 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .O(\rgf/c0bus_sel_0 [2]));
  LUT3 #(
    .INIT(8'h04)) 
    \grn[15]_i_4__1 
       (.I0(\grn[15]_i_3__30_n_0 ),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .O(\rgf/c0bus_sel_0 [1]));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_4__2 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [0]),
        .O(\grn[15]_i_4__2_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4__3 
       (.I0(\grn[15]_i_6__0_n_0 ),
        .I1(\rgf/rctl/p_0_in [1]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\rgf/rctl/p_0_in [2]),
        .O(\rgf/c0bus_sel_0 [5]));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \grn[15]_i_4__4 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\iv[15]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn03/grn1__0 ));
  LUT6 #(
    .INIT(64'hB8BBB888B888B888)) 
    \grn[15]_i_4__5 
       (.I0(\rgf/rgf_c0bus_0 [31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(c0bus[15]),
        .I3(fch_wrbufn0),
        .I4(fch_term),
        .I5(\grn[15]_i_5_n_0 ),
        .O(\rgf/c0bus_bk2 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \grn[15]_i_4__6 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_4__6_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \grn[15]_i_4__7 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [1]),
        .O(\grn[15]_i_4__7_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \grn[15]_i_4__8 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\grn[15]_i_6__0_n_0 ),
        .I2(\rgf/rctl/p_0_in [2]),
        .I3(\rgf/rctl/p_0_in [1]),
        .O(\rgf/c0bus_sel_0 [4]));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_4__9 
       (.I0(\rgf/rctl/p_0_in [0]),
        .I1(\grn[15]_i_6__0_n_0 ),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\rgf/rctl/p_0_in [2]),
        .O(\rgf/c0bus_sel_0 [6]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBB8)) 
    \grn[15]_i_5 
       (.I0(\rgf/rctl/rgf_c0bus_wb [15]),
        .I1(\rgf/rctl/rgf_selc0_stat ),
        .I2(\grn[15]_i_6_n_0 ),
        .I3(\grn[15]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .O(\grn[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000000D)) 
    \grn[15]_i_5__0 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\tr[31]_i_4_n_0 ),
        .I4(\rgf/rctl/rgf_selc1_rn [2]),
        .I5(\grn[15]_i_7__0_n_0 ),
        .O(\rgf/bank02/grn00/grn1__0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \grn[15]_i_6 
       (.I0(cbus_i[15]),
        .I1(ccmd[4]),
        .O(\grn[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h1B1F5F1FFFFFFFFF)) 
    \grn[15]_i_6__0 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(ctl_selc0[0]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_wb [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\grn[15]_i_6__0_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \grn[15]_i_7 
       (.I0(bdatr[15]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\grn[15]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_7__0 
       (.I0(\rgf/rctl/rgf_selc1 [1]),
        .I1(\rgf/rctl/rgf_selc1 [0]),
        .O(\grn[15]_i_7__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [1]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[1]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[1]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[1]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[1]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[1]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[1]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[1]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[1]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[1]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[1]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[1]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[1]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[1]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[1]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[1]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[1]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[1]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[1]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[1]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[1]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[1]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[1]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[1]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[1]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[1]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [1]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c0bus_0 [1]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[1]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[1]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[1]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[1]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[1]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[1]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[1]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/rgf_c0bus_0 [1]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[1]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [2]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[2]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[2]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[2]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[2]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[2]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[2]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[2]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__15 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[2]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__16 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[2]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__17 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[2]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__18 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[2]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__19 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[2]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[2]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__20 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[2]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__21 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[2]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__22 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[2]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__23 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[2]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__24 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[2]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__25 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[2]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__26 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[2]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__27 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[2]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__28 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[2]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__29 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[2]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[2]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[2]_i_1__30 
       (.I0(\rgf/rgf_c0bus_0 [18]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[2]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[2]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[2]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[2]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[2]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[2]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[2]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/rgf_c0bus_0 [2]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[2]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [3]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[3]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[3]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[3]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[3]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[3]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[3]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[3]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[3]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[3]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[3]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[3]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[3]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[3]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[3]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[3]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[3]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[3]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[3]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[3]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[3]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[3]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[3]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[3]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[3]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[3]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [3]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c0bus_0 [3]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[3]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[3]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[3]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[3]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[3]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[3]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[3]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/rgf_c0bus_0 [3]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[3]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [4]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[4]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[4]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[4]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[4]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[4]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[4]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[4]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__15 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[4]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__16 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[4]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__17 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[4]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__18 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[4]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__19 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[4]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[4]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__20 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[4]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__21 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[4]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__22 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[4]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__23 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[4]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__24 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[4]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__25 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[4]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__26 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[4]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__27 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[4]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__28 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[4]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__29 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[4]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[4]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[4]_i_1__30 
       (.I0(\rgf/rgf_c0bus_0 [20]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[4]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[4]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[4]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[4]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[4]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[4]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[4]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/rgf_c0bus_0 [4]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[4]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [5]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[5]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[5]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[5]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[5]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[5]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[5]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[5]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__15 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[5]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__16 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[5]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__17 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[5]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__18 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[5]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__19 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[5]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[5]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__20 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[5]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__21 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[5]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__22 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[5]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__23 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[5]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__24 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[5]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__25 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[5]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__26 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[5]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__27 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[5]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__28 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[5]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__29 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[5]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[5]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \grn[5]_i_1__30 
       (.I0(\rgf/rgf_c0bus_0 [21]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[5]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[5]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[5]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[5]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[5]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[5]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[5]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/rgf_c0bus_0 [5]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[5]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [6]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[6]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[6]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[6]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[6]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[6]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[6]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[6]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[6]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[6]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[6]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[6]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[6]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[6]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[6]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[6]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[6]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[6]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[6]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[6]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[6]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[6]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[6]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[6]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[6]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[6]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [6]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c0bus_0 [6]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[6]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[6]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[6]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[6]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[6]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[6]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[6]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[6]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [7]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[7]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[7]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[7]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[7]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[7]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[7]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[7]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[7]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[7]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[7]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[7]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[7]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[7]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[7]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[7]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[7]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[7]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[7]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[7]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[7]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[7]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[7]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[7]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[7]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[7]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [7]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c0bus_0 [7]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[7]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[7]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[7]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[7]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[7]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[7]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[7]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/rgf_c0bus_0 [7]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[7]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [8]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[8]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[8]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[8]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[8]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[8]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[8]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[8]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[8]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[8]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[8]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[8]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[8]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[8]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[8]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[8]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[8]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[8]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[8]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[8]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[8]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[8]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[8]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[8]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[8]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[8]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [8]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c0bus_0 [8]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[8]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[8]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[8]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[8]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[8]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[8]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[8]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/rgf_c0bus_0 [8]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[8]_i_1__9_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn00/grn1__0 ),
        .O(\rgf/p_2_in [9]));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__0 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn01/grn1__0 ),
        .O(\grn[9]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn02/grn1__0 ),
        .O(\grn[9]_i_1__1_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__10 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn01/grn1__0 ),
        .O(\grn[9]_i_1__10_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__11 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn00/grn1__0 ),
        .O(\grn[9]_i_1__11_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__12 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn02/grn1__0 ),
        .O(\grn[9]_i_1__12_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__13 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn04/grn1__0 ),
        .O(\grn[9]_i_1__13_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__14 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn06/grn1__0 ),
        .O(\grn[9]_i_1__14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__15 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn20/grn1__0 ),
        .O(\grn[9]_i_1__15_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__16 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn21/grn1__0 ),
        .O(\grn[9]_i_1__16_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__17 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn22/grn1__0 ),
        .O(\grn[9]_i_1__17_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__18 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn23/grn1__0 ),
        .O(\grn[9]_i_1__18_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__19 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn24/grn1__0 ),
        .O(\grn[9]_i_1__19_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__2 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn03/grn1__0 ),
        .O(\grn[9]_i_1__2_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__20 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn25/grn1__0 ),
        .O(\grn[9]_i_1__20_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__21 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn26/grn1__0 ),
        .O(\grn[9]_i_1__21_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__22 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank02/grn27/grn1__0 ),
        .O(\grn[9]_i_1__22_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__23 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn20/grn1__0 ),
        .O(\grn[9]_i_1__23_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__24 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn21/grn1__0 ),
        .O(\grn[9]_i_1__24_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__25 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn22/grn1__0 ),
        .O(\grn[9]_i_1__25_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__26 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn23/grn1__0 ),
        .O(\grn[9]_i_1__26_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__27 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn24/grn1__0 ),
        .O(\grn[9]_i_1__27_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__28 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn25/grn1__0 ),
        .O(\grn[9]_i_1__28_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__29 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn26/grn1__0 ),
        .O(\grn[9]_i_1__29_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__3 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn04/grn1__0 ),
        .O(\grn[9]_i_1__3_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \grn[9]_i_1__30 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/rgf_c1bus_0 [9]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c0bus_0 [9]),
        .I5(\rgf/bank13/grn27/grn1__0 ),
        .O(\grn[9]_i_1__30_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__4 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn05/grn1__0 ),
        .O(\grn[9]_i_1__4_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__5 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn06/grn1__0 ),
        .O(\grn[9]_i_1__5_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__6 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank02/grn07/grn1__0 ),
        .O(\grn[9]_i_1__6_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__7 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn07/grn1__0 ),
        .O(\grn[9]_i_1__7_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__8 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn05/grn1__0 ),
        .O(\grn[9]_i_1__8_n_0 ));
  LUT3 #(
    .INIT(8'hAC)) 
    \grn[9]_i_1__9 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/rgf_c0bus_0 [9]),
        .I2(\rgf/bank13/grn03/grn1__0 ),
        .O(\grn[9]_i_1__9_n_0 ));
  LUT4 #(
    .INIT(16'hE200)) 
    \ir0_id_fl[20]_i_1 
       (.I0(\fch/ir0_id_fl [20]),
        .I1(\fch/fch_term_fl ),
        .I2(\ir0_id_fl[20]_i_2_n_0 ),
        .I3(\fch/rst_n_fl ),
        .O(\ir0_id_fl[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEFAFAAAFF)) 
    \ir0_id_fl[20]_i_2 
       (.I0(\fch/fch_irq_req_fl ),
        .I1(\fch/nir_id [20]),
        .I2(\nir_id[20]_i_1_n_0 ),
        .I3(\ir0_id_fl[20]_i_3_n_0 ),
        .I4(\fch/fadr_1_fl ),
        .I5(fch_issu1_inferred_i_13_n_0),
        .O(\ir0_id_fl[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFFFAAAA)) 
    \ir0_id_fl[20]_i_3 
       (.I0(fdat[31]),
        .I1(\ir0_id_fl[20]_i_4_n_0 ),
        .I2(fdat[28]),
        .I3(fdat[26]),
        .I4(\ir0_id_fl[20]_i_5_n_0 ),
        .O(\ir0_id_fl[20]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hBBBAAAFB)) 
    \ir0_id_fl[20]_i_4 
       (.I0(\ir0_id_fl[20]_i_6_n_0 ),
        .I1(fdat[25]),
        .I2(fdat[23]),
        .I3(fdat[24]),
        .I4(fdat[27]),
        .O(\ir0_id_fl[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA2082AAAAAAAA)) 
    \ir0_id_fl[20]_i_5 
       (.I0(fch_issu1_inferred_i_88_n_0),
        .I1(fdat[17]),
        .I2(fdat[19]),
        .I3(fdat[16]),
        .I4(fdat[26]),
        .I5(\ir0_id_fl[20]_i_7_n_0 ),
        .O(\ir0_id_fl[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0020010000000100)) 
    \ir0_id_fl[20]_i_6 
       (.I0(fdat[21]),
        .I1(\ir0_id_fl[20]_i_8_n_0 ),
        .I2(fdat[22]),
        .I3(fdat[23]),
        .I4(fdat[20]),
        .I5(fdat[19]),
        .O(\ir0_id_fl[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \ir0_id_fl[20]_i_7 
       (.I0(fdat[24]),
        .I1(fdat[18]),
        .I2(fch_issu1_inferred_i_149_n_0),
        .I3(fdat[25]),
        .I4(fdat[29]),
        .I5(fch_issu1_inferred_i_138_n_0),
        .O(\ir0_id_fl[20]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ir0_id_fl[20]_i_8 
       (.I0(fdat[24]),
        .I1(fdat[27]),
        .O(\ir0_id_fl[20]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hEEE20000)) 
    \ir0_id_fl[21]_i_1 
       (.I0(\fch/ir0_id_fl [21]),
        .I1(\fch/fch_term_fl ),
        .I2(\ir0_id_fl[21]_i_2_n_0 ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/rst_n_fl ),
        .O(\ir0_id_fl[21]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \ir0_id_fl[21]_i_10 
       (.I0(fdat[22]),
        .I1(fdat[20]),
        .I2(fdat[21]),
        .O(\ir0_id_fl[21]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \ir0_id_fl[21]_i_11 
       (.I0(fdat[28]),
        .I1(fdat[18]),
        .I2(fdat[27]),
        .I3(fdat[26]),
        .O(\ir0_id_fl[21]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    \ir0_id_fl[21]_i_2 
       (.I0(\fch/nir_id [21]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/lir_id_0 [21]),
        .I4(\fch/fadr_1_fl ),
        .I5(\ir0_id_fl[21]_i_3_n_0 ),
        .O(\ir0_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000AEAEAE)) 
    \ir0_id_fl[21]_i_3 
       (.I0(\ir0_id_fl[21]_i_4_n_0 ),
        .I1(\ir0_id_fl[21]_i_5_n_0 ),
        .I2(\ir0_id_fl[21]_i_6_n_0 ),
        .I3(\ir0_id_fl[21]_i_7_n_0 ),
        .I4(\ir0_id_fl[21]_i_8_n_0 ),
        .I5(fdat[31]),
        .O(\ir0_id_fl[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h80C0CC0000000000)) 
    \ir0_id_fl[21]_i_4 
       (.I0(\ir0_id_fl[21]_i_9_n_0 ),
        .I1(fch_issu1_inferred_i_89_n_0),
        .I2(fdat[24]),
        .I3(fdat[26]),
        .I4(fdat[27]),
        .I5(fdat[25]),
        .O(\ir0_id_fl[21]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ir0_id_fl[21]_i_5 
       (.I0(fdat[24]),
        .I1(fdat[25]),
        .O(\ir0_id_fl[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7777FFF07777FFFF)) 
    \ir0_id_fl[21]_i_6 
       (.I0(fch_issu1_inferred_i_48_n_0),
        .I1(fch_issu1_inferred_i_89_n_0),
        .I2(\ir0_id_fl[21]_i_10_n_0 ),
        .I3(fch_issu1_inferred_i_76_n_0),
        .I4(fdat[23]),
        .I5(\ir0_id_fl[21]_i_11_n_0 ),
        .O(\ir0_id_fl[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ir0_id_fl[21]_i_7 
       (.I0(fdat[24]),
        .I1(fdat[18]),
        .I2(fdat[21]),
        .I3(fdat[20]),
        .I4(fdat[26]),
        .I5(fdat[25]),
        .O(\ir0_id_fl[21]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h41)) 
    \ir0_id_fl[21]_i_8 
       (.I0(fdat[16]),
        .I1(fdat[19]),
        .I2(fdat[17]),
        .O(\ir0_id_fl[21]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hCC028CC0)) 
    \ir0_id_fl[21]_i_9 
       (.I0(fdat[19]),
        .I1(fdat[22]),
        .I2(fdat[20]),
        .I3(fdat[21]),
        .I4(fdat[23]),
        .O(\ir0_id_fl[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_1
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_17_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [15]),
        .O(\fch/ir0 [15]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_10
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_26_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [6]),
        .O(\fch/ir0 [6]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_11
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_27_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [5]),
        .O(\fch/ir0 [5]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_12
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_28_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [4]),
        .O(\fch/ir0 [4]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_13
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_29_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [3]),
        .O(\fch/ir0 [3]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_14
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_30_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [2]),
        .O(\fch/ir0 [2]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_15
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_31_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [1]),
        .O(\fch/ir0 [1]));
  LUT6 #(
    .INIT(64'hAA08AA08AA080008)) 
    ir0_inferred_i_16
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir0_fl [0]),
        .I2(\fch/ctl_fetch0_fl ),
        .I3(\fch/fch_term_fl ),
        .I4(ir0_inferred_i_32_n_0),
        .I5(\fch/fch_irq_req_fl ),
        .O(\fch/ir0 [0]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_17
       (.I0(\fch/data0 [15]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[15]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[31]),
        .O(ir0_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_18
       (.I0(\fch/data0 [14]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[14]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[30]),
        .O(ir0_inferred_i_18_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_19
       (.I0(\fch/data0 [13]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[13]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[29]),
        .O(ir0_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_2
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_18_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [14]),
        .O(\fch/ir0 [14]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_20
       (.I0(\fch/data0 [12]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[12]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[28]),
        .O(ir0_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_21
       (.I0(\fch/data0 [11]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[11]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[27]),
        .O(ir0_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_22
       (.I0(\fch/data0 [10]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[10]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[26]),
        .O(ir0_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_23
       (.I0(\fch/data0 [9]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[9]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[25]),
        .O(ir0_inferred_i_23_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_24
       (.I0(\fch/data0 [8]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[8]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[24]),
        .O(ir0_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_25
       (.I0(\fch/data0 [7]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[7]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[23]),
        .O(ir0_inferred_i_25_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_26
       (.I0(\fch/data0 [6]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[6]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[22]),
        .O(ir0_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_27
       (.I0(\fch/data0 [5]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[5]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[21]),
        .O(ir0_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_28
       (.I0(\fch/data0 [4]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[4]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[20]),
        .O(ir0_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_29
       (.I0(\fch/data0 [3]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[3]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[19]),
        .O(ir0_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_3
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_19_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [13]),
        .O(\fch/ir0 [13]));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_30
       (.I0(\fch/data0 [2]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[2]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[18]),
        .O(ir0_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_31
       (.I0(\fch/data0 [1]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[1]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[17]),
        .O(ir0_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hFB08FBFBFB080808)) 
    ir0_inferred_i_32
       (.I0(\fch/data0 [0]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[0]),
        .I4(\fch/fadr_1_fl ),
        .I5(fdat[16]),
        .O(ir0_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_4
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_20_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [12]),
        .O(\fch/ir0 [12]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_5
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_21_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [11]),
        .O(\fch/ir0 [11]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_6
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_22_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [10]),
        .O(\fch/ir0 [10]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_7
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_23_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [9]),
        .O(\fch/ir0 [9]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_8
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_24_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [8]),
        .O(\fch/ir0 [8]));
  LUT6 #(
    .INIT(64'h00800A8A00800080)) 
    ir0_inferred_i_9
       (.I0(\fch/rst_n_fl ),
        .I1(ir0_inferred_i_25_n_0),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_irq_req_fl ),
        .I4(\fch/ctl_fetch0_fl ),
        .I5(\fch/ir0_fl [7]),
        .O(\fch/ir0 [7]));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[20]_i_1 
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir1_id_fl [20]),
        .I2(\fch/fch_term_fl ),
        .I3(\ir1_id_fl[20]_i_2_n_0 ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(\fch/fch_issu1 ),
        .O(fch_wrbufn1));
  LUT5 #(
    .INIT(32'hDDDDF0DD)) 
    \ir1_id_fl[20]_i_2 
       (.I0(\nir_id[20]_i_1_n_0 ),
        .I1(\fch/fadr_1_fl ),
        .I2(\ir0_id_fl[20]_i_3_n_0 ),
        .I3(\fch/stat [1]),
        .I4(\fch/stat [0]),
        .O(\ir1_id_fl[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h080808A808080808)) 
    \ir1_id_fl[21]_i_1 
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir1_id_fl [21]),
        .I2(\fch/fch_term_fl ),
        .I3(\ir1_id_fl[21]_i_2_n_0 ),
        .I4(\fch/fch_irq_req_fl ),
        .I5(\fch/fch_issu1 ),
        .O(fch_memacc1));
  LUT5 #(
    .INIT(32'hC5CCF5FF)) 
    \ir1_id_fl[21]_i_2 
       (.I0(\ir0_id_fl[21]_i_3_n_0 ),
        .I1(\fch/fadr_1_fl ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(\fch/lir_id_0 [21]),
        .O(\ir1_id_fl[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA000800080008)) 
    ir1_inferred_i_1
       (.I0(\fch/rst_n_fl ),
        .I1(\fch/ir1_fl [15]),
        .I2(\fch/ctl_fetch1_fl ),
        .I3(\fch/fch_term_fl ),
        .I4(ir1_inferred_i_17_n_0),
        .I5(ir1_inferred_i_18_n_0),
        .O(\fch/ir1 [15]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_10
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_27_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [6]),
        .O(\fch/ir1 [6]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_11
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_28_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [5]),
        .O(\fch/ir1 [5]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_12
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_29_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [4]),
        .O(\fch/ir1 [4]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_13
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_30_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [3]),
        .O(\fch/ir1 [3]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_14
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_31_n_0),
        .I2(\fch/ctl_fetch1_fl ),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/ir1_fl [2]),
        .O(\fch/ir1 [2]));
  LUT5 #(
    .INIT(32'h888A8888)) 
    ir1_inferred_i_15
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_32_n_0),
        .I2(\fch/ctl_fetch1_fl ),
        .I3(\fch/fch_term_fl ),
        .I4(\fch/ir1_fl [1]),
        .O(\fch/ir1 [1]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_16
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_33_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [0]),
        .O(\fch/ir1 [0]));
  LUT3 #(
    .INIT(8'h08)) 
    ir1_inferred_i_17
       (.I0(\fch/fch_issu1 ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_irq_req_fl ),
        .O(ir1_inferred_i_17_n_0));
  LUT5 #(
    .INIT(32'h0808FB08)) 
    ir1_inferred_i_18
       (.I0(fdat[31]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(fdat[15]),
        .I4(\fch/fadr_1_fl ),
        .O(ir1_inferred_i_18_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_19
       (.I0(fdat[30]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[14]),
        .O(ir1_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_2
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_19_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [14]),
        .O(\fch/ir1 [14]));
  LUT5 #(
    .INIT(32'hDD0DDDFD)) 
    ir1_inferred_i_20
       (.I0(fdat[13]),
        .I1(\fch/fadr_1_fl ),
        .I2(\fch/stat [1]),
        .I3(\fch/stat [0]),
        .I4(fdat[29]),
        .O(ir1_inferred_i_20_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_21
       (.I0(fdat[28]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[12]),
        .O(ir1_inferred_i_21_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_22
       (.I0(fdat[27]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[11]),
        .O(ir1_inferred_i_22_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_23
       (.I0(fdat[26]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[10]),
        .O(ir1_inferred_i_23_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_24
       (.I0(fdat[25]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[9]),
        .O(ir1_inferred_i_24_n_0));
  LUT5 #(
    .INIT(32'hC5CCF5FF)) 
    ir1_inferred_i_25
       (.I0(fdat[24]),
        .I1(\fch/fadr_1_fl ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(fdat[8]),
        .O(ir1_inferred_i_25_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_26
       (.I0(fdat[23]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[7]),
        .O(ir1_inferred_i_26_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_27
       (.I0(fdat[22]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[6]),
        .O(ir1_inferred_i_27_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_28
       (.I0(fdat[21]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[5]),
        .O(ir1_inferred_i_28_n_0));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_29
       (.I0(fdat[20]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[4]),
        .O(ir1_inferred_i_29_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_3
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_20_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [13]),
        .O(\fch/ir1 [13]));
  LUT5 #(
    .INIT(32'hF704F7F7)) 
    ir1_inferred_i_30
       (.I0(fdat[19]),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [0]),
        .I3(\fch/fadr_1_fl ),
        .I4(fdat[3]),
        .O(ir1_inferred_i_30_n_0));
  LUT6 #(
    .INIT(64'h40CC404040004040)) 
    ir1_inferred_i_31
       (.I0(\fch/fadr_1_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(fdat[2]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fdat[18]),
        .O(ir1_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'h40CC404040004040)) 
    ir1_inferred_i_32
       (.I0(\fch/fadr_1_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(fdat[1]),
        .I3(\fch/stat [0]),
        .I4(\fch/stat [1]),
        .I5(fdat[17]),
        .O(ir1_inferred_i_32_n_0));
  LUT5 #(
    .INIT(32'hC5CCF5FF)) 
    ir1_inferred_i_33
       (.I0(fdat[16]),
        .I1(\fch/fadr_1_fl ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(fdat[0]),
        .O(ir1_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_4
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_21_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [12]),
        .O(\fch/ir1 [12]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_5
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_22_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [11]),
        .O(\fch/ir1 [11]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_6
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_23_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [10]),
        .O(\fch/ir1 [10]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_7
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_24_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [9]),
        .O(\fch/ir1 [9]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_8
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_25_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [8]),
        .O(\fch/ir1 [8]));
  LUT6 #(
    .INIT(64'h080808AA08080808)) 
    ir1_inferred_i_9
       (.I0(\fch/rst_n_fl ),
        .I1(ir1_inferred_i_17_n_0),
        .I2(ir1_inferred_i_26_n_0),
        .I3(\fch/ctl_fetch1_fl ),
        .I4(\fch/fch_term_fl ),
        .I5(\fch/ir1_fl [7]),
        .O(\fch/ir1 [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [0]),
        .O(\rgf/ivec/p_1_in [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [10]),
        .O(\rgf/ivec/p_1_in [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [11]),
        .O(\rgf/ivec/p_1_in [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [12]),
        .O(\rgf/ivec/p_1_in [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [13]),
        .O(\rgf/ivec/p_1_in [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [14]),
        .O(\rgf/ivec/p_1_in [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [15]),
        .O(\rgf/ivec/p_1_in [15]));
  LUT4 #(
    .INIT(16'h0004)) 
    \iv[15]_i_2 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .I2(\iv[15]_i_4_n_0 ),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/c1bus_sel_cr [3]));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_3 
       (.I0(\grn[15]_i_3_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\pc[15]_i_11_n_0 ),
        .O(\rgf/c0bus_sel_cr [3]));
  LUT2 #(
    .INIT(4'h7)) 
    \iv[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\iv[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [1]),
        .O(\rgf/ivec/p_1_in [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [2]),
        .O(\rgf/ivec/p_1_in [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [3]),
        .O(\rgf/ivec/p_1_in [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [4]),
        .O(\rgf/ivec/p_1_in [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [5]),
        .O(\rgf/ivec/p_1_in [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [6]),
        .O(\rgf/ivec/p_1_in [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [7]),
        .O(\rgf/ivec/p_1_in [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [8]),
        .O(\rgf/ivec/p_1_in [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [3]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [3]),
        .I4(\rgf/ivec/iv [9]),
        .O(\rgf/ivec/p_1_in [9]));
  FDRE \mem/bctl/ctl/stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\stat[0]_i_1__2_n_0 ),
        .Q(\mem/bctl/ctl/p_0_in [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \mem/bctl/ctl/stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\mem/bctl/ctl/stat_nx ),
        .Q(\mem/bctl/ctl/p_0_in [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \mem/bctl/fch_term_fl_reg 
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_term),
        .Q(\mem/bctl/fch_term_fl ),
        .R(\<const0> ));
  FDRE \mem/bctl/read_cyc_reg[0] 
       (.C(clk),
        .CE(brdy),
        .D(badr[0]),
        .Q(\mem/read_cyc [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \mem/bctl/read_cyc_reg[1] 
       (.C(clk),
        .CE(brdy),
        .D(bcmd[2]),
        .Q(\mem/read_cyc [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \mem/bctl/read_cyc_reg[2] 
       (.C(clk),
        .CE(brdy),
        .D(bcmd[0]),
        .Q(\mem/read_cyc [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \mem/bctl/read_cyc_reg[3] 
       (.C(clk),
        .CE(brdy),
        .D(\mem/mem_accslot ),
        .Q(\mem/read_cyc [3]),
        .R(\alu1/div/p_0_in__0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \mul_a[15]_i_1 
       (.I0(rst_n),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\mul_a[15]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \mul_a[15]_i_1__0 
       (.I0(rst_n),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\mul_a[15]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[16]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[16]),
        .O(\mul_a[16]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[16]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[16]),
        .O(\mul_a[16]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[17]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[17]),
        .O(\alu0/mul_a_i [17]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[17]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[17]),
        .O(\alu1/mul_a_i [17]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[18]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[18]),
        .O(\alu0/mul_a_i [18]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[18]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[18]),
        .O(\alu1/mul_a_i [18]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[19]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[19]),
        .O(\alu0/mul_a_i [19]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[19]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[19]),
        .O(\alu1/mul_a_i [19]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[20]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[20]),
        .O(\alu0/mul_a_i [20]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[20]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[20]),
        .O(\alu1/mul_a_i [20]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[21]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[21]),
        .O(\alu0/mul_a_i [21]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[21]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[21]),
        .O(\alu1/mul_a_i [21]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[22]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[22]),
        .O(\alu0/mul_a_i [22]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[22]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[22]),
        .O(\alu1/mul_a_i [22]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[23]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[23]),
        .O(\alu0/mul_a_i [23]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[23]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[23]),
        .O(\alu1/mul_a_i [23]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[24]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[24]),
        .O(\alu0/mul_a_i [24]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[24]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[24]),
        .O(\alu1/mul_a_i [24]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[25]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[25]),
        .O(\alu0/mul_a_i [25]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[25]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[25]),
        .O(\alu1/mul_a_i [25]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[26]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[26]),
        .O(\alu0/mul_a_i [26]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[26]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[26]),
        .O(\alu1/mul_a_i [26]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[27]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[27]),
        .O(\alu0/mul_a_i [27]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[27]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[27]),
        .O(\alu1/mul_a_i [27]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[28]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[28]),
        .O(\alu0/mul_a_i [28]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[28]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[28]),
        .O(\alu1/mul_a_i [28]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[29]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[29]),
        .O(\alu0/mul_a_i [29]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[29]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[29]),
        .O(\alu1/mul_a_i [29]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[30]_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[30]),
        .O(\alu0/mul_a_i [30]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[30]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[30]),
        .O(\alu1/mul_a_i [30]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[31]_i_1 
       (.I0(\alu1/mul_a_i [31]),
        .I1(rst_n),
        .O(\mul_a[31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_a[31]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(rst_n),
        .O(\mul_a[31]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_a[32]_i_1 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(rst_n),
        .I2(\alu1/mul_a_i [31]),
        .O(\mul_a[32]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_a[32]_i_1__0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(rst_n),
        .O(\mul_a[32]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[32]_i_2 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[31]),
        .O(\alu1/mul_a_i [31]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[0]_i_1 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(b1bus_0[0]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[0]_i_1__0 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(b0bus_0[0]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[1]_i_1 
       (.I0(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .O(b1bus_0[1]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[1]_i_1__0 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(b0bus_0[1]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[2]_i_1 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .O(b1bus_0[2]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[2]_i_1__0 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(b0bus_0[2]));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_b[31]_i_1 
       (.I0(b0bus_0[31]),
        .I1(rst_n),
        .I2(\rgf/sreg/sr [8]),
        .O(\mul_b[31]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_b[31]_i_1__0 
       (.I0(b1bus_0[31]),
        .I1(rst_n),
        .I2(\rgf/sreg/sr [8]),
        .O(\mul_b[31]_i_1__0_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_b[32]_i_1 
       (.I0(b0bus_0[31]),
        .I1(rst_n),
        .I2(\rgf/sreg/sr [8]),
        .I3(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .O(\mul_b[32]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_b[32]_i_1__0 
       (.I0(b1bus_0[31]),
        .I1(rst_n),
        .I2(\rgf/sreg/sr [8]),
        .I3(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .O(\mul_b[32]_i_1__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[3]_i_1 
       (.I0(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .O(b1bus_0[3]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[3]_i_1__0 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(b0bus_0[3]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[4]_i_1 
       (.I0(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(b1bus_0[4]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[4]_i_1__0 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(b0bus_0[4]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[5]_i_1 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(b1bus_0[5]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[5]_i_1__0 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(b0bus_0[5]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[6]_i_1 
       (.I0(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .O(b1bus_0[6]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[6]_i_1__0 
       (.I0(\bbus_o[6]_INST_0_i_1_n_0 ),
        .O(b0bus_0[6]));
  LUT2 #(
    .INIT(4'h2)) 
    mul_rslt_i_1
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .O(\alu0/mul/mul_rslt0 ));
  LUT2 #(
    .INIT(4'h2)) 
    mul_rslt_i_1__0
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .O(\alu1/mul/mul_rslt0 ));
  LUT3 #(
    .INIT(8'h75)) 
    \mulh[15]_i_1 
       (.I0(rst_n),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\mulh[15]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h75)) 
    \mulh[15]_i_1__0 
       (.I0(rst_n),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\mulh[15]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \mulh[15]_i_2 
       (.I0(rst_n),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .O(\alu0/mul/mul_b ));
  LUT2 #(
    .INIT(4'h7)) 
    \mulh[15]_i_2__0 
       (.I0(rst_n),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .O(\alu1/mul/mul_b ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[12]_i_1 
       (.I0(\nir_id[12]_i_2_n_0 ),
        .O(\fch/lir_id_0 [12]));
  LUT6 #(
    .INIT(64'hBFBFFFBFAAAAAAAA)) 
    \nir_id[12]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[12]_i_3_n_0 ),
        .I2(fdat[14]),
        .I3(\nir_id[14]_i_5_n_0 ),
        .I4(\nir_id[12]_i_4_n_0 ),
        .I5(\nir_id[14]_i_7_n_0 ),
        .O(\nir_id[12]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAEAAA)) 
    \nir_id[12]_i_3 
       (.I0(\nir_id[14]_i_8_n_0 ),
        .I1(fdat[0]),
        .I2(fdat[8]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .O(\nir_id[12]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hA008AA08AAA8AAA8)) 
    \nir_id[12]_i_4 
       (.I0(fdat[10]),
        .I1(fdat[0]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[12]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[13]_i_1 
       (.I0(\nir_id[13]_i_2_n_0 ),
        .O(\fch/lir_id_0 [13]));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAABFBB)) 
    \nir_id[13]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[13]_i_3_n_0 ),
        .I2(\nir_id[13]_i_4_n_0 ),
        .I3(\nir_id[14]_i_5_n_0 ),
        .I4(fdat[15]),
        .I5(\nir_id[13]_i_5_n_0 ),
        .O(\nir_id[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAEAAFAAAFAAA)) 
    \nir_id[13]_i_3 
       (.I0(\nir_id[13]_i_6_n_0 ),
        .I1(fdat[1]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(\nir_id[13]_i_7_n_0 ),
        .I5(fdat[10]),
        .O(\nir_id[13]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hA20AAAAAA200AAA0)) 
    \nir_id[13]_i_4 
       (.I0(fdat[10]),
        .I1(fdat[6]),
        .I2(fdat[9]),
        .I3(fdat[8]),
        .I4(fdat[7]),
        .I5(fdat[1]),
        .O(\nir_id[13]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[13]_i_5 
       (.I0(fdat[14]),
        .I1(fdat[13]),
        .O(\nir_id[13]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[13]_i_6 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .O(\nir_id[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7CEFFFF)) 
    \nir_id[13]_i_7 
       (.I0(fdat[6]),
        .I1(fdat[5]),
        .I2(fdat[3]),
        .I3(fdat[4]),
        .I4(\nir_id[13]_i_8_n_0 ),
        .I5(\nir_id[13]_i_9_n_0 ),
        .O(\nir_id[13]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \nir_id[13]_i_8 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .O(\nir_id[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h08880880FFFFFFFF)) 
    \nir_id[13]_i_9 
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[6]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fdat[9]),
        .O(\nir_id[13]_i_9_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[14]_i_1 
       (.I0(\nir_id[14]_i_2_n_0 ),
        .O(\fch/lir_id_0 [14]));
  LUT3 #(
    .INIT(8'h09)) 
    \nir_id[14]_i_10 
       (.I0(fdat[3]),
        .I1(fdat[1]),
        .I2(fdat[0]),
        .O(\nir_id[14]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \nir_id[14]_i_11 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .I2(fdat[10]),
        .O(\nir_id[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AAA8A8A882)) 
    \nir_id[14]_i_12 
       (.I0(fdat[8]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(fdat[3]),
        .O(\nir_id[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBFBFFFBFAAAAAAAA)) 
    \nir_id[14]_i_2 
       (.I0(\nir_id[14]_i_3_n_0 ),
        .I1(\nir_id[14]_i_4_n_0 ),
        .I2(fdat[14]),
        .I3(\nir_id[14]_i_5_n_0 ),
        .I4(\nir_id[14]_i_6_n_0 ),
        .I5(\nir_id[14]_i_7_n_0 ),
        .O(\nir_id[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00B0F030)) 
    \nir_id[14]_i_3 
       (.I0(fdat[11]),
        .I1(fdat[14]),
        .I2(fdat[15]),
        .I3(fdat[13]),
        .I4(fdat[12]),
        .O(\nir_id[14]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBAAAAAAEAAAAA)) 
    \nir_id[14]_i_4 
       (.I0(\nir_id[14]_i_8_n_0 ),
        .I1(fdat[8]),
        .I2(fdat[2]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(fdat[7]),
        .O(\nir_id[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA00002000)) 
    \nir_id[14]_i_5 
       (.I0(\nir_id[14]_i_9_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[9]),
        .I3(fdat[7]),
        .I4(fdat[8]),
        .I5(fdat[10]),
        .O(\nir_id[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hA2A0AAA8AAA8AAA8)) 
    \nir_id[14]_i_6 
       (.I0(fdat[10]),
        .I1(fdat[8]),
        .I2(fdat[9]),
        .I3(fdat[2]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0A000A030A000A00)) 
    \nir_id[14]_i_7 
       (.I0(fdat[13]),
        .I1(\nir_id[14]_i_10_n_0 ),
        .I2(fdat[15]),
        .I3(fdat[14]),
        .I4(\nir_id[14]_i_11_n_0 ),
        .I5(\nir_id[20]_i_5_n_0 ),
        .O(\nir_id[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h3FFF3F3FBFBF3F3F)) 
    \nir_id[14]_i_8 
       (.I0(fdat[8]),
        .I1(fdat[12]),
        .I2(fdat[11]),
        .I3(\nir_id[14]_i_12_n_0 ),
        .I4(fdat[9]),
        .I5(fdat[10]),
        .O(\nir_id[14]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \nir_id[14]_i_9 
       (.I0(fdat[12]),
        .I1(fdat[11]),
        .O(\nir_id[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hF6FFFFFFFFFFFFFF)) 
    \nir_id[15]_i_1 
       (.I0(fdat[8]),
        .I1(fdat[11]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(fdat[12]),
        .I5(\nir_id[15]_i_2_n_0 ),
        .O(\fch/lir_id_0 [15]));
  LUT3 #(
    .INIT(8'h40)) 
    \nir_id[15]_i_2 
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .O(\nir_id[15]_i_2_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[16]_i_1 
       (.I0(\nir_id[16]_i_2_n_0 ),
        .O(\fch/lir_id_0 [16]));
  LUT6 #(
    .INIT(64'h111F111111111111)) 
    \nir_id[16]_i_2 
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(fdat[8]),
        .I2(\nir_id[16]_i_3_n_0 ),
        .I3(fdat[15]),
        .I4(fdat[13]),
        .I5(fdat[14]),
        .O(\nir_id[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hA8AAAAAA)) 
    \nir_id[16]_i_3 
       (.I0(\nir_id[16]_i_4_n_0 ),
        .I1(fdat[3]),
        .I2(fdat[11]),
        .I3(fdat[12]),
        .I4(\nir_id[17]_i_6_n_0 ),
        .O(\nir_id[16]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFD000)) 
    \nir_id[16]_i_4 
       (.I0(\nir_id[18]_i_6_n_0 ),
        .I1(fdat[0]),
        .I2(fdat[9]),
        .I3(fdat[10]),
        .I4(\nir_id[16]_i_5_n_0 ),
        .I5(\nir_id[17]_i_7_n_0 ),
        .O(\nir_id[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h5CDCFFFFFFFFFFFF)) 
    \nir_id[16]_i_5 
       (.I0(\nir_id[16]_i_6_n_0 ),
        .I1(fdat[3]),
        .I2(fdat[10]),
        .I3(fdat[9]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[16]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \nir_id[16]_i_6 
       (.I0(fdat[9]),
        .I1(fdat[8]),
        .I2(fdat[6]),
        .I3(fdat[7]),
        .O(\nir_id[16]_i_6_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[17]_i_1 
       (.I0(\nir_id[17]_i_2_n_0 ),
        .O(\fch/lir_id_0 [17]));
  LUT6 #(
    .INIT(64'hAAAABBABAAAAAAAB)) 
    \nir_id[17]_i_2 
       (.I0(\nir_id[17]_i_3_n_0 ),
        .I1(\nir_id[17]_i_4_n_0 ),
        .I2(fdat[4]),
        .I3(\nir_id[21]_i_9_n_0 ),
        .I4(fdat[15]),
        .I5(\nir_id[17]_i_5_n_0 ),
        .O(\nir_id[17]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0551555500000000)) 
    \nir_id[17]_i_3 
       (.I0(fdat[9]),
        .I1(fdat[11]),
        .I2(fdat[12]),
        .I3(fdat[14]),
        .I4(fdat[13]),
        .I5(fdat[15]),
        .O(\nir_id[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF3FFF7FFF7FFF)) 
    \nir_id[17]_i_4 
       (.I0(\nir_id[17]_i_6_n_0 ),
        .I1(fdat[12]),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .I4(\nir_id[17]_i_7_n_0 ),
        .I5(fdat[11]),
        .O(\nir_id[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h03A303A303A300A0)) 
    \nir_id[17]_i_5 
       (.I0(\nir_id[18]_i_6_n_0 ),
        .I1(fdat[4]),
        .I2(fdat[9]),
        .I3(fdat[1]),
        .I4(fdat[8]),
        .I5(\nir_id[18]_i_7_n_0 ),
        .O(\nir_id[17]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h0A5BD5FF)) 
    \nir_id[17]_i_6 
       (.I0(fdat[10]),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[9]),
        .O(\nir_id[17]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h30002020)) 
    \nir_id[17]_i_7 
       (.I0(fdat[7]),
        .I1(fdat[10]),
        .I2(fdat[9]),
        .I3(fdat[6]),
        .I4(fdat[8]),
        .O(\nir_id[17]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[18]_i_1 
       (.I0(\nir_id[18]_i_2_n_0 ),
        .O(\fch/lir_id_0 [18]));
  LUT6 #(
    .INIT(64'hD1FF1111113F1111)) 
    \nir_id[18]_i_2 
       (.I0(\nir_id[18]_i_3_n_0 ),
        .I1(fdat[10]),
        .I2(fdat[11]),
        .I3(fdat[5]),
        .I4(\nir_id[18]_i_4_n_0 ),
        .I5(\nir_id[18]_i_5_n_0 ),
        .O(\nir_id[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hD55DD555)) 
    \nir_id[18]_i_3 
       (.I0(fdat[15]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .I3(fdat[12]),
        .I4(fdat[11]),
        .O(\nir_id[18]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[18]_i_4 
       (.I0(fdat[15]),
        .I1(\nir_id[17]_i_4_n_0 ),
        .O(\nir_id[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h202F202F202F2020)) 
    \nir_id[18]_i_5 
       (.I0(\nir_id[18]_i_6_n_0 ),
        .I1(fdat[2]),
        .I2(fdat[9]),
        .I3(fdat[5]),
        .I4(fdat[8]),
        .I5(\nir_id[18]_i_7_n_0 ),
        .O(\nir_id[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8C804880CC000C04)) 
    \nir_id[18]_i_6 
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[5]),
        .I3(fdat[6]),
        .I4(fdat[3]),
        .I5(fdat[4]),
        .O(\nir_id[18]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \nir_id[18]_i_7 
       (.I0(fdat[7]),
        .I1(fdat[6]),
        .O(\nir_id[18]_i_7_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \nir_id[19]_i_1 
       (.I0(\nir_id[19]_i_2_n_0 ),
        .O(\fch/lir_id_0 [19]));
  LUT6 #(
    .INIT(64'hAEEEEAAEAAEEEEEE)) 
    \nir_id[19]_i_2 
       (.I0(\nir_id[19]_i_3_n_0 ),
        .I1(fdat[15]),
        .I2(fdat[13]),
        .I3(fdat[14]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[19]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0222222222222222)) 
    \nir_id[19]_i_3 
       (.I0(\nir_id[18]_i_4_n_0 ),
        .I1(\nir_id[19]_i_4_n_0 ),
        .I2(\nir_id[19]_i_5_n_0 ),
        .I3(\nir_id[19]_i_6_n_0 ),
        .I4(\nir_id[19]_i_7_n_0 ),
        .I5(fdat[11]),
        .O(\nir_id[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0020010000000000)) 
    \nir_id[19]_i_4 
       (.I0(fdat[7]),
        .I1(fdat[9]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[10]),
        .I5(fdat[11]),
        .O(\nir_id[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF77FF77F77FFF7FF)) 
    \nir_id[19]_i_5 
       (.I0(fdat[7]),
        .I1(fdat[8]),
        .I2(fdat[5]),
        .I3(fdat[6]),
        .I4(fdat[3]),
        .I5(fdat[4]),
        .O(\nir_id[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFDFFFFFFFDDFD)) 
    \nir_id[19]_i_6 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[3]),
        .I3(fdat[6]),
        .I4(fdat[5]),
        .I5(fdat[4]),
        .O(\nir_id[19]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[19]_i_7 
       (.I0(fdat[9]),
        .I1(fdat[10]),
        .O(\nir_id[19]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h44445444)) 
    \nir_id[20]_i_1 
       (.I0(fdat[15]),
        .I1(\nir_id[20]_i_2_n_0 ),
        .I2(fdat[12]),
        .I3(fdat[10]),
        .I4(\nir_id[20]_i_3_n_0 ),
        .O(\nir_id[20]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEFBEAAAAAAAA)) 
    \nir_id[20]_i_2 
       (.I0(\nir_id[20]_i_4_n_0 ),
        .I1(fdat[1]),
        .I2(fdat[3]),
        .I3(fdat[0]),
        .I4(fdat[10]),
        .I5(\nir_id[20]_i_5_n_0 ),
        .O(\nir_id[20]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAFFFFEE)) 
    \nir_id[20]_i_3 
       (.I0(\nir_id[20]_i_6_n_0 ),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[5]),
        .I4(fdat[4]),
        .I5(\nir_id[20]_i_7_n_0 ),
        .O(\nir_id[20]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h7776)) 
    \nir_id[20]_i_4 
       (.I0(fdat[14]),
        .I1(fdat[13]),
        .I2(fdat[12]),
        .I3(fdat[11]),
        .O(\nir_id[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \nir_id[20]_i_5 
       (.I0(fdat[13]),
        .I1(fdat[7]),
        .I2(fdat[2]),
        .I3(\nir_id[20]_i_8_n_0 ),
        .I4(fdat[8]),
        .I5(fdat[9]),
        .O(\nir_id[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h11F1FFFFFFFFFFFF)) 
    \nir_id[20]_i_6 
       (.I0(fdat[6]),
        .I1(fdat[7]),
        .I2(fdat[4]),
        .I3(fdat[3]),
        .I4(fdat[8]),
        .I5(fdat[11]),
        .O(\nir_id[20]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0E45)) 
    \nir_id[20]_i_7 
       (.I0(fdat[8]),
        .I1(fdat[7]),
        .I2(fdat[9]),
        .I3(fdat[11]),
        .O(\nir_id[20]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \nir_id[20]_i_8 
       (.I0(fdat[6]),
        .I1(fdat[4]),
        .I2(fdat[5]),
        .O(\nir_id[20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AAAB)) 
    \nir_id[21]_i_1 
       (.I0(\nir_id[21]_i_2_n_0 ),
        .I1(fdat[9]),
        .I2(fdat[8]),
        .I3(\nir_id[21]_i_3_n_0 ),
        .I4(\nir_id[21]_i_4_n_0 ),
        .I5(fdat[15]),
        .O(\fch/lir_id_0 [21]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \nir_id[21]_i_10 
       (.I0(fdat[4]),
        .I1(fdat[5]),
        .I2(fdat[2]),
        .I3(fdat[8]),
        .O(\nir_id[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8FC0000000000000)) 
    \nir_id[21]_i_2 
       (.I0(\nir_id[21]_i_5_n_0 ),
        .I1(fdat[8]),
        .I2(fdat[11]),
        .I3(fdat[10]),
        .I4(\nir_id[21]_i_6_n_0 ),
        .I5(fdat[9]),
        .O(\nir_id[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00DFDFDFDFDFDFDF)) 
    \nir_id[21]_i_3 
       (.I0(\nir_id[21]_i_7_n_0 ),
        .I1(fdat[14]),
        .I2(\nir_id[21]_i_8_n_0 ),
        .I3(fdat[7]),
        .I4(\nir_id[21]_i_9_n_0 ),
        .I5(\nir_id[21]_i_6_n_0 ),
        .O(\nir_id[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000041)) 
    \nir_id[21]_i_4 
       (.I0(fdat[0]),
        .I1(fdat[1]),
        .I2(fdat[3]),
        .I3(fdat[9]),
        .I4(fdat[10]),
        .I5(\nir_id[21]_i_10_n_0 ),
        .O(\nir_id[21]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hC8CC0C20)) 
    \nir_id[21]_i_5 
       (.I0(fdat[3]),
        .I1(fdat[6]),
        .I2(fdat[7]),
        .I3(fdat[4]),
        .I4(fdat[5]),
        .O(\nir_id[21]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \nir_id[21]_i_6 
       (.I0(fdat[12]),
        .I1(fdat[13]),
        .I2(fdat[14]),
        .O(\nir_id[21]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \nir_id[21]_i_7 
       (.I0(fdat[2]),
        .I1(fdat[7]),
        .I2(fdat[13]),
        .O(\nir_id[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \nir_id[21]_i_8 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .I2(fdat[6]),
        .I3(fdat[10]),
        .I4(fdat[11]),
        .I5(fdat[12]),
        .O(\nir_id[21]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \nir_id[21]_i_9 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .O(\nir_id[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h8A888A888A888A8A)) 
    \nir_id[24]_i_1 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\nir_id[24]_i_3_n_0 ),
        .I2(\nir_id[24]_i_4_n_0 ),
        .I3(\nir_id[24]_i_5_n_0 ),
        .I4(\nir_id[24]_i_6_n_0 ),
        .I5(\nir_id[24]_i_7_n_0 ),
        .O(\fch/fctl/fch_nir_lir ));
  LUT6 #(
    .INIT(64'h0000000000008002)) 
    \nir_id[24]_i_10 
       (.I0(\nir_id[24]_i_16_n_0 ),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [12]),
        .I4(\nir_id[24]_i_17_n_0 ),
        .I5(\nir_id[24]_i_18_n_0 ),
        .O(ctl_fetch_ext1));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_11 
       (.I0(fdat[8]),
        .I1(fdat[9]),
        .O(\nir_id[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFEAAAAABAAAAAAAA)) 
    \nir_id[24]_i_12 
       (.I0(\nir_id[24]_i_19_n_0 ),
        .I1(fdat[7]),
        .I2(fdat[6]),
        .I3(fdat[10]),
        .I4(fdat[9]),
        .I5(\nir_id[24]_i_20_n_0 ),
        .O(\nir_id[24]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000C1C00001C0C0)) 
    \nir_id[24]_i_13 
       (.I0(\bdatw[8]_INST_0_i_21_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [6]),
        .I3(stat[2]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [0]),
        .O(\nir_id[24]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFFFFFFFFFFFFE)) 
    \nir_id[24]_i_14 
       (.I0(\bdatw[31]_INST_0_i_79_n_0 ),
        .I1(stat[1]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [8]),
        .O(\nir_id[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDFFADFFFFFFA)) 
    \nir_id[24]_i_15 
       (.I0(\fch/ir0 [12]),
        .I1(stat[2]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [11]),
        .I4(stat[0]),
        .I5(\rgf/sreg/sr [9]),
        .O(\nir_id[24]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0F0000000F000018)) 
    \nir_id[24]_i_16 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [6]),
        .I5(\bdatw[9]_INST_0_i_10_n_0 ),
        .O(\nir_id[24]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBFFFFFFFFFFB)) 
    \nir_id[24]_i_17 
       (.I0(\fch/ir1 [4]),
        .I1(\fch_irq_lev[1]_i_8_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [10]),
        .I4(\nir_id[24]_i_21_n_0 ),
        .I5(\fch/ir1 [8]),
        .O(\nir_id[24]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDFFADFFFFFFA)) 
    \nir_id[24]_i_18 
       (.I0(\fch/ir1 [12]),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [11]),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\rgf/sreg/sr [9]),
        .O(\nir_id[24]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0F0000010F000000)) 
    \nir_id[24]_i_19 
       (.I0(\nir_id[24]_i_22_n_0 ),
        .I1(fdat[13]),
        .I2(\nir_id[24]_i_23_n_0 ),
        .I3(fdat[7]),
        .I4(fdat[12]),
        .I5(\nir_id[24]_i_24_n_0 ),
        .O(\nir_id[24]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h003C000055FFFFFD)) 
    \nir_id[24]_i_2 
       (.I0(\nir_id[24]_i_8_n_0 ),
        .I1(fdat[11]),
        .I2(fdat[12]),
        .I3(fdat[13]),
        .I4(fdat[14]),
        .I5(fdat[15]),
        .O(\fch/lir_id_0 [24]));
  LUT6 #(
    .INIT(64'h000000008B778BFF)) 
    \nir_id[24]_i_20 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .I2(fdat[7]),
        .I3(fdat[6]),
        .I4(fdat[9]),
        .I5(\nir_id[24]_i_25_n_0 ),
        .O(\nir_id[24]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_21 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .O(\nir_id[24]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \nir_id[24]_i_22 
       (.I0(fdat[5]),
        .I1(fdat[4]),
        .O(\nir_id[24]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFEFE)) 
    \nir_id[24]_i_23 
       (.I0(fdat[10]),
        .I1(fdat[11]),
        .I2(fdat[8]),
        .I3(fdat[9]),
        .I4(fdat[6]),
        .I5(fdat[7]),
        .O(\nir_id[24]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_24 
       (.I0(fdat[2]),
        .I1(fdat[9]),
        .O(\nir_id[24]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h60FFFFFFFFFFFFFF)) 
    \nir_id[24]_i_25 
       (.I0(fdat[3]),
        .I1(fdat[5]),
        .I2(fdat[6]),
        .I3(fdat[8]),
        .I4(fdat[12]),
        .I5(fdat[11]),
        .O(\nir_id[24]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000030C0C03939)) 
    \nir_id[24]_i_3 
       (.I0(\fch/fch_issu1_ir ),
        .I1(\fch/stat [1]),
        .I2(\fch/stat [2]),
        .I3(fch_leir_nir_i_2_n_0),
        .I4(\fch/stat [0]),
        .I5(\fadr[15]_INST_0_i_16_n_0 ),
        .O(\nir_id[24]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \nir_id[24]_i_4 
       (.I0(fch_term),
        .I1(\fch/stat [2]),
        .I2(\fch/stat [0]),
        .O(\nir_id[24]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h45401015)) 
    \nir_id[24]_i_5 
       (.I0(fch_heir_nir_i_3_n_0),
        .I1(\fch/fch_issu1 ),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_issu1_fl ),
        .I4(\fch/stat [1]),
        .O(\nir_id[24]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \nir_id[24]_i_6 
       (.I0(ctl_fetch_ext0),
        .I1(ctl_fetch_ext1),
        .O(\nir_id[24]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \nir_id[24]_i_7 
       (.I0(\fch/fch_issu1_fl ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_issu1 ),
        .I3(\fch/stat [1]),
        .O(\nir_id[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h01000001FFFFFFFF)) 
    \nir_id[24]_i_8 
       (.I0(fdat[4]),
        .I1(\nir_id[24]_i_11_n_0 ),
        .I2(fdat[1]),
        .I3(fdat[0]),
        .I4(fdat[3]),
        .I5(\nir_id[24]_i_12_n_0 ),
        .O(\nir_id[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008002)) 
    \nir_id[24]_i_9 
       (.I0(\nir_id[24]_i_13_n_0 ),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [12]),
        .I4(\nir_id[24]_i_14_n_0 ),
        .I5(\nir_id[24]_i_15_n_0 ),
        .O(ctl_fetch_ext0));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[0]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[0]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [0]),
        .O(niss_dsp_a0[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[10]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [10]),
        .O(niss_dsp_a0[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[11]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [11]),
        .O(niss_dsp_a0[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[12]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [12]),
        .O(niss_dsp_a0[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[13]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [13]),
        .O(niss_dsp_a0[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[14]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[14]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [14]),
        .O(niss_dsp_a0[14]));
  LUT5 #(
    .INIT(32'h80FF8080)) 
    \niss_dsp_a0[15]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu0/mul/mul_rslt ),
        .I2(\alu0/mul/mul_a [15]),
        .I3(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .O(niss_dsp_a0[15]));
  LUT4 #(
    .INIT(16'hFD7F)) 
    \niss_dsp_a0[15]_INST_0_i_1 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\niss_dsp_a0[15]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[16]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [16]),
        .O(niss_dsp_a0[16]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[17]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [17]),
        .O(niss_dsp_a0[17]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[18]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [18]),
        .O(niss_dsp_a0[18]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[19]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [19]),
        .O(niss_dsp_a0[19]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[1]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [1]),
        .O(niss_dsp_a0[1]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[20]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [20]),
        .O(niss_dsp_a0[20]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[21]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [21]),
        .O(niss_dsp_a0[21]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[22]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [22]),
        .O(niss_dsp_a0[22]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[23]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [23]),
        .O(niss_dsp_a0[23]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[24]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [24]),
        .O(niss_dsp_a0[24]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[25]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [25]),
        .O(niss_dsp_a0[25]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[26]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [26]),
        .O(niss_dsp_a0[26]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[27]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [27]),
        .O(niss_dsp_a0[27]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[28]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [28]),
        .O(niss_dsp_a0[28]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[29]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [29]),
        .O(niss_dsp_a0[29]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[2]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [2]),
        .O(niss_dsp_a0[2]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[30]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [30]),
        .O(niss_dsp_a0[30]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[31]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [31]),
        .O(niss_dsp_a0[31]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a0[32]_INST_0 
       (.I0(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [32]),
        .O(niss_dsp_a0[32]));
  LUT4 #(
    .INIT(16'h1000)) 
    \niss_dsp_a0[32]_INST_0_i_1 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hD3)) 
    \niss_dsp_a0[32]_INST_0_i_10 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .O(\niss_dsp_a0[32]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    \niss_dsp_a0[32]_INST_0_i_11 
       (.I0(\rgf_selc0_wb[1]_i_15_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [11]),
        .I3(\niss_dsp_a0[32]_INST_0_i_12_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_13_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_14_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF0FFF7F0070)) 
    \niss_dsp_a0[32]_INST_0_i_12 
       (.I0(crdy),
        .I1(div_crdy0),
        .I2(\fch/ir0 [7]),
        .I3(stat[1]),
        .I4(stat[0]),
        .I5(\fch/ir0 [8]),
        .O(\niss_dsp_a0[32]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF282A2A2A)) 
    \niss_dsp_a0[32]_INST_0_i_13 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(ctl_fetch0_fl_i_28_n_0),
        .I4(\fch/ir0 [9]),
        .I5(\niss_dsp_a0[32]_INST_0_i_15_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0080888A0000880A)) 
    \niss_dsp_a0[32]_INST_0_i_14 
       (.I0(\rgf_selc0_rn_wb[2]_i_26_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(stat[1]),
        .I4(stat[0]),
        .I5(\ccmd[2]_INST_0_i_10_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \niss_dsp_a0[32]_INST_0_i_15 
       (.I0(ctl_fetch0_fl_i_40_n_0),
        .I1(\fch/ir0 [8]),
        .I2(stat[0]),
        .I3(\ccmd[2]_INST_0_i_9_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\niss_dsp_a0[32]_INST_0_i_16_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \niss_dsp_a0[32]_INST_0_i_16 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [4]),
        .O(\niss_dsp_a0[32]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a0[32]_INST_0_i_2 
       (.I0(a0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .O(\niss_dsp_a0[32]_INST_0_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_3 
       (.I0(ccmd[4]),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_4 
       (.I0(ccmd[4]),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a0[32]_INST_0_i_5 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_6 
       (.I0(ccmd[4]),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0010001000001111)) 
    \niss_dsp_a0[32]_INST_0_i_7 
       (.I0(ccmd[4]),
        .I1(\niss_dsp_a0[32]_INST_0_i_9_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_10_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_11_n_0 ),
        .I5(\fch/ir0 [15]),
        .O(\niss_dsp_a0[32]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a0[32]_INST_0_i_8 
       (.I0(ccmd[4]),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(\niss_dsp_a0[32]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4F5F4FFF5FFF5FFF)) 
    \niss_dsp_a0[32]_INST_0_i_9 
       (.I0(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I1(stat[2]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [12]),
        .O(\niss_dsp_a0[32]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[3]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [3]),
        .O(niss_dsp_a0[3]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[4]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [4]),
        .O(niss_dsp_a0[4]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[5]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [5]),
        .O(niss_dsp_a0[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[6]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [6]),
        .O(niss_dsp_a0[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[7]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [7]),
        .O(niss_dsp_a0[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[8]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [8]),
        .O(niss_dsp_a0[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a0[9]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_a [9]),
        .O(niss_dsp_a0[9]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[0]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [0]),
        .O(niss_dsp_a1[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[10]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[10]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [10]),
        .O(niss_dsp_a1[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[11]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[11]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [11]),
        .O(niss_dsp_a1[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[12]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [12]),
        .O(niss_dsp_a1[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[13]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[13]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [13]),
        .O(niss_dsp_a1[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[14]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[14]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [14]),
        .O(niss_dsp_a1[14]));
  LUT5 #(
    .INIT(32'h80FF8080)) 
    \niss_dsp_a1[15]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu1/mul/mul_rslt ),
        .I2(\alu1/mul/mul_a [15]),
        .I3(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(niss_dsp_a1[15]));
  LUT4 #(
    .INIT(16'h070F)) 
    \niss_dsp_a1[15]_INST_0_i_1 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(acmd1[0]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hC000000000000080)) 
    \niss_dsp_a1[15]_INST_0_i_10 
       (.I0(\fch/ir1 [7]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\niss_dsp_a1[15]_INST_0_i_22_n_0 ),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [6]),
        .O(\niss_dsp_a1[15]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h44114F1100000000)) 
    \niss_dsp_a1[15]_INST_0_i_11 
       (.I0(\fch/ir1 [14]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\niss_dsp_a1[15]_INST_0_i_23_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [8]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5000000)) 
    \niss_dsp_a1[15]_INST_0_i_12 
       (.I0(\fch/ir1 [8]),
        .I1(div_crdy1),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\niss_dsp_a1[15]_INST_0_i_24_n_0 ),
        .I5(\niss_dsp_a1[15]_INST_0_i_25_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000001AB)) 
    \niss_dsp_a1[15]_INST_0_i_13 
       (.I0(\fch/ir1 [10]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\niss_dsp_a1[15]_INST_0_i_26_n_0 ),
        .I3(\niss_dsp_a1[15]_INST_0_i_27_n_0 ),
        .I4(\niss_dsp_a1[15]_INST_0_i_28_n_0 ),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\niss_dsp_a1[15]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEEEEFFFFFEF)) 
    \niss_dsp_a1[15]_INST_0_i_14 
       (.I0(\rgf_selc1_wb[1]_i_38_n_0 ),
        .I1(\fch/ir1 [15]),
        .I2(\bcmd[2]_INST_0_i_5_n_0 ),
        .I3(\rgf/sreg/sr [7]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [14]),
        .O(\niss_dsp_a1[15]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0F04)) 
    \niss_dsp_a1[15]_INST_0_i_15 
       (.I0(\fch/ir1 [14]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [15]),
        .O(\niss_dsp_a1[15]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \niss_dsp_a1[15]_INST_0_i_16 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [7]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\fch/ir1 [9]),
        .I5(\niss_dsp_a1[15]_INST_0_i_29_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \niss_dsp_a1[15]_INST_0_i_17 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [7]),
        .O(\niss_dsp_a1[15]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \niss_dsp_a1[15]_INST_0_i_18 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [15]),
        .O(\niss_dsp_a1[15]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \niss_dsp_a1[15]_INST_0_i_19 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [10]),
        .O(\niss_dsp_a1[15]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8AAA888A8AAA8AA)) 
    \niss_dsp_a1[15]_INST_0_i_2 
       (.I0(\niss_dsp_a1[15]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a1[15]_INST_0_i_5_n_0 ),
        .I2(\niss_dsp_a1[15]_INST_0_i_6_n_0 ),
        .I3(\niss_dsp_a1[15]_INST_0_i_7_n_0 ),
        .I4(\niss_dsp_a1[15]_INST_0_i_8_n_0 ),
        .I5(\niss_dsp_a1[15]_INST_0_i_9_n_0 ),
        .O(acmd1[0]));
  LUT3 #(
    .INIT(8'h78)) 
    \niss_dsp_a1[15]_INST_0_i_20 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir1 [12]),
        .I2(\rgf/sreg/sr [5]),
        .O(\niss_dsp_a1[15]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h00000633)) 
    \niss_dsp_a1[15]_INST_0_i_21 
       (.I0(\rgf/sreg/sr [4]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [14]),
        .O(\niss_dsp_a1[15]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \niss_dsp_a1[15]_INST_0_i_22 
       (.I0(\bcmd[1]_INST_0_i_13_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [8]),
        .O(\niss_dsp_a1[15]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \niss_dsp_a1[15]_INST_0_i_23 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .O(\niss_dsp_a1[15]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[15]_INST_0_i_24 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .O(\niss_dsp_a1[15]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \niss_dsp_a1[15]_INST_0_i_25 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [9]),
        .O(\niss_dsp_a1[15]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEF00EFFFEF)) 
    \niss_dsp_a1[15]_INST_0_i_26 
       (.I0(\fch/ir1 [6]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(div_crdy1),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [9]),
        .O(\niss_dsp_a1[15]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FDDF7775)) 
    \niss_dsp_a1[15]_INST_0_i_27 
       (.I0(\bdatw[31]_INST_0_i_107_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(\niss_dsp_a1[15]_INST_0_i_30_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h80C0C0408000C080)) 
    \niss_dsp_a1[15]_INST_0_i_28 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [6]),
        .O(\niss_dsp_a1[15]_INST_0_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[15]_INST_0_i_29 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [3]),
        .O(\niss_dsp_a1[15]_INST_0_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[15]_INST_0_i_3 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0A0A0A0A88828082)) 
    \niss_dsp_a1[15]_INST_0_i_30 
       (.I0(\niss_dsp_a1[15]_INST_0_i_31_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(div_crdy1),
        .I5(\ctl1/stat_reg_n_0_[1] ),
        .O(\niss_dsp_a1[15]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[15]_INST_0_i_31 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [8]),
        .O(\niss_dsp_a1[15]_INST_0_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[15]_INST_0_i_4 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\niss_dsp_a1[32]_INST_0_i_9_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFF4)) 
    \niss_dsp_a1[15]_INST_0_i_5 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\niss_dsp_a1[15]_INST_0_i_10_n_0 ),
        .I2(\niss_dsp_a1[15]_INST_0_i_11_n_0 ),
        .I3(\niss_dsp_a1[15]_INST_0_i_12_n_0 ),
        .I4(\niss_dsp_a1[15]_INST_0_i_13_n_0 ),
        .I5(\niss_dsp_a1[15]_INST_0_i_14_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \niss_dsp_a1[15]_INST_0_i_6 
       (.I0(\fch/ir1 [11]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\rgf/sreg/sr [6]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [14]),
        .O(\niss_dsp_a1[15]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hA88AAAAA)) 
    \niss_dsp_a1[15]_INST_0_i_7 
       (.I0(\fch/ir1 [13]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [15]),
        .I4(\niss_dsp_a1[15]_INST_0_i_15_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EAAA0000)) 
    \niss_dsp_a1[15]_INST_0_i_8 
       (.I0(\niss_dsp_a1[15]_INST_0_i_16_n_0 ),
        .I1(\niss_dsp_a1[15]_INST_0_i_17_n_0 ),
        .I2(\bdatw[8]_INST_0_i_10_n_0 ),
        .I3(\bcmd[2]_INST_0_i_5_n_0 ),
        .I4(\niss_dsp_a1[15]_INST_0_i_18_n_0 ),
        .I5(\niss_dsp_a1[15]_INST_0_i_19_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF9A00FFFF)) 
    \niss_dsp_a1[15]_INST_0_i_9 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [15]),
        .I2(\niss_dsp_a1[15]_INST_0_i_20_n_0 ),
        .I3(\fch/ir1 [14]),
        .I4(\bcmd[2]_INST_0_i_5_n_0 ),
        .I5(\niss_dsp_a1[15]_INST_0_i_21_n_0 ),
        .O(\niss_dsp_a1[15]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[16]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [16]),
        .O(niss_dsp_a1[16]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[17]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [17]),
        .O(niss_dsp_a1[17]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[18]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [18]),
        .O(niss_dsp_a1[18]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[19]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [19]),
        .O(niss_dsp_a1[19]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[1]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[1]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [1]),
        .O(niss_dsp_a1[1]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[20]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [20]),
        .O(niss_dsp_a1[20]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[21]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [21]),
        .O(niss_dsp_a1[21]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[22]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [22]),
        .O(niss_dsp_a1[22]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[23]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [23]),
        .O(niss_dsp_a1[23]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[24]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [24]),
        .O(niss_dsp_a1[24]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[25]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [25]),
        .O(niss_dsp_a1[25]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[26]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [26]),
        .O(niss_dsp_a1[26]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[27]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [27]),
        .O(niss_dsp_a1[27]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[28]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [28]),
        .O(niss_dsp_a1[28]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[29]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [29]),
        .O(niss_dsp_a1[29]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[2]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[2]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [2]),
        .O(niss_dsp_a1[2]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[30]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [30]),
        .O(niss_dsp_a1[30]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[31]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [31]),
        .O(niss_dsp_a1[31]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niss_dsp_a1[32]_INST_0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [32]),
        .O(niss_dsp_a1[32]));
  LUT3 #(
    .INIT(8'h80)) 
    \niss_dsp_a1[32]_INST_0_i_1 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00A0707000000000)) 
    \niss_dsp_a1[32]_INST_0_i_10 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [13]),
        .I5(\rgf_selc1_wb[0]_i_6_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \niss_dsp_a1[32]_INST_0_i_11 
       (.I0(\niss_dsp_a1[32]_INST_0_i_24_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\rgf_selc1_wb[1]_i_5_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_25_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_26_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_11_n_0 ));
  MUXF7 \niss_dsp_a1[32]_INST_0_i_12 
       (.I0(\niss_dsp_a1[32]_INST_0_i_27_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_28_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_12_n_0 ),
        .S(\fch/ir1 [8]));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[32]_INST_0_i_13 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .O(\niss_dsp_a1[32]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFFFFFBFFFBFFF)) 
    \niss_dsp_a1[32]_INST_0_i_14 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [10]),
        .I5(\ctl1/stat_reg_n_0_[1] ),
        .O(\niss_dsp_a1[32]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8A00000088000000)) 
    \niss_dsp_a1[32]_INST_0_i_15 
       (.I0(\niss_dsp_a1[32]_INST_0_i_29_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [11]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h28282828282A2A2A)) 
    \niss_dsp_a1[32]_INST_0_i_16 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [10]),
        .O(\niss_dsp_a1[32]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0002020000020000)) 
    \niss_dsp_a1[32]_INST_0_i_17 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [11]),
        .O(\niss_dsp_a1[32]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000000002000A822)) 
    \niss_dsp_a1[32]_INST_0_i_18 
       (.I0(\niss_dsp_a1[32]_INST_0_i_30_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(div_crdy1),
        .I3(\niss_dsp_a1[32]_INST_0_i_31_n_0 ),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\niss_dsp_a1[32]_INST_0_i_32_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hA7FF5FFFFFFF5FFF)) 
    \niss_dsp_a1[32]_INST_0_i_19 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [15]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \niss_dsp_a1[32]_INST_0_i_2 
       (.I0(\rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ),
        .I1(\rgf/a1bus_b13 [15]),
        .I2(\rgf/a1bus_sr [15]),
        .I3(\rgf/a1bus_b02 [15]),
        .I4(\rgf/a1bus_out/badr[15]_INST_0_i_3_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\niss_dsp_a1[32]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4044)) 
    \niss_dsp_a1[32]_INST_0_i_20 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .I2(\niss_dsp_a1[32]_INST_0_i_33_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_34_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_35_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\niss_dsp_a1[32]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FFDF)) 
    \niss_dsp_a1[32]_INST_0_i_21 
       (.I0(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [9]),
        .I3(\niss_dsp_a1[32]_INST_0_i_36_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_37_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_38_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFF777F77F7FFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_22 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [14]),
        .O(\niss_dsp_a1[32]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000200200)) 
    \niss_dsp_a1[32]_INST_0_i_23 
       (.I0(\niss_dsp_a1[15]_INST_0_i_18_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_39_n_0 ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\niss_dsp_a1[32]_INST_0_i_40_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \niss_dsp_a1[32]_INST_0_i_24 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [15]),
        .O(\niss_dsp_a1[32]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hEFFF)) 
    \niss_dsp_a1[32]_INST_0_i_25 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [0]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .O(\niss_dsp_a1[32]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \niss_dsp_a1[32]_INST_0_i_26 
       (.I0(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [9]),
        .O(\niss_dsp_a1[32]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAAAA2A)) 
    \niss_dsp_a1[32]_INST_0_i_27 
       (.I0(\niss_dsp_a1[32]_INST_0_i_41_n_0 ),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_42_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [7]),
        .I5(\niss_dsp_a1[32]_INST_0_i_43_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDDD0DDDD)) 
    \niss_dsp_a1[32]_INST_0_i_28 
       (.I0(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_44_n_0 ),
        .I2(\bcmd[1]_INST_0_i_13_n_0 ),
        .I3(\fch/ir1 [9]),
        .I4(div_crdy1),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h111111111F111111)) 
    \niss_dsp_a1[32]_INST_0_i_29 
       (.I0(\niss_dsp_a1[32]_INST_0_i_45_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\niss_dsp_a1[32]_INST_0_i_46_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [8]),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\niss_dsp_a1[32]_INST_0_i_29_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_3 
       (.I0(acmd1[4]),
        .I1(acmd1[3]),
        .O(\niss_dsp_a1[32]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0504)) 
    \niss_dsp_a1[32]_INST_0_i_30 
       (.I0(\fch/ir1 [9]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(div_crdy1),
        .O(\niss_dsp_a1[32]_INST_0_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_31 
       (.I0(\fch/ir1 [7]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .O(\niss_dsp_a1[32]_INST_0_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \niss_dsp_a1[32]_INST_0_i_32 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [10]),
        .O(\niss_dsp_a1[32]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00000E0000000000)) 
    \niss_dsp_a1[32]_INST_0_i_33 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\fch/ir1 [6]),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\fch/ir1 [8]),
        .O(\niss_dsp_a1[32]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF07FFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_34 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [10]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(\fch/ir1 [8]),
        .O(\niss_dsp_a1[32]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \niss_dsp_a1[32]_INST_0_i_35 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [8]),
        .I4(div_crdy1),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\niss_dsp_a1[32]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hF7CEFFBFFFDFDFEF)) 
    \niss_dsp_a1[32]_INST_0_i_36 
       (.I0(\fch/ir1 [4]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [3]),
        .O(\niss_dsp_a1[32]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h00000020FFFFFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_37 
       (.I0(\bcmd[1]_INST_0_i_26_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [6]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [11]),
        .O(\niss_dsp_a1[32]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h6200000022003300)) 
    \niss_dsp_a1[32]_INST_0_i_38 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(div_crdy1),
        .I3(\rgf_selc1_rn_wb[1]_i_24_n_0 ),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [10]),
        .O(\niss_dsp_a1[32]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \niss_dsp_a1[32]_INST_0_i_39 
       (.I0(\bcmd[0]_INST_0_i_12_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [1]),
        .O(\niss_dsp_a1[32]_INST_0_i_39_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[32]_INST_0_i_4 
       (.I0(acmd1[0]),
        .I1(dctl_sign_f_i_2_n_0),
        .O(\niss_dsp_a1[32]_INST_0_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \niss_dsp_a1[32]_INST_0_i_40 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [7]),
        .O(\niss_dsp_a1[32]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h5F5F7FFF55D57FFF)) 
    \niss_dsp_a1[32]_INST_0_i_41 
       (.I0(\niss_dsp_a1[32]_INST_0_i_47_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [9]),
        .O(\niss_dsp_a1[32]_INST_0_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_a1[32]_INST_0_i_42 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [9]),
        .O(\niss_dsp_a1[32]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h2220000002000000)) 
    \niss_dsp_a1[32]_INST_0_i_43 
       (.I0(\niss_dsp_a1[32]_INST_0_i_30_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [10]),
        .I5(div_crdy1),
        .O(\niss_dsp_a1[32]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFF03AAAAFFFFAAAA)) 
    \niss_dsp_a1[32]_INST_0_i_44 
       (.I0(\niss_dsp_a1[32]_INST_0_i_48_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(div_crdy1),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\fch/ir1 [7]),
        .I5(\niss_dsp_a1[32]_INST_0_i_49_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF704)) 
    \niss_dsp_a1[32]_INST_0_i_45 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [7]),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .O(\niss_dsp_a1[32]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF7FFFFFF)) 
    \niss_dsp_a1[32]_INST_0_i_46 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [9]),
        .I5(\ctl1/stat_reg_n_0_[1] ),
        .O(\niss_dsp_a1[32]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_a1[32]_INST_0_i_47 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [10]),
        .O(\niss_dsp_a1[32]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAAAAAAAFDFD)) 
    \niss_dsp_a1[32]_INST_0_i_48 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\fch/ir1 [6]),
        .O(\niss_dsp_a1[32]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'h5D557FF5)) 
    \niss_dsp_a1[32]_INST_0_i_49 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [6]),
        .O(\niss_dsp_a1[32]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h5454545454555454)) 
    \niss_dsp_a1[32]_INST_0_i_5 
       (.I0(\niss_dsp_a1[32]_INST_0_i_9_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_10_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_11_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_12_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_13_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_14_n_0 ),
        .O(\niss_dsp_a1[32]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \niss_dsp_a1[32]_INST_0_i_6 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf/sreg/sr [15]),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_14_n_0 ),
        .O(\rgf/a1bus_sr [15]));
  LUT6 #(
    .INIT(64'h00000000FFFE0000)) 
    \niss_dsp_a1[32]_INST_0_i_7 
       (.I0(\niss_dsp_a1[32]_INST_0_i_15_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_16_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_17_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_18_n_0 ),
        .I4(\niss_dsp_a1[15]_INST_0_i_4_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_19_n_0 ),
        .O(acmd1[4]));
  LUT6 #(
    .INIT(64'hAAAAAAAA0008AAAA)) 
    \niss_dsp_a1[32]_INST_0_i_8 
       (.I0(\niss_dsp_a1[15]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_20_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_21_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_14_n_0 ),
        .I4(\niss_dsp_a1[32]_INST_0_i_22_n_0 ),
        .I5(\niss_dsp_a1[32]_INST_0_i_23_n_0 ),
        .O(acmd1[3]));
  LUT5 #(
    .INIT(32'h00000008)) 
    \niss_dsp_a1[32]_INST_0_i_9 
       (.I0(\niss_dsp_a1[32]_INST_0_i_16_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [11]),
        .O(\niss_dsp_a1[32]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[3]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[3]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [3]),
        .O(niss_dsp_a1[3]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[4]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[4]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [4]),
        .O(niss_dsp_a1[4]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[5]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[5]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [5]),
        .O(niss_dsp_a1[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[6]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[6]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [6]),
        .O(niss_dsp_a1[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[7]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[7]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [7]),
        .O(niss_dsp_a1[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[8]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [8]),
        .O(niss_dsp_a1[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_a1[9]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[9]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_a [9]),
        .O(niss_dsp_a1[9]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[0]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[0] ),
        .O(niss_dsp_b0[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[10]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[10]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[10] ),
        .O(niss_dsp_b0[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[11]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[11]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[11] ),
        .O(niss_dsp_b0[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[12]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[12]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[12] ),
        .O(niss_dsp_b0[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[13]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[13]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[13] ),
        .O(niss_dsp_b0[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[14]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[14]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[14] ),
        .O(niss_dsp_b0[14]));
  LUT5 #(
    .INIT(32'hC000E222)) 
    \niss_dsp_b0[15]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/mul/mul_rslt ),
        .I3(\alu0/mul/mul_b_reg_n_0_[15] ),
        .I4(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .O(niss_dsp_b0[15]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[16]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[16] ),
        .O(niss_dsp_b0[16]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[17]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[17] ),
        .O(niss_dsp_b0[17]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[18]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[18] ),
        .O(niss_dsp_b0[18]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[19]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[19] ),
        .O(niss_dsp_b0[19]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[1]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[1] ),
        .O(niss_dsp_b0[1]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[20]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[20] ),
        .O(niss_dsp_b0[20]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[21]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[21] ),
        .O(niss_dsp_b0[21]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[22]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[22] ),
        .O(niss_dsp_b0[22]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[23]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[23] ),
        .O(niss_dsp_b0[23]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[24]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[24] ),
        .O(niss_dsp_b0[24]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[25]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[25] ),
        .O(niss_dsp_b0[25]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[26]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[26] ),
        .O(niss_dsp_b0[26]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[27]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[27] ),
        .O(niss_dsp_b0[27]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[28]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[28] ),
        .O(niss_dsp_b0[28]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[29]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[29] ),
        .O(niss_dsp_b0[29]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[2]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[2] ),
        .O(niss_dsp_b0[2]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[30]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[30] ),
        .O(niss_dsp_b0[30]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[31]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[31] ),
        .O(niss_dsp_b0[31]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b0[32]_INST_0 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a0[32]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[32] ),
        .O(niss_dsp_b0[32]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[3]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[3] ),
        .O(niss_dsp_b0[3]));
  LUT5 #(
    .INIT(32'h808080FF)) 
    \niss_dsp_b0[4]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu0/mul/mul_rslt ),
        .I2(\alu0/mul/mul_b_reg_n_0_[4] ),
        .I3(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .O(niss_dsp_b0[4]));
  LUT2 #(
    .INIT(4'hE)) 
    \niss_dsp_b0[4]_INST_0_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\niss_dsp_b0[4]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[5]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[5] ),
        .O(niss_dsp_b0[5]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b0[6]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[6] ),
        .O(niss_dsp_b0[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[7]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[7]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[7] ),
        .O(niss_dsp_b0[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[8]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[8]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[8] ),
        .O(niss_dsp_b0[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b0[9]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(b0bus_0[9]),
        .I3(\alu0/mul/mul_rslt ),
        .I4(\alu0/mul/mul_b_reg_n_0_[9] ),
        .O(niss_dsp_b0[9]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[0]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[0] ),
        .O(niss_dsp_b1[0]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \niss_dsp_b1[0]_INST_0_i_1 
       (.I0(\niss_dsp_b1[0]_INST_0_i_2_n_0 ),
        .I1(\rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_5_n_0 ),
        .I4(\rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_6_n_0 ),
        .I5(p_2_in4_in[0]),
        .O(\niss_dsp_b1[0]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \niss_dsp_b1[0]_INST_0_i_12 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \niss_dsp_b1[0]_INST_0_i_13 
       (.I0(\rgf/b1bus_sel_0 [6]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/bank02/gr26 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFDFF5F5F5755FFFF)) 
    \niss_dsp_b1[0]_INST_0_i_2 
       (.I0(ctl_selb1_0[2]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [0]),
        .I3(\niss_dsp_b1[0]_INST_0_i_8_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(\niss_dsp_b1[0]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \niss_dsp_b1[0]_INST_0_i_22 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sr [0]));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_23 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr03 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_24 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_25 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr07 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_26 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_27 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr23 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_28 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr21 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_29 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr27 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[0]_INST_0_i_30 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [0]),
        .O(\niss_dsp_b1[0]_INST_0_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \niss_dsp_b1[0]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [0]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[0]));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_b1[0]_INST_0_i_8 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [3]),
        .O(\niss_dsp_b1[0]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[10]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[10]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[10] ),
        .O(niss_dsp_b1[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[11]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[11]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[11] ),
        .O(niss_dsp_b1[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[12]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[12]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[12] ),
        .O(niss_dsp_b1[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[13]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[13]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[13] ),
        .O(niss_dsp_b1[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[14]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[14]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[14] ),
        .O(niss_dsp_b1[14]));
  LUT5 #(
    .INIT(32'hC000E222)) 
    \niss_dsp_b1[15]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/mul/mul_rslt ),
        .I3(\alu1/mul/mul_b_reg_n_0_[15] ),
        .I4(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .O(niss_dsp_b1[15]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[16]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[16] ),
        .O(niss_dsp_b1[16]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[17]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[17] ),
        .O(niss_dsp_b1[17]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[18]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[18] ),
        .O(niss_dsp_b1[18]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[19]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[19] ),
        .O(niss_dsp_b1[19]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[1]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[1] ),
        .O(niss_dsp_b1[1]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \niss_dsp_b1[1]_INST_0_i_1 
       (.I0(\niss_dsp_b1[1]_INST_0_i_2_n_0 ),
        .I1(\rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_5_n_0 ),
        .I4(\rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_6_n_0 ),
        .I5(p_2_in4_in[1]),
        .O(\niss_dsp_b1[1]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \niss_dsp_b1[1]_INST_0_i_12 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \niss_dsp_b1[1]_INST_0_i_13 
       (.I0(\rgf/b1bus_sel_0 [6]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/bank02/gr26 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \niss_dsp_b1[1]_INST_0_i_2 
       (.I0(\fch/ir1 [0]),
        .I1(ctl_selb1_0[1]),
        .I2(\niss_dsp_b1[1]_INST_0_i_8_n_0 ),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(\fch/ir1 [1]),
        .I5(ctl_selb1_0[2]),
        .O(\niss_dsp_b1[1]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \niss_dsp_b1[1]_INST_0_i_22 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sr [1]));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_23 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr03 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_24 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_25 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr07 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_26 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_27 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr23 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_28 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr21 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_29 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr27 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[1]_INST_0_i_30 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\niss_dsp_b1[1]_INST_0_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \niss_dsp_b1[1]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [1]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[1]));
  LUT4 #(
    .INIT(16'h0004)) 
    \niss_dsp_b1[1]_INST_0_i_8 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [2]),
        .O(\niss_dsp_b1[1]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[20]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[20] ),
        .O(niss_dsp_b1[20]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[21]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[21] ),
        .O(niss_dsp_b1[21]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[22]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[22] ),
        .O(niss_dsp_b1[22]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[23]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[23] ),
        .O(niss_dsp_b1[23]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[24]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[24] ),
        .O(niss_dsp_b1[24]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[25]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[25] ),
        .O(niss_dsp_b1[25]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[26]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[26] ),
        .O(niss_dsp_b1[26]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[27]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[27] ),
        .O(niss_dsp_b1[27]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[28]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[28] ),
        .O(niss_dsp_b1[28]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[29]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[29] ),
        .O(niss_dsp_b1[29]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[2]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[2] ),
        .O(niss_dsp_b1[2]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \niss_dsp_b1[2]_INST_0_i_1 
       (.I0(\niss_dsp_b1[2]_INST_0_i_2_n_0 ),
        .I1(\rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_3_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_4_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_5_n_0 ),
        .I4(\rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_6_n_0 ),
        .I5(p_2_in4_in[2]),
        .O(\niss_dsp_b1[2]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \niss_dsp_b1[2]_INST_0_i_13 
       (.I0(\bank02/b1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00080000)) 
    \niss_dsp_b1[2]_INST_0_i_14 
       (.I0(\rgf/b1bus_sel_0 [6]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/bank02/gr26 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0CD13FD1FFFFFFFF)) 
    \niss_dsp_b1[2]_INST_0_i_2 
       (.I0(\fch/ir1 [1]),
        .I1(ctl_selb1_0[1]),
        .I2(\niss_dsp_b1[2]_INST_0_i_8_n_0 ),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(\fch/ir1 [2]),
        .I5(ctl_selb1_0[2]),
        .O(\niss_dsp_b1[2]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \niss_dsp_b1[2]_INST_0_i_24 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\rgf/sreg/sr [2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sr [2]));
  LUT6 #(
    .INIT(64'h5151FF51FFFFFFFF)) 
    \niss_dsp_b1[2]_INST_0_i_27 
       (.I0(\niss_dsp_b1[2]_INST_0_i_36_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_53_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_56_n_0 ),
        .I3(\niss_dsp_b1[2]_INST_0_i_37_n_0 ),
        .I4(\niss_dsp_b1[2]_INST_0_i_38_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_49_n_0 ),
        .O(\niss_dsp_b1[2]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_28 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr03 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_29 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_30 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr07 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_31 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_32 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr23 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_33 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr21 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_34 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr27 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[2]_INST_0_i_35 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h5555400040004000)) 
    \niss_dsp_b1[2]_INST_0_i_36 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I2(\niss_dsp_b1[2]_INST_0_i_39_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_31_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_74_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_73_n_0 ),
        .O(\niss_dsp_b1[2]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h555555557F777F7F)) 
    \niss_dsp_b1[2]_INST_0_i_37 
       (.I0(\rgf_selc1_rn_wb[0]_i_4_n_0 ),
        .I1(ctl_fetch1_fl_i_16_n_0),
        .I2(\niss_dsp_b1[5]_INST_0_i_69_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_68_n_0 ),
        .I4(\fch/ir1 [0]),
        .I5(\badr[31]_INST_0_i_101_n_0 ),
        .O(\niss_dsp_b1[2]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \niss_dsp_b1[2]_INST_0_i_38 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [0]),
        .I3(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .O(\niss_dsp_b1[2]_INST_0_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \niss_dsp_b1[2]_INST_0_i_39 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [2]),
        .O(\niss_dsp_b1[2]_INST_0_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \niss_dsp_b1[2]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [2]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[2]));
  LUT4 #(
    .INIT(16'h0100)) 
    \niss_dsp_b1[2]_INST_0_i_8 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [1]),
        .O(\niss_dsp_b1[2]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[30]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[30] ),
        .O(niss_dsp_b1[30]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[31]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[31] ),
        .O(niss_dsp_b1[31]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niss_dsp_b1[32]_INST_0 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\niss_dsp_a1[32]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[32] ),
        .O(niss_dsp_b1[32]));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[3]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[3] ),
        .O(niss_dsp_b1[3]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \niss_dsp_b1[3]_INST_0_i_1 
       (.I0(\niss_dsp_b1[3]_INST_0_i_2_n_0 ),
        .I1(\niss_dsp_b1[3]_INST_0_i_3_n_0 ),
        .I2(p_2_in4_in[3]),
        .I3(\rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_5_n_0 ),
        .I4(\rgf/b1bus_b02 [3]),
        .I5(\rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_7_n_0 ),
        .O(\niss_dsp_b1[3]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \niss_dsp_b1[3]_INST_0_i_13 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\rgf/sreg/sr [3]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sr [3]));
  LUT6 #(
    .INIT(64'hAAAABBBBAAAAFBBB)) 
    \niss_dsp_b1[3]_INST_0_i_2 
       (.I0(\niss_dsp_b1[5]_INST_0_i_8_n_0 ),
        .I1(ctl_selb1_0[1]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_20 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr03 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_21 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_22 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr07 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_23 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_24 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr23 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_25 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr21 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_26 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr27 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_27 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_28 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr07 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_29 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h2222222200008000)) 
    \niss_dsp_b1[3]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(ctl_selb1_0[1]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_30 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr27 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[3]_INST_0_i_31 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr25 [3]),
        .O(\niss_dsp_b1[3]_INST_0_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \niss_dsp_b1[3]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [3]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[3]));
  LUT5 #(
    .INIT(32'h808080FF)) 
    \niss_dsp_b1[4]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu1/mul/mul_rslt ),
        .I2(\alu1/mul/mul_b_reg_n_0_[4] ),
        .I3(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .O(niss_dsp_b1[4]));
  LUT2 #(
    .INIT(4'hE)) 
    \niss_dsp_b1[4]_INST_0_i_1 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\niss_dsp_b1[4]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[5]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[5] ),
        .O(niss_dsp_b1[5]));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \niss_dsp_b1[5]_INST_0_i_1 
       (.I0(\niss_dsp_b1[5]_INST_0_i_2_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_3_n_0 ),
        .I2(p_2_in4_in[5]),
        .I3(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_5_n_0 ),
        .I4(\rgf/b1bus_b02 [5]),
        .I5(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_7_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \niss_dsp_b1[5]_INST_0_i_15 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_rn[0]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .I4(ctl_selb1_rn[1]),
        .O(\rgf/b1bus_sr [5]));
  LUT6 #(
    .INIT(64'hABABABFBABABABAB)) 
    \niss_dsp_b1[5]_INST_0_i_2 
       (.I0(\niss_dsp_b1[5]_INST_0_i_8_n_0 ),
        .I1(\fch/ir1 [4]),
        .I2(ctl_selb1_0[1]),
        .I3(\niss_dsp_b1[5]_INST_0_i_9_n_0 ),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [0]),
        .O(\niss_dsp_b1[5]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF40FF40404040)) 
    \niss_dsp_b1[5]_INST_0_i_22 
       (.I0(\niss_dsp_b1[5]_INST_0_i_48_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_49_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_51_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_52_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_53_n_0 ),
        .O(ctl_selb1_rn[1]));
  LUT6 #(
    .INIT(64'h808080AA80808080)) 
    \niss_dsp_b1[5]_INST_0_i_23 
       (.I0(\niss_dsp_b1[5]_INST_0_i_49_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_54_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [15]),
        .I5(\niss_dsp_b1[5]_INST_0_i_55_n_0 ),
        .O(ctl_selb1_rn[0]));
  LUT6 #(
    .INIT(64'h040004000400FFFF)) 
    \niss_dsp_b1[5]_INST_0_i_24 
       (.I0(\niss_dsp_b1[5]_INST_0_i_56_n_0 ),
        .I1(\bcmd[0]_INST_0_i_4_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(ctl_fetch1_fl_i_16_n_0),
        .I4(\niss_dsp_b1[5]_INST_0_i_57_n_0 ),
        .I5(\ctl1/stat_reg_n_0_[2] ),
        .O(ctl_selb1_rn[2]));
  LUT3 #(
    .INIT(8'hBF)) 
    \niss_dsp_b1[5]_INST_0_i_25 
       (.I0(ctl_selb1_0[2]),
        .I1(\bdatw[31]_INST_0_i_12_n_0 ),
        .I2(ctl_selb1_0[1]),
        .O(\niss_dsp_b1[5]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_26 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr03 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_28 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr01 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h080808080808A808)) 
    \niss_dsp_b1[5]_INST_0_i_3 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(ctl_selb1_0[1]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [1]),
        .I5(\niss_dsp_b1[5]_INST_0_i_9_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_30 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr07 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_31 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_33 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr23 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_35 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr21 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_37 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr27 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_38 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_38_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \niss_dsp_b1[5]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_11_n_0 ),
        .I1(\fch/eir [5]),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(p_2_in4_in[5]));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_40 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr07 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_42 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_45 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr27 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_46 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr25 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \niss_dsp_b1[5]_INST_0_i_48 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [6]),
        .O(\niss_dsp_b1[5]_INST_0_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niss_dsp_b1[5]_INST_0_i_49 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .O(\niss_dsp_b1[5]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000600000)) 
    \niss_dsp_b1[5]_INST_0_i_50 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [8]),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hD0D5D5DDFFFFFFFF)) 
    \niss_dsp_b1[5]_INST_0_i_51 
       (.I0(\fch/ir1 [1]),
        .I1(\niss_dsp_b1[5]_INST_0_i_63_n_0 ),
        .I2(\stat[1]_i_22_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(\badr[31]_INST_0_i_102_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAA200AAAAAAAA)) 
    \niss_dsp_b1[5]_INST_0_i_52 
       (.I0(\sr[15]_i_6_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_64_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_65_n_0 ),
        .I3(\fch/ir1 [1]),
        .I4(\niss_dsp_b1[5]_INST_0_i_66_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_67_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_53 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [14]),
        .O(\niss_dsp_b1[5]_INST_0_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \niss_dsp_b1[5]_INST_0_i_54 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .O(\niss_dsp_b1[5]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFAEAAAAAAAAAAAA)) 
    \niss_dsp_b1[5]_INST_0_i_55 
       (.I0(\badr[31]_INST_0_i_101_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\niss_dsp_b1[5]_INST_0_i_68_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_69_n_0 ),
        .I4(\fch/ir1 [13]),
        .I5(\fch/ir1 [14]),
        .O(\niss_dsp_b1[5]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h000000D5DDDDDDDD)) 
    \niss_dsp_b1[5]_INST_0_i_56 
       (.I0(\fch/ir1 [2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_68_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_70_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_71_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_72_n_0 ),
        .I5(\sr[15]_i_6_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h0777777777777777)) 
    \niss_dsp_b1[5]_INST_0_i_57 
       (.I0(\niss_dsp_b1[5]_INST_0_i_73_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_74_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_31_n_0 ),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [6]),
        .I5(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFF54FFFFFF54FF54)) 
    \niss_dsp_b1[5]_INST_0_i_58 
       (.I0(\niss_dsp_b1[5]_INST_0_i_75_n_0 ),
        .I1(\bdatw[31]_INST_0_i_43_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_76_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_77_n_0 ),
        .I4(\bdatw[31]_INST_0_i_102_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_78_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFF0FFFBFBF0FF)) 
    \niss_dsp_b1[5]_INST_0_i_59 
       (.I0(\niss_dsp_b1[5]_INST_0_i_52_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_51_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_79_n_0 ),
        .I3(\niss_dsp_b1[2]_INST_0_i_36_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_53_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_56_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hBBFAFBFAFFFFFFFF)) 
    \niss_dsp_b1[5]_INST_0_i_60 
       (.I0(\bdatw[15]_INST_0_i_90_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_48_n_0 ),
        .I2(\niss_dsp_b1[2]_INST_0_i_37_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_54_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_49_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hDF5F0F0FDD5F0F0F)) 
    \niss_dsp_b1[5]_INST_0_i_61 
       (.I0(\niss_dsp_b1[2]_INST_0_i_37_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_54_n_0 ),
        .I2(\bdatw[15]_INST_0_i_90_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_49_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_48_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h454545454FFF4F4F)) 
    \niss_dsp_b1[5]_INST_0_i_62 
       (.I0(\niss_dsp_b1[2]_INST_0_i_36_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_56_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_53_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_52_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_51_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_79_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAA888AAAA)) 
    \niss_dsp_b1[5]_INST_0_i_63 
       (.I0(\badr[31]_INST_0_i_167_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(div_crdy1),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_63_n_0 ));
  LUT5 #(
    .INIT(32'hCDFDCECC)) 
    \niss_dsp_b1[5]_INST_0_i_64 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [8]),
        .O(\niss_dsp_b1[5]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'h00F70000)) 
    \niss_dsp_b1[5]_INST_0_i_65 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(div_crdy1),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .O(\niss_dsp_b1[5]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEAAAAAAA)) 
    \niss_dsp_b1[5]_INST_0_i_66 
       (.I0(\niss_dsp_b1[5]_INST_0_i_80_n_0 ),
        .I1(\bdatw[31]_INST_0_i_113_n_0 ),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [6]),
        .I4(\bdatw[31]_INST_0_i_139_n_0 ),
        .I5(\fch/ir1 [3]),
        .O(\niss_dsp_b1[5]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hB7FF47FFFFFFFFFF)) 
    \niss_dsp_b1[5]_INST_0_i_67 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [3]),
        .I5(\stat[2]_i_13_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'hFFFB0000FFFFFFFF)) 
    \niss_dsp_b1[5]_INST_0_i_68 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(div_crdy1),
        .I2(\bdatw[31]_INST_0_i_151_n_0 ),
        .I3(\fch/ir1 [8]),
        .I4(\niss_dsp_b1[5]_INST_0_i_81_n_0 ),
        .I5(\badr[31]_INST_0_i_102_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h080808080808AA08)) 
    \niss_dsp_b1[5]_INST_0_i_69 
       (.I0(\sr[15]_i_6_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\niss_dsp_b1[5]_INST_0_i_82_n_0 ),
        .I3(\fch/ir1 [8]),
        .I4(\stat[1]_i_22_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_83_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hAA82AAAAAAAAAAAA)) 
    \niss_dsp_b1[5]_INST_0_i_70 
       (.I0(\niss_dsp_b1[5]_INST_0_i_64_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [6]),
        .I5(\bdatw[31]_INST_0_i_113_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h0888008080000080)) 
    \niss_dsp_b1[5]_INST_0_i_71 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h4000444444044444)) 
    \niss_dsp_b1[5]_INST_0_i_72 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [8]),
        .I3(div_crdy1),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [6]),
        .O(\niss_dsp_b1[5]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \niss_dsp_b1[5]_INST_0_i_73 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [15]),
        .I3(\rgf_selc1_rn_wb[1]_i_21_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \niss_dsp_b1[5]_INST_0_i_74 
       (.I0(\fch/ir1 [6]),
        .I1(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [0]),
        .I5(\fch/ir1 [1]),
        .O(\niss_dsp_b1[5]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'hFFAE00AE00000000)) 
    \niss_dsp_b1[5]_INST_0_i_75 
       (.I0(\stat[1]_i_12__0_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_84_n_0 ),
        .I2(\bdatw[31]_INST_0_i_115_n_0 ),
        .I3(\fch/ir1 [12]),
        .I4(\bdatw[31]_INST_0_i_114_n_0 ),
        .I5(\bdatw[31]_INST_0_i_44_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000005575)) 
    \niss_dsp_b1[5]_INST_0_i_76 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\bdatw[31]_INST_0_i_105_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_85_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_86_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_87_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_88_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'hBFBFBFBABFBFBFBF)) 
    \niss_dsp_b1[5]_INST_0_i_77 
       (.I0(\bcmd[3]_INST_0_i_4_n_0 ),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [2]),
        .I4(\niss_dsp_b1[5]_INST_0_i_89_n_0 ),
        .I5(\bcmd[1]_INST_0_i_24_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAEF)) 
    \niss_dsp_b1[5]_INST_0_i_78 
       (.I0(\bdatw[31]_INST_0_i_100_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_90_n_0 ),
        .I2(\bdatw[31]_INST_0_i_146_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_91_n_0 ),
        .I4(\bdatw[31]_INST_0_i_144_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_92_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \niss_dsp_b1[5]_INST_0_i_79 
       (.I0(\niss_dsp_b1[5]_INST_0_i_50_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [6]),
        .O(\niss_dsp_b1[5]_INST_0_i_79_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \niss_dsp_b1[5]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_12_n_0 ),
        .I1(ctl_selb1_0[2]),
        .O(\niss_dsp_b1[5]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \niss_dsp_b1[5]_INST_0_i_80 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [9]),
        .O(\niss_dsp_b1[5]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h3FF33F3F3F77FF33)) 
    \niss_dsp_b1[5]_INST_0_i_81 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [9]),
        .O(\niss_dsp_b1[5]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF40E022224A4A)) 
    \niss_dsp_b1[5]_INST_0_i_82 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [7]),
        .I3(div_crdy1),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [10]),
        .O(\niss_dsp_b1[5]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h9B5FFF3F7FBFDD7F)) 
    \niss_dsp_b1[5]_INST_0_i_83 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [5]),
        .O(\niss_dsp_b1[5]_INST_0_i_83_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \niss_dsp_b1[5]_INST_0_i_84 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir1 [13]),
        .O(\niss_dsp_b1[5]_INST_0_i_84_n_0 ));
  LUT4 #(
    .INIT(16'h4FFF)) 
    \niss_dsp_b1[5]_INST_0_i_85 
       (.I0(\bdatw[31]_INST_0_i_152_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_93_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [11]),
        .O(\niss_dsp_b1[5]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABAAABAAABBBB)) 
    \niss_dsp_b1[5]_INST_0_i_86 
       (.I0(\bdatw[31]_INST_0_i_110_n_0 ),
        .I1(\bdatw[31]_INST_0_i_109_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_94_n_0 ),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \niss_dsp_b1[5]_INST_0_i_87 
       (.I0(\bdatw[31]_INST_0_i_113_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_95_n_0 ),
        .I2(\bdatw[31]_INST_0_i_153_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [11]),
        .O(\niss_dsp_b1[5]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h0000000060000000)) 
    \niss_dsp_b1[5]_INST_0_i_88 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [11]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\bcmd[1]_INST_0_i_13_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_31_n_0 ),
        .I5(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \niss_dsp_b1[5]_INST_0_i_89 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [5]),
        .I3(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I4(\bdatw[31]_INST_0_i_173_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_96_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_89_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \niss_dsp_b1[5]_INST_0_i_9 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [2]),
        .O(\niss_dsp_b1[5]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hAAFB)) 
    \niss_dsp_b1[5]_INST_0_i_90 
       (.I0(\fch/ir1 [11]),
        .I1(div_crdy1),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\fch/ir1 [10]),
        .O(\niss_dsp_b1[5]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'hAA20AA20AA20AAAA)) 
    \niss_dsp_b1[5]_INST_0_i_91 
       (.I0(\fch/ir1 [11]),
        .I1(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I2(\bdatw[31]_INST_0_i_172_n_0 ),
        .I3(\bdatw[31]_INST_0_i_171_n_0 ),
        .I4(\bdatw[31]_INST_0_i_170_n_0 ),
        .I5(\bdatw[31]_INST_0_i_169_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000F202F2)) 
    \niss_dsp_b1[5]_INST_0_i_92 
       (.I0(div_crdy1),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [6]),
        .I5(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .O(\niss_dsp_b1[5]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hE6FDFFFFFFFFFFFF)) 
    \niss_dsp_b1[5]_INST_0_i_93 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [6]),
        .O(\niss_dsp_b1[5]_INST_0_i_93_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \niss_dsp_b1[5]_INST_0_i_94 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(div_crdy1),
        .O(\niss_dsp_b1[5]_INST_0_i_94_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niss_dsp_b1[5]_INST_0_i_95 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .O(\niss_dsp_b1[5]_INST_0_i_95_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \niss_dsp_b1[5]_INST_0_i_96 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [6]),
        .O(\niss_dsp_b1[5]_INST_0_i_96_n_0 ));
  LUT5 #(
    .INIT(32'hAB010101)) 
    \niss_dsp_b1[6]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[6] ),
        .O(niss_dsp_b1[6]));
  LUT6 #(
    .INIT(64'h0202020200020202)) 
    \niss_dsp_b1[6]_INST_0_i_1 
       (.I0(\niss_dsp_b1[6]_INST_0_i_2_n_0 ),
        .I1(\rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_3_n_0 ),
        .I2(\rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [6]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(\niss_dsp_b1[6]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h52A257A7FFFFFFFF)) 
    \niss_dsp_b1[6]_INST_0_i_2 
       (.I0(\bdatw[31]_INST_0_i_12_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(ctl_selb1_0[1]),
        .I3(\niss_dsp_b1[6]_INST_0_i_5_n_0 ),
        .I4(\fch/ir1 [5]),
        .I5(ctl_selb1_0[2]),
        .O(\niss_dsp_b1[6]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \niss_dsp_b1[6]_INST_0_i_5 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [3]),
        .O(\niss_dsp_b1[6]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[7]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[7]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[7] ),
        .O(niss_dsp_b1[7]));
  LUT6 #(
    .INIT(64'hFEFEFEFEFFFEFEFE)) 
    \niss_dsp_b1[7]_INST_0_i_1 
       (.I0(\niss_dsp_b1[7]_INST_0_i_2_n_0 ),
        .I1(\rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_3_n_0 ),
        .I2(\rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_4_n_0 ),
        .I3(\bdatw[31]_INST_0_i_11_n_0 ),
        .I4(\fch/eir [7]),
        .I5(\bdatw[31]_INST_0_i_12_n_0 ),
        .O(b1bus_0[7]));
  LUT6 #(
    .INIT(64'hAA0A08A8A00008A8)) 
    \niss_dsp_b1[7]_INST_0_i_2 
       (.I0(ctl_selb1_0[2]),
        .I1(\fch/ir1 [6]),
        .I2(ctl_selb1_0[1]),
        .I3(\niss_dsp_b1[7]_INST_0_i_5_n_0 ),
        .I4(\bdatw[31]_INST_0_i_12_n_0 ),
        .I5(\fch/ir1 [7]),
        .O(\niss_dsp_b1[7]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \niss_dsp_b1[7]_INST_0_i_5 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [2]),
        .I3(\fch/ir1 [3]),
        .O(\niss_dsp_b1[7]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[8]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[8]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[8] ),
        .O(niss_dsp_b1[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niss_dsp_b1[9]_INST_0 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(b1bus_0[9]),
        .I3(\alu1/mul/mul_rslt ),
        .I4(\alu1/mul/mul_b_reg_n_0_[9] ),
        .O(niss_dsp_b1[9]));
  LUT4 #(
    .INIT(16'hBA8A)) 
    \pc0[0]_i_1 
       (.I0(\rgf/pcnt/pc [0]),
        .I1(fch_irq_req),
        .I2(\pc0[15]_i_4_n_0 ),
        .I3(\fch/p_2_in0_in [0]),
        .O(fch_pc[0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[10]_i_1 
       (.I0(\pc0[10]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [10]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[10]_i_3_n_0 ),
        .O(fch_pc[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[10]_i_2 
       (.I0(\fch/p_2_in [10]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [10]),
        .O(\pc0[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[10]_i_3 
       (.I0(\fch/p_2_in [10]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[12]_INST_0_i_1_n_6 ),
        .O(\pc0[10]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[11]_i_1 
       (.I0(\pc0[11]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [11]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[11]_i_4_n_0 ),
        .O(fch_pc[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[11]_i_2 
       (.I0(\fch/p_2_in [11]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [11]),
        .O(\pc0[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[11]_i_4 
       (.I0(\fch/p_2_in [11]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[12]_INST_0_i_1_n_5 ),
        .O(\pc0[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[12]_i_1 
       (.I0(\pc0[12]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [12]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[12]_i_3_n_0 ),
        .O(fch_pc[12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[12]_i_2 
       (.I0(\fch/p_2_in [12]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [12]),
        .O(\pc0[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[12]_i_3 
       (.I0(\fch/p_2_in [12]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[12]_INST_0_i_1_n_4 ),
        .O(\pc0[12]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[13]_i_1 
       (.I0(\pc0[13]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [13]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[13]_i_3_n_0 ),
        .O(fch_pc[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[13]_i_2 
       (.I0(\fch/p_2_in [13]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [13]),
        .O(\pc0[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[13]_i_3 
       (.I0(\fch/p_2_in [13]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[15]_INST_0_i_4_n_7 ),
        .O(\pc0[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[14]_i_1 
       (.I0(\pc0[14]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [14]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[14]_i_3_n_0 ),
        .O(fch_pc[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[14]_i_2 
       (.I0(\fch/p_2_in [14]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [14]),
        .O(\pc0[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[14]_i_3 
       (.I0(\fch/p_2_in [14]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[15]_INST_0_i_4_n_6 ),
        .O(\pc0[14]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[15]_i_1 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [15]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[15]_i_5_n_0 ),
        .O(fch_pc[15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[15]_i_2 
       (.I0(\fch/p_2_in [15]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [15]),
        .O(\pc0[15]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000A808)) 
    \pc0[15]_i_4 
       (.I0(fch_heir_nir_i_2_n_0),
        .I1(\fch/fch_issu1_fl ),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_issu1 ),
        .I4(\fch/stat [1]),
        .I5(fch_heir_nir_i_3_n_0),
        .O(\pc0[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[15]_i_5 
       (.I0(\fch/p_2_in [15]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[15]_INST_0_i_4_n_5 ),
        .O(\pc0[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0222222200000000)) 
    \pc0[15]_i_6 
       (.I0(\fch/fch_issu1 ),
        .I1(\fch/ctl_bcc_take0_fl ),
        .I2(stat[0]),
        .I3(stat[2]),
        .I4(stat[1]),
        .I5(\fadr[15]_INST_0_i_15_n_0 ),
        .O(\pc0[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h08000888)) 
    \pc0[15]_i_7 
       (.I0(\fadr[15]_INST_0_i_7_n_0 ),
        .I1(\fadr[15]_INST_0_i_6_n_0 ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(\fch/fch_issu1_ir ),
        .O(\pc0[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \pc0[15]_i_8 
       (.I0(\fadr[15]_INST_0_i_6_n_0 ),
        .I1(\fch/fch_issu1_ir ),
        .I2(\fch/stat [2]),
        .I3(\fch/stat [0]),
        .I4(\fadr[15]_INST_0_i_8_n_0 ),
        .O(\pc0[15]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[1]_i_1 
       (.I0(\pc0[1]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [1]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[1]_i_3_n_0 ),
        .O(fch_pc[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[1]_i_2 
       (.I0(\fch/p_2_in [1]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [1]),
        .O(\pc0[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[1]_i_3 
       (.I0(\fch/p_2_in [1]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[4]_INST_0_i_1_n_7 ),
        .O(\pc0[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[2]_i_1 
       (.I0(\pc0[2]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [2]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[2]_i_3_n_0 ),
        .O(fch_pc[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[2]_i_2 
       (.I0(\fch/p_2_in [2]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [2]),
        .O(\pc0[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[2]_i_3 
       (.I0(\fch/p_2_in [2]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[4]_INST_0_i_1_n_6 ),
        .O(\pc0[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[3]_i_1 
       (.I0(\pc0[3]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [3]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[3]_i_4_n_0 ),
        .O(fch_pc[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[3]_i_2 
       (.I0(\fch/p_2_in [3]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [3]),
        .O(\pc0[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[3]_i_4 
       (.I0(\fch/p_2_in [3]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[4]_INST_0_i_1_n_5 ),
        .O(\pc0[3]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \pc0[3]_i_5 
       (.I0(\rgf/pcnt/pc [2]),
        .O(\pc0[3]_i_5_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \pc0[3]_i_6 
       (.I0(\rgf/pcnt/pc [1]),
        .O(\pc0[3]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[4]_i_1 
       (.I0(\pc0[4]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [4]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[4]_i_3_n_0 ),
        .O(fch_pc[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[4]_i_2 
       (.I0(\fch/p_2_in [4]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [4]),
        .O(\pc0[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[4]_i_3 
       (.I0(\fch/p_2_in [4]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[4]_INST_0_i_1_n_4 ),
        .O(\pc0[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[5]_i_1 
       (.I0(\pc0[5]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [5]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[5]_i_3_n_0 ),
        .O(fch_pc[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[5]_i_2 
       (.I0(\fch/p_2_in [5]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [5]),
        .O(\pc0[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[5]_i_3 
       (.I0(\fch/p_2_in [5]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[8]_INST_0_i_1_n_7 ),
        .O(\pc0[5]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[6]_i_1 
       (.I0(\pc0[6]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [6]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[6]_i_3_n_0 ),
        .O(fch_pc[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[6]_i_2 
       (.I0(\fch/p_2_in [6]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [6]),
        .O(\pc0[6]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[6]_i_3 
       (.I0(\fch/p_2_in [6]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[8]_INST_0_i_1_n_6 ),
        .O(\pc0[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[7]_i_1 
       (.I0(\pc0[7]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [7]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[7]_i_4_n_0 ),
        .O(fch_pc[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[7]_i_2 
       (.I0(\fch/p_2_in [7]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [7]),
        .O(\pc0[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[7]_i_4 
       (.I0(\fch/p_2_in [7]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[8]_INST_0_i_1_n_5 ),
        .O(\pc0[7]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[8]_i_1 
       (.I0(\pc0[8]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [8]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[8]_i_3_n_0 ),
        .O(fch_pc[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[8]_i_2 
       (.I0(\fch/p_2_in [8]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [8]),
        .O(\pc0[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[8]_i_3 
       (.I0(\fch/p_2_in [8]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[8]_INST_0_i_1_n_4 ),
        .O(\pc0[8]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc0[9]_i_1 
       (.I0(\pc0[9]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [9]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[9]_i_3_n_0 ),
        .O(fch_pc[9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \pc0[9]_i_2 
       (.I0(\fch/p_2_in [9]),
        .I1(\pc0[15]_i_6_n_0 ),
        .I2(\rgf/pcnt/pc [9]),
        .O(\pc0[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAA0200AAAA)) 
    \pc0[9]_i_3 
       (.I0(\fch/p_2_in [9]),
        .I1(\pc0[15]_i_7_n_0 ),
        .I2(\fadr[15]_INST_0_i_9_n_0 ),
        .I3(\pc0[15]_i_8_n_0 ),
        .I4(\fadr[15]_INST_0_i_5_n_0 ),
        .I5(\fadr[12]_INST_0_i_1_n_7 ),
        .O(\pc0[9]_i_3_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[11]_i_3 
       (.CI(\pc0_reg[7]_i_3_n_0 ),
        .CO({\pc0_reg[11]_i_3_n_0 ,\pc0_reg[11]_i_3_n_1 ,\pc0_reg[11]_i_3_n_2 ,\pc0_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in0_in [11:8]),
        .S(\rgf/pcnt/pc [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[15]_i_3 
       (.CI(\pc0_reg[11]_i_3_n_0 ),
        .CO({\pc0_reg[15]_i_3_n_1 ,\pc0_reg[15]_i_3_n_2 ,\pc0_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in0_in [15:12]),
        .S(\rgf/pcnt/pc [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[3]_i_3 
       (.CI(\<const0> ),
        .CO({\pc0_reg[3]_i_3_n_0 ,\pc0_reg[3]_i_3_n_1 ,\pc0_reg[3]_i_3_n_2 ,\pc0_reg[3]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rgf/pcnt/pc [2:1],\<const0> }),
        .O({\fch/p_2_in0_in [3:1],\NLW_pc0_reg[3]_i_3_O_UNCONNECTED [0]}),
        .S({\rgf/pcnt/pc [3],\pc0[3]_i_5_n_0 ,\pc0[3]_i_6_n_0 ,\rgf/pcnt/pc [0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc0_reg[7]_i_3 
       (.CI(\pc0_reg[3]_i_3_n_0 ),
        .CO({\pc0_reg[7]_i_3_n_0 ,\pc0_reg[7]_i_3_n_1 ,\pc0_reg[7]_i_3_n_2 ,\pc0_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\fch/p_2_in0_in [7:4]),
        .S(\rgf/pcnt/pc [7:4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_2 
       (.I0(\pc0[11]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [11]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[11]_i_4_n_0 ),
        .O(\pc1[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_3 
       (.I0(\pc0[10]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [10]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[10]_i_3_n_0 ),
        .O(\pc1[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_4 
       (.I0(\pc0[9]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [9]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[9]_i_3_n_0 ),
        .O(\pc1[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[11]_i_5 
       (.I0(\pc0[8]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [8]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[8]_i_3_n_0 ),
        .O(\pc1[11]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_2 
       (.I0(\pc0[15]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [15]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[15]_i_5_n_0 ),
        .O(\pc1[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_3 
       (.I0(\pc0[14]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [14]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[14]_i_3_n_0 ),
        .O(\pc1[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_4 
       (.I0(\pc0[13]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [13]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[13]_i_3_n_0 ),
        .O(\pc1[15]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[15]_i_5 
       (.I0(\pc0[12]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [12]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[12]_i_3_n_0 ),
        .O(\pc1[15]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[3]_i_2 
       (.I0(\pc0[3]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [3]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[3]_i_4_n_0 ),
        .O(\pc1[3]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[3]_i_3 
       (.I0(\pc0[2]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [2]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[2]_i_3_n_0 ),
        .O(\pc1[3]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h111DDD1D)) 
    \pc1[3]_i_4 
       (.I0(\pc1[3]_i_6_n_0 ),
        .I1(fch_irq_req),
        .I2(\rgf/pcnt/pc [1]),
        .I3(\pc0[15]_i_6_n_0 ),
        .I4(\fch/p_2_in [1]),
        .O(\pc1[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hBA8A)) 
    \pc1[3]_i_5 
       (.I0(\rgf/pcnt/pc [0]),
        .I1(fch_irq_req),
        .I2(\pc0[15]_i_4_n_0 ),
        .I3(\fch/p_2_in0_in [0]),
        .O(\pc1[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[3]_i_6 
       (.I0(\fch/p_2_in0_in [1]),
        .I1(\pc0[15]_i_4_n_0 ),
        .I2(\fch/p_2_in [1]),
        .I3(\pc1[3]_i_7_n_0 ),
        .I4(\fadr[4]_INST_0_i_1_n_7 ),
        .O(\pc1[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h008C00BFFFFFFFFF)) 
    \pc1[3]_i_7 
       (.I0(\pc1[3]_i_8_n_0 ),
        .I1(\fadr[15]_INST_0_i_6_n_0 ),
        .I2(\fadr[15]_INST_0_i_7_n_0 ),
        .I3(\fadr[15]_INST_0_i_9_n_0 ),
        .I4(\fadr[15]_INST_0_i_11_n_0 ),
        .I5(\fadr[15]_INST_0_i_5_n_0 ),
        .O(\pc1[3]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \pc1[3]_i_8 
       (.I0(\fch/fch_issu1 ),
        .I1(\fch/fch_term_fl ),
        .I2(\fch/fch_issu1_fl ),
        .I3(\fch/stat [1]),
        .I4(\fch/stat [0]),
        .O(\pc1[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_2 
       (.I0(\pc0[7]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [7]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[7]_i_4_n_0 ),
        .O(\pc1[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_3 
       (.I0(\pc0[6]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [6]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[6]_i_3_n_0 ),
        .O(\pc1[7]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_4 
       (.I0(\pc0[5]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [5]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[5]_i_3_n_0 ),
        .O(\pc1[7]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \pc1[7]_i_5 
       (.I0(\pc0[4]_i_2_n_0 ),
        .I1(fch_irq_req),
        .I2(\fch/p_2_in0_in [4]),
        .I3(\pc0[15]_i_4_n_0 ),
        .I4(\pc0[4]_i_3_n_0 ),
        .O(\pc1[7]_i_5_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[11]_i_1 
       (.CI(\pc1_reg[7]_i_1_n_0 ),
        .CO({\pc1_reg[11]_i_1_n_0 ,\pc1_reg[11]_i_1_n_1 ,\pc1_reg[11]_i_1_n_2 ,\pc1_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\pc1_reg[11]_i_1_n_4 ,\pc1_reg[11]_i_1_n_5 ,\pc1_reg[11]_i_1_n_6 ,\pc1_reg[11]_i_1_n_7 }),
        .S({\pc1[11]_i_2_n_0 ,\pc1[11]_i_3_n_0 ,\pc1[11]_i_4_n_0 ,\pc1[11]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[15]_i_1 
       (.CI(\pc1_reg[11]_i_1_n_0 ),
        .CO({\pc1_reg[15]_i_1_n_1 ,\pc1_reg[15]_i_1_n_2 ,\pc1_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\pc1_reg[15]_i_1_n_4 ,\pc1_reg[15]_i_1_n_5 ,\pc1_reg[15]_i_1_n_6 ,\pc1_reg[15]_i_1_n_7 }),
        .S({\pc1[15]_i_2_n_0 ,\pc1[15]_i_3_n_0 ,\pc1[15]_i_4_n_0 ,\pc1[15]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\pc1_reg[3]_i_1_n_0 ,\pc1_reg[3]_i_1_n_1 ,\pc1_reg[3]_i_1_n_2 ,\pc1_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,fch_pc[1],\<const0> }),
        .O({\pc1_reg[3]_i_1_n_4 ,\pc1_reg[3]_i_1_n_5 ,\pc1_reg[3]_i_1_n_6 ,\pc1_reg[3]_i_1_n_7 }),
        .S({\pc1[3]_i_2_n_0 ,\pc1[3]_i_3_n_0 ,\pc1[3]_i_4_n_0 ,\pc1[3]_i_5_n_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc1_reg[7]_i_1 
       (.CI(\pc1_reg[3]_i_1_n_0 ),
        .CO({\pc1_reg[7]_i_1_n_0 ,\pc1_reg[7]_i_1_n_1 ,\pc1_reg[7]_i_1_n_2 ,\pc1_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\pc1_reg[7]_i_1_n_4 ,\pc1_reg[7]_i_1_n_5 ,\pc1_reg[7]_i_1_n_6 ,\pc1_reg[7]_i_1_n_7 }),
        .S({\pc1[7]_i_2_n_0 ,\pc1[7]_i_3_n_0 ,\pc1[7]_i_4_n_0 ,\pc1[7]_i_5_n_0 }));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[0]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/rgf_c1bus_0 [0]),
        .I4(\pc[0]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[0]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[0]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [0]),
        .O(\rgf/rgf_c1bus_0 [0]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[0]_i_3 
       (.I0(fch_pc[0]),
        .I1(\rgf/pcnt/pc [0]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[10]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/rgf_c1bus_0 [10]),
        .I4(\pc[10]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [10]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[10]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[10]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [10]),
        .O(\rgf/rgf_c1bus_0 [10]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[10]_i_3 
       (.I0(fch_pc[10]),
        .I1(\rgf/pcnt/pc [10]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[10]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[11]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/rgf_c1bus_0 [11]),
        .I4(\pc[11]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[11]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[11]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [11]),
        .O(\rgf/rgf_c1bus_0 [11]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[11]_i_3 
       (.I0(fch_pc[11]),
        .I1(\rgf/pcnt/pc [11]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[11]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[12]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/rgf_c1bus_0 [12]),
        .I4(\pc[12]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[12]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [12]),
        .O(\rgf/rgf_c0bus_0 [12]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[12]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[12]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [12]),
        .O(\rgf/rgf_c1bus_0 [12]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[12]_i_4 
       (.I0(fch_pc[12]),
        .I1(\rgf/pcnt/pc [12]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[12]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[13]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/rgf_c1bus_0 [13]),
        .I4(\pc[13]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[13]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [13]),
        .O(\rgf/rgf_c0bus_0 [13]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[13]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[13]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [13]),
        .O(\rgf/rgf_c1bus_0 [13]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[13]_i_4 
       (.I0(fch_pc[13]),
        .I1(\rgf/pcnt/pc [13]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[13]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[14]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/rgf_c1bus_0 [14]),
        .I4(\pc[14]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[14]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [14]),
        .O(\rgf/rgf_c0bus_0 [14]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[14]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[14]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [14]),
        .O(\rgf/rgf_c1bus_0 [14]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[14]_i_4 
       (.I0(fch_pc[14]),
        .I1(\rgf/pcnt/pc [14]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[14]_i_4_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \pc[15]_i_1 
       (.I0(rst_n),
        .O(\alu1/div/p_0_in__0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_10 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(ctl_selc0_rn),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_rn_wb [0]),
        .O(\rgf/rctl/p_0_in [0]));
  LUT6 #(
    .INIT(64'hE4E0A0E0FFFFFFFF)) 
    \pc[15]_i_11 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(ctl_selc0[0]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_wb [0]),
        .I5(\rgf/rctl/p_0_in [4]),
        .O(\pc[15]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \pc[15]_i_12 
       (.I0(fch_term),
        .I1(ctl_fetch_lng0),
        .I2(ctl_fetch_ext0),
        .I3(ctl_fetch_lng1),
        .I4(ctl_fetch_ext1),
        .O(\pc[15]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_13 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(ctl_selc0[1]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_wb [1]),
        .O(\rgf/rctl/p_0_in [4]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[15]_i_2 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/rgf_c1bus_0 [15]),
        .I4(\pc[15]_i_7_n_0 ),
        .O(\rgf/pcnt/p_1_in [15]));
  LUT4 #(
    .INIT(16'h0010)) 
    \pc[15]_i_3 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_11_n_0 ),
        .O(\rgf/c0bus_sel_cr [1]));
  LUT5 #(
    .INIT(32'h00001000)) 
    \pc[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1 [1]),
        .I4(\rgf/rctl/rgf_selc1 [0]),
        .O(\rgf/c1bus_sel_cr [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_5 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[15]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [15]),
        .O(\rgf/rgf_c0bus_0 [15]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_6 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[15]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [15]),
        .O(\rgf/rgf_c1bus_0 [15]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[15]_i_7 
       (.I0(fch_pc[15]),
        .I1(\rgf/pcnt/pc [15]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_8 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\rgf_selc0_rn_wb[1]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_rn_wb [1]),
        .O(\rgf/rctl/p_0_in [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[15]_i_9 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\rgf_selc0_rn_wb[2]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_selc0_rn_wb [2]),
        .O(\rgf/rctl/p_0_in [2]));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[1]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/rgf_c1bus_0 [1]),
        .I4(\pc[1]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [1]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[1]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[1]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [1]),
        .O(\rgf/rgf_c1bus_0 [1]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[1]_i_3 
       (.I0(fch_pc[1]),
        .I1(\rgf/pcnt/pc [1]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[2]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/rgf_c1bus_0 [2]),
        .I4(\pc[2]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[2]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[2]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [2]),
        .O(\rgf/rgf_c0bus_0 [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[2]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[2]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [2]),
        .O(\rgf/rgf_c1bus_0 [2]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[2]_i_4 
       (.I0(fch_pc[2]),
        .I1(\rgf/pcnt/pc [2]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[2]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[3]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/rgf_c1bus_0 [3]),
        .I4(\pc[3]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[3]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[3]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [3]),
        .O(\rgf/rgf_c0bus_0 [3]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[3]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[3]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [3]),
        .O(\rgf/rgf_c1bus_0 [3]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[3]_i_4 
       (.I0(fch_pc[3]),
        .I1(\rgf/pcnt/pc [3]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[3]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[4]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/rgf_c1bus_0 [4]),
        .I4(\pc[4]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [4]));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \pc[4]_i_10 
       (.I0(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\pc[4]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \pc[4]_i_11 
       (.I0(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I3(\pc[4]_i_13_n_0 ),
        .O(\pc[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0D0800000F0F0F0F)) 
    \pc[4]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_25_n_0 ),
        .O(\pc[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000C880C440CCC0C)) 
    \pc[4]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_28_n_0 ),
        .O(\pc[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \pc[4]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\pc[4]_i_5_n_0 ),
        .I3(\pc[4]_i_6_n_0 ),
        .I4(\rgf/rctl/rgf_selc0_stat ),
        .I5(\rgf/rctl/rgf_c0bus_wb [4]),
        .O(\rgf/rgf_c0bus_0 [4]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[4]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[4]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [4]),
        .O(\rgf/rgf_c1bus_0 [4]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[4]_i_4 
       (.I0(fch_pc[4]),
        .I1(\rgf/pcnt/pc [4]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[4]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFEEEE)) 
    \pc[4]_i_5 
       (.I0(\rgf_c0bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .I2(\pc[4]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_2_n_0 ),
        .O(\pc[4]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \pc[4]_i_6 
       (.I0(cbus_i[4]),
        .I1(ccmd[4]),
        .O(\pc[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1F100FFFFFFFF)) 
    \pc[4]_i_7 
       (.I0(\pc[4]_i_8_n_0 ),
        .I1(\pc[4]_i_9_n_0 ),
        .I2(\pc[4]_i_10_n_0 ),
        .I3(\pc[4]_i_11_n_0 ),
        .I4(\pc[4]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\pc[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h4444F44444F4F4F4)) 
    \pc[4]_i_8 
       (.I0(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_13_n_0 ),
        .O(\pc[4]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \pc[4]_i_9 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .O(\pc[4]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[5]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/rgf_c1bus_0 [5]),
        .I4(\pc[5]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [5]));
  LUT2 #(
    .INIT(4'h1)) 
    \pc[5]_i_10 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_20_n_0 ),
        .O(\pc[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \pc[5]_i_11 
       (.I0(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\pc[5]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \pc[5]_i_12 
       (.I0(\rgf_c0bus_wb[5]_i_20_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_18_n_0 ),
        .I3(\pc[5]_i_15_n_0 ),
        .O(\pc[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0D0800000F0F0F0F)) 
    \pc[5]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_28_n_0 ),
        .O(\pc[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \pc[5]_i_14 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\pc[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h000C880C440CCC0C)) 
    \pc[5]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[21]_i_27_n_0 ),
        .O(\pc[5]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \pc[5]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\pc[5]_i_5_n_0 ),
        .I3(\pc[5]_i_6_n_0 ),
        .I4(\rgf/rctl/rgf_selc0_stat ),
        .I5(\rgf/rctl/rgf_c0bus_wb [5]),
        .O(\rgf/rgf_c0bus_0 [5]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[5]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[5]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [5]),
        .O(\rgf/rgf_c1bus_0 [5]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[5]_i_4 
       (.I0(fch_pc[5]),
        .I1(\rgf/pcnt/pc [5]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEFEEEE)) 
    \pc[5]_i_5 
       (.I0(\rgf_c0bus_wb[5]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .I2(\pc[5]_i_7_n_0 ),
        .I3(\pc[5]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_2_n_0 ),
        .O(\pc[5]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \pc[5]_i_6 
       (.I0(cbus_i[5]),
        .I1(ccmd[4]),
        .O(\pc[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF1F1F100FFFFFFFF)) 
    \pc[5]_i_7 
       (.I0(\pc[5]_i_9_n_0 ),
        .I1(\pc[5]_i_10_n_0 ),
        .I2(\pc[5]_i_11_n_0 ),
        .I3(\pc[5]_i_12_n_0 ),
        .I4(\pc[5]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\pc[5]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \pc[5]_i_8 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\pc[5]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_15_n_0 ),
        .O(\pc[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4444F44444F4F4F4)) 
    \pc[5]_i_9 
       (.I0(\rgf_c0bus_wb[5]_i_18_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[21]_i_13_n_0 ),
        .O(\pc[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[6]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/rgf_c1bus_0 [6]),
        .I4(\pc[6]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [6]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[6]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[6]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [6]),
        .O(\rgf/rgf_c1bus_0 [6]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[6]_i_3 
       (.I0(fch_pc[6]),
        .I1(\rgf/pcnt/pc [6]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[7]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/rgf_c1bus_0 [7]),
        .I4(\pc[7]_i_4_n_0 ),
        .O(\rgf/pcnt/p_1_in [7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[7]_i_2 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[7]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [7]),
        .O(\rgf/rgf_c0bus_0 [7]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[7]_i_3 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[7]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [7]),
        .O(\rgf/rgf_c1bus_0 [7]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[7]_i_4 
       (.I0(fch_pc[7]),
        .I1(\rgf/pcnt/pc [7]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[7]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[8]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/rgf_c1bus_0 [8]),
        .I4(\pc[8]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [8]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[8]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[8]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [8]),
        .O(\rgf/rgf_c1bus_0 [8]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[8]_i_3 
       (.I0(fch_pc[8]),
        .I1(\rgf/pcnt/pc [8]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[8]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEC20)) 
    \pc[9]_i_1 
       (.I0(\rgf/c0bus_sel_cr [1]),
        .I1(\rgf/c1bus_sel_cr [1]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/rgf_c1bus_0 [9]),
        .I4(\pc[9]_i_3_n_0 ),
        .O(\rgf/pcnt/p_1_in [9]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \pc[9]_i_2 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[9]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [9]),
        .O(\rgf/rgf_c1bus_0 [9]));
  LUT5 #(
    .INIT(32'h000A000C)) 
    \pc[9]_i_3 
       (.I0(fch_pc[9]),
        .I1(\rgf/pcnt/pc [9]),
        .I2(\rgf/c0bus_sel_cr [1]),
        .I3(\rgf/c1bus_sel_cr [1]),
        .I4(\pc[15]_i_12_n_0 ),
        .O(\pc[9]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[0]_i_1 
       (.I0(\alu0/div/add_out [0]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_in0 ),
        .O(\alu0/div/p_2_in [0]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[0]_i_1__0 
       (.I0(\alu1/div/add_out [0]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_in0 ),
        .O(\alu1/div/p_2_in [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[10]_i_1 
       (.I0(\alu0/div/add_out [10]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [6]),
        .O(\alu0/div/p_2_in [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[10]_i_1__0 
       (.I0(\alu1/div/add_out [10]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [6]),
        .O(\alu1/div/p_2_in [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[11]_i_1 
       (.I0(\alu0/div/add_out [11]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [7]),
        .O(\alu0/div/p_2_in [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[11]_i_1__0 
       (.I0(\alu1/div/add_out [11]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [7]),
        .O(\alu1/div/p_2_in [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[12]_i_1 
       (.I0(\alu0/div/add_out [12]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [8]),
        .O(\alu0/div/p_2_in [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[12]_i_1__0 
       (.I0(\alu1/div/add_out [12]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [8]),
        .O(\alu1/div/p_2_in [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[13]_i_1 
       (.I0(\alu0/div/add_out [13]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [9]),
        .O(\alu0/div/p_2_in [13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[13]_i_1__0 
       (.I0(\alu1/div/add_out [13]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [9]),
        .O(\alu1/div/p_2_in [13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[14]_i_1 
       (.I0(\alu0/div/add_out [14]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [10]),
        .O(\alu0/div/p_2_in [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[14]_i_1__0 
       (.I0(\alu1/div/add_out [14]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [10]),
        .O(\alu1/div/p_2_in [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[15]_i_1 
       (.I0(\alu0/div/add_out [15]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [11]),
        .O(\alu0/div/p_2_in [15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[15]_i_1__0 
       (.I0(\alu1/div/add_out [15]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [11]),
        .O(\alu1/div/p_2_in [15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[16]_i_1 
       (.I0(\alu0/div/add_out [16]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [12]),
        .O(\alu0/div/p_2_in [16]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[16]_i_1__0 
       (.I0(\alu1/div/add_out [16]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [12]),
        .O(\alu1/div/p_2_in [16]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[17]_i_1 
       (.I0(\alu0/div/add_out [17]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [13]),
        .O(\alu0/div/p_2_in [17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[17]_i_1__0 
       (.I0(\alu1/div/add_out [17]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [13]),
        .O(\alu1/div/p_2_in [17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[18]_i_1 
       (.I0(\alu0/div/add_out [18]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [14]),
        .O(\alu0/div/p_2_in [18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[18]_i_1__0 
       (.I0(\alu1/div/add_out [18]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [14]),
        .O(\alu1/div/p_2_in [18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[19]_i_1 
       (.I0(\alu0/div/add_out [19]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [15]),
        .O(\alu0/div/p_2_in [19]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[19]_i_1__0 
       (.I0(\alu1/div/add_out [19]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [15]),
        .O(\alu1/div/p_2_in [19]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[1]_i_1 
       (.I0(\alu0/div/add_out [1]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/rem1 ),
        .O(\alu0/div/p_2_in [1]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[1]_i_1__0 
       (.I0(\alu1/div/add_out [1]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem1 ),
        .O(\alu1/div/p_2_in [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[20]_i_1 
       (.I0(\alu0/div/add_out [20]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [16]),
        .O(\alu0/div/p_2_in [20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[20]_i_1__0 
       (.I0(\alu1/div/add_out [20]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [16]),
        .O(\alu1/div/p_2_in [20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[21]_i_1 
       (.I0(\alu0/div/add_out [21]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [17]),
        .O(\alu0/div/p_2_in [21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[21]_i_1__0 
       (.I0(\alu1/div/add_out [21]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [17]),
        .O(\alu1/div/p_2_in [21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[22]_i_1 
       (.I0(\alu0/div/add_out [22]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [18]),
        .O(\alu0/div/p_2_in [22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[22]_i_1__0 
       (.I0(\alu1/div/add_out [22]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [18]),
        .O(\alu1/div/p_2_in [22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[23]_i_1 
       (.I0(\alu0/div/add_out [23]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [19]),
        .O(\alu0/div/p_2_in [23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[23]_i_1__0 
       (.I0(\alu1/div/add_out [23]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [19]),
        .O(\alu1/div/p_2_in [23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[24]_i_1 
       (.I0(\alu0/div/add_out [24]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [20]),
        .O(\alu0/div/p_2_in [24]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[24]_i_1__0 
       (.I0(\alu1/div/add_out [24]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [20]),
        .O(\alu1/div/p_2_in [24]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[25]_i_1 
       (.I0(\alu0/div/add_out [25]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [21]),
        .O(\alu0/div/p_2_in [25]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[25]_i_1__0 
       (.I0(\alu1/div/add_out [25]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [21]),
        .O(\alu1/div/p_2_in [25]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[26]_i_1 
       (.I0(\alu0/div/add_out [26]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [22]),
        .O(\alu0/div/p_2_in [26]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[26]_i_1__0 
       (.I0(\alu1/div/add_out [26]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [22]),
        .O(\alu1/div/p_2_in [26]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[27]_i_1 
       (.I0(\alu0/div/add_out [27]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [23]),
        .O(\alu0/div/p_2_in [27]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[27]_i_1__0 
       (.I0(\alu1/div/add_out [27]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [23]),
        .O(\alu1/div/p_2_in [27]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[28]_i_1 
       (.I0(\alu0/div/add_out [28]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [24]),
        .O(\alu0/div/p_2_in [28]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[28]_i_1__0 
       (.I0(\alu1/div/add_out [28]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [24]),
        .O(\alu1/div/p_2_in [28]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[29]_i_1 
       (.I0(\alu0/div/add_out [29]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [25]),
        .O(\alu0/div/p_2_in [29]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[29]_i_1__0 
       (.I0(\alu1/div/add_out [29]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [25]),
        .O(\alu1/div/p_2_in [29]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[2]_i_1 
       (.I0(\alu0/div/add_out [2]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/rem2 ),
        .O(\alu0/div/p_2_in [2]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[2]_i_1__0 
       (.I0(\alu1/div/add_out [2]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem2 ),
        .O(\alu1/div/p_2_in [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[30]_i_1 
       (.I0(\alu0/div/add_out [30]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [26]),
        .O(\alu0/div/p_2_in [30]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[30]_i_1__0 
       (.I0(\alu1/div/add_out [30]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [26]),
        .O(\alu1/div/p_2_in [30]));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFEE)) 
    \quo[31]_i_1 
       (.I0(\quo[31]_i_3_n_0 ),
        .I1(\quo[31]_i_4_n_0 ),
        .I2(\alu0/div/dctl_stat [3]),
        .I3(\alu0/div/dctl_stat [2]),
        .I4(\alu0/div/dctl_stat [1]),
        .I5(\alu0/div/dctl_stat [0]),
        .O(\quo[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFEE)) 
    \quo[31]_i_1__0 
       (.I0(\quo[31]_i_3__0_n_0 ),
        .I1(\quo[31]_i_4__0_n_0 ),
        .I2(\alu1/div/dctl_stat [3]),
        .I3(\alu1/div/dctl_stat [2]),
        .I4(\alu1/div/dctl_stat [1]),
        .I5(\alu1/div/dctl_stat [0]),
        .O(\quo[31]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[31]_i_2 
       (.I0(\alu0/div/add_out [31]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [27]),
        .O(\alu0/div/p_2_in [31]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[31]_i_2__0 
       (.I0(\alu1/div/add_out [31]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [27]),
        .O(\alu1/div/p_2_in [31]));
  LUT2 #(
    .INIT(4'h2)) 
    \quo[31]_i_3 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\dso[31]_i_4_n_0 ),
        .O(\quo[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \quo[31]_i_3__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\dso[31]_i_4__0_n_0 ),
        .O(\quo[31]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h0200222233223322)) 
    \quo[31]_i_4 
       (.I0(\alu0/div/dctl_stat [0]),
        .I1(\quo[31]_i_5_n_0 ),
        .I2(\alu0/div/den2 ),
        .I3(chg_quo_sgn_i_2_n_0),
        .I4(\alu0/div/dctl/dctl_sign ),
        .I5(\alu0/div/dctl_stat [2]),
        .O(\quo[31]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0200222233223322)) 
    \quo[31]_i_4__0 
       (.I0(\alu1/div/dctl_stat [0]),
        .I1(\quo[31]_i_5__0_n_0 ),
        .I2(\alu1/div/den2 ),
        .I3(chg_quo_sgn_i_2__0_n_0),
        .I4(\alu1/div/dctl/dctl_sign ),
        .I5(\alu1/div/dctl_stat [2]),
        .O(\quo[31]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \quo[31]_i_5 
       (.I0(\alu0/div/dctl_stat [1]),
        .I1(\alu0/div/dctl_stat [3]),
        .O(\quo[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \quo[31]_i_5__0 
       (.I0(\alu1/div/dctl_stat [1]),
        .I1(\alu1/div/dctl_stat [3]),
        .O(\quo[31]_i_5__0_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[3]_i_1 
       (.I0(\alu0/div/add_out [3]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/rem3 ),
        .O(\alu0/div/p_2_in [3]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[3]_i_1__0 
       (.I0(\alu1/div/add_out [3]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem3 ),
        .O(\alu1/div/p_2_in [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[4]_i_1 
       (.I0(\alu0/div/add_out [4]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [0]),
        .O(\alu0/div/p_2_in [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[4]_i_1__0 
       (.I0(\alu1/div/add_out [4]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [0]),
        .O(\alu1/div/p_2_in [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[5]_i_1 
       (.I0(\alu0/div/add_out [5]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [1]),
        .O(\alu0/div/p_2_in [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[5]_i_1__0 
       (.I0(\alu1/div/add_out [5]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [1]),
        .O(\alu1/div/p_2_in [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[6]_i_1 
       (.I0(\alu0/div/add_out [6]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [2]),
        .O(\alu0/div/p_2_in [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[6]_i_1__0 
       (.I0(\alu1/div/add_out [6]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [2]),
        .O(\alu1/div/p_2_in [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[7]_i_1 
       (.I0(\alu0/div/add_out [7]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [3]),
        .O(\alu0/div/p_2_in [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[7]_i_1__0 
       (.I0(\alu1/div/add_out [7]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [3]),
        .O(\alu1/div/p_2_in [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[8]_i_1 
       (.I0(\alu0/div/add_out [8]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [4]),
        .O(\alu0/div/p_2_in [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[8]_i_1__0 
       (.I0(\alu1/div/add_out [8]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [4]),
        .O(\alu1/div/p_2_in [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[9]_i_1 
       (.I0(\alu0/div/add_out [9]),
        .I1(\quo[31]_i_3_n_0 ),
        .I2(\alu0/div/quo [5]),
        .O(\alu0/div/p_2_in [9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[9]_i_1__0 
       (.I0(\alu1/div/add_out [9]),
        .I1(\quo[31]_i_3__0_n_0 ),
        .I2(\alu1/div/quo [5]),
        .O(\alu1/div/p_2_in [9]));
  LUT1 #(
    .INIT(2'h1)) 
    \read_cyc[3]_i_1 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(\mem/mem_accslot ));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_1
       (.I0(\alu0/div/rem1__0 [7]),
        .I1(\alu0/div/dso_0 [7]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_1__0
       (.I0(\alu1/div/rem1__0 [7]),
        .I1(\alu1/div/dso_0 [7]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_2
       (.I0(\alu0/div/rem1__0 [6]),
        .I1(\alu0/div/dso_0 [6]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_2__0
       (.I0(\alu1/div/rem1__0 [6]),
        .I1(\alu1/div/dso_0 [6]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_3
       (.I0(\alu0/div/rem1__0 [5]),
        .I1(\alu0/div/dso_0 [5]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_3__0
       (.I0(\alu1/div/rem1__0 [5]),
        .I1(\alu1/div/dso_0 [5]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_4
       (.I0(\alu0/div/rem1__0 [4]),
        .I1(\alu0/div/dso_0 [4]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_4__0
       (.I0(\alu1/div/rem1__0 [4]),
        .I1(\alu1/div/dso_0 [4]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__0_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_1
       (.I0(\alu0/div/rem1__0 [11]),
        .I1(\alu0/div/dso_0 [11]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_1__0
       (.I0(\alu1/div/rem1__0 [11]),
        .I1(\alu1/div/dso_0 [11]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_2
       (.I0(\alu0/div/rem1__0 [10]),
        .I1(\alu0/div/dso_0 [10]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_2__0
       (.I0(\alu1/div/rem1__0 [10]),
        .I1(\alu1/div/dso_0 [10]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_3
       (.I0(\alu0/div/rem1__0 [9]),
        .I1(\alu0/div/dso_0 [9]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_3__0
       (.I0(\alu1/div/rem1__0 [9]),
        .I1(\alu1/div/dso_0 [9]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_4
       (.I0(\alu0/div/rem1__0 [8]),
        .I1(\alu0/div/dso_0 [8]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_4__0
       (.I0(\alu1/div/rem1__0 [8]),
        .I1(\alu1/div/dso_0 [8]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__1_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_1
       (.I0(\alu0/div/rem1__0 [15]),
        .I1(\alu0/div/rem1 ),
        .I2(\alu0/div/dso_0 [15]),
        .O(rem0_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_1__0
       (.I0(\alu1/div/rem1__0 [15]),
        .I1(\alu1/div/rem1 ),
        .I2(\alu1/div/dso_0 [15]),
        .O(rem0_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_2
       (.I0(\alu0/div/rem1__0 [14]),
        .I1(\alu0/div/dso_0 [14]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_2__0
       (.I0(\alu1/div/rem1__0 [14]),
        .I1(\alu1/div/dso_0 [14]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_3
       (.I0(\alu0/div/rem1__0 [13]),
        .I1(\alu0/div/dso_0 [13]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_3__0
       (.I0(\alu1/div/rem1__0 [13]),
        .I1(\alu1/div/dso_0 [13]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_4
       (.I0(\alu0/div/rem1__0 [12]),
        .I1(\alu0/div/dso_0 [12]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_4__0
       (.I0(\alu1/div/rem1__0 [12]),
        .I1(\alu1/div/dso_0 [12]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__2_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_1
       (.I0(\alu0/div/rem1__0 [19]),
        .I1(\alu0/div/dso_0 [19]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_1__0
       (.I0(\alu1/div/rem1__0 [19]),
        .I1(\alu1/div/dso_0 [19]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_2
       (.I0(\alu0/div/rem1__0 [18]),
        .I1(\alu0/div/dso_0 [18]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_2__0
       (.I0(\alu1/div/rem1__0 [18]),
        .I1(\alu1/div/dso_0 [18]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_3
       (.I0(\alu0/div/rem1__0 [17]),
        .I1(\alu0/div/dso_0 [17]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_3__0
       (.I0(\alu1/div/rem1__0 [17]),
        .I1(\alu1/div/dso_0 [17]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_4
       (.I0(\alu0/div/rem1__0 [16]),
        .I1(\alu0/div/dso_0 [16]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_4__0
       (.I0(\alu1/div/rem1__0 [16]),
        .I1(\alu1/div/dso_0 [16]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__3_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_1
       (.I0(\alu0/div/rem1__0 [23]),
        .I1(\alu0/div/dso_0 [23]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_1__0
       (.I0(\alu1/div/rem1__0 [23]),
        .I1(\alu1/div/dso_0 [23]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__4_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_2
       (.I0(\alu0/div/rem1__0 [22]),
        .I1(\alu0/div/dso_0 [22]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_2__0
       (.I0(\alu1/div/rem1__0 [22]),
        .I1(\alu1/div/dso_0 [22]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__4_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_3
       (.I0(\alu0/div/rem1__0 [21]),
        .I1(\alu0/div/dso_0 [21]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_3__0
       (.I0(\alu1/div/rem1__0 [21]),
        .I1(\alu1/div/dso_0 [21]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__4_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_4
       (.I0(\alu0/div/rem1__0 [20]),
        .I1(\alu0/div/dso_0 [20]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_4__0
       (.I0(\alu1/div/rem1__0 [20]),
        .I1(\alu1/div/dso_0 [20]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__4_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_1
       (.I0(\alu0/div/rem1__0 [27]),
        .I1(\alu0/div/dso_0 [27]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_1__0
       (.I0(\alu1/div/rem1__0 [27]),
        .I1(\alu1/div/dso_0 [27]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__5_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_2
       (.I0(\alu0/div/rem1__0 [26]),
        .I1(\alu0/div/dso_0 [26]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_2__0
       (.I0(\alu1/div/rem1__0 [26]),
        .I1(\alu1/div/dso_0 [26]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__5_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_3
       (.I0(\alu0/div/rem1__0 [25]),
        .I1(\alu0/div/dso_0 [25]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_3__0
       (.I0(\alu1/div/rem1__0 [25]),
        .I1(\alu1/div/dso_0 [25]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__5_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_4
       (.I0(\alu0/div/rem1__0 [24]),
        .I1(\alu0/div/dso_0 [24]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_4__0
       (.I0(\alu1/div/rem1__0 [24]),
        .I1(\alu1/div/dso_0 [24]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__5_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_1
       (.I0(\alu0/div/rem1__0 [31]),
        .I1(\alu0/div/rem1 ),
        .I2(\alu0/div/dso_0 [31]),
        .O(rem0_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_1__0
       (.I0(\alu1/div/rem1__0 [31]),
        .I1(\alu1/div/rem1 ),
        .I2(\alu1/div/dso_0 [31]),
        .O(rem0_carry__6_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_2
       (.I0(\alu0/div/rem1__0 [30]),
        .I1(\alu0/div/dso_0 [30]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_2__0
       (.I0(\alu1/div/rem1__0 [30]),
        .I1(\alu1/div/dso_0 [30]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__6_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_3
       (.I0(\alu0/div/rem1__0 [29]),
        .I1(\alu0/div/dso_0 [29]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_3__0
       (.I0(\alu1/div/rem1__0 [29]),
        .I1(\alu1/div/dso_0 [29]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__6_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_4
       (.I0(\alu0/div/rem1__0 [28]),
        .I1(\alu0/div/dso_0 [28]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry__6_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_4__0
       (.I0(\alu1/div/rem1__0 [28]),
        .I1(\alu1/div/dso_0 [28]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry__6_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem0_carry__7_i_1
       (.I0(\alu0/div/rem1 ),
        .I1(\alu0/div/rem1__0 [32]),
        .O(rem0_carry__7_i_1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem0_carry__7_i_1__0
       (.I0(\alu1/div/rem1 ),
        .I1(\alu1/div/rem1__0 [32]),
        .O(rem0_carry__7_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem0_carry_i_1
       (.I0(\alu0/div/rem1 ),
        .O(rem0_carry_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem0_carry_i_1__0
       (.I0(\alu1/div/rem1 ),
        .O(rem0_carry_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_2
       (.I0(\alu0/div/rem1__0 [3]),
        .I1(\alu0/div/dso_0 [3]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_2__0
       (.I0(\alu1/div/rem1__0 [3]),
        .I1(\alu1/div/dso_0 [3]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_3
       (.I0(\alu0/div/rem1__0 [2]),
        .I1(\alu0/div/dso_0 [2]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_3__0
       (.I0(\alu1/div/rem1__0 [2]),
        .I1(\alu1/div/dso_0 [2]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_4
       (.I0(\alu0/div/rem1__0 [1]),
        .I1(\alu0/div/dso_0 [1]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_4__0
       (.I0(\alu1/div/rem1__0 [1]),
        .I1(\alu1/div/dso_0 [1]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_5
       (.I0(\alu0/div/den [28]),
        .I1(\alu0/div/dso_0 [0]),
        .I2(\alu0/div/rem1 ),
        .O(rem0_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_5__0
       (.I0(\alu1/div/den [28]),
        .I1(\alu1/div/dso_0 [0]),
        .I2(\alu1/div/rem1 ),
        .O(rem0_carry_i_5__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_1
       (.I0(\alu0/div/rem2__0 [7]),
        .I1(\alu0/div/dso_0 [7]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_1__0
       (.I0(\alu1/div/rem2__0 [7]),
        .I1(\alu1/div/dso_0 [7]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_2
       (.I0(\alu0/div/rem2__0 [6]),
        .I1(\alu0/div/dso_0 [6]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_2__0
       (.I0(\alu1/div/rem2__0 [6]),
        .I1(\alu1/div/dso_0 [6]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_3
       (.I0(\alu0/div/rem2__0 [5]),
        .I1(\alu0/div/dso_0 [5]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_3__0
       (.I0(\alu1/div/rem2__0 [5]),
        .I1(\alu1/div/dso_0 [5]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_4
       (.I0(\alu0/div/rem2__0 [4]),
        .I1(\alu0/div/dso_0 [4]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_4__0
       (.I0(\alu1/div/rem2__0 [4]),
        .I1(\alu1/div/dso_0 [4]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__0_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_1
       (.I0(\alu0/div/rem2__0 [11]),
        .I1(\alu0/div/dso_0 [11]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_1__0
       (.I0(\alu1/div/rem2__0 [11]),
        .I1(\alu1/div/dso_0 [11]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_2
       (.I0(\alu0/div/rem2__0 [10]),
        .I1(\alu0/div/dso_0 [10]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_2__0
       (.I0(\alu1/div/rem2__0 [10]),
        .I1(\alu1/div/dso_0 [10]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_3
       (.I0(\alu0/div/rem2__0 [9]),
        .I1(\alu0/div/dso_0 [9]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_3__0
       (.I0(\alu1/div/rem2__0 [9]),
        .I1(\alu1/div/dso_0 [9]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_4
       (.I0(\alu0/div/rem2__0 [8]),
        .I1(\alu0/div/dso_0 [8]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_4__0
       (.I0(\alu1/div/rem2__0 [8]),
        .I1(\alu1/div/dso_0 [8]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__1_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_1
       (.I0(\alu0/div/rem2__0 [15]),
        .I1(\alu0/div/rem2 ),
        .I2(\alu0/div/dso_0 [15]),
        .O(rem1_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_1__0
       (.I0(\alu1/div/rem2__0 [15]),
        .I1(\alu1/div/rem2 ),
        .I2(\alu1/div/dso_0 [15]),
        .O(rem1_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_2
       (.I0(\alu0/div/rem2__0 [14]),
        .I1(\alu0/div/dso_0 [14]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_2__0
       (.I0(\alu1/div/rem2__0 [14]),
        .I1(\alu1/div/dso_0 [14]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_3
       (.I0(\alu0/div/rem2__0 [13]),
        .I1(\alu0/div/dso_0 [13]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_3__0
       (.I0(\alu1/div/rem2__0 [13]),
        .I1(\alu1/div/dso_0 [13]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_4
       (.I0(\alu0/div/rem2__0 [12]),
        .I1(\alu0/div/dso_0 [12]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_4__0
       (.I0(\alu1/div/rem2__0 [12]),
        .I1(\alu1/div/dso_0 [12]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__2_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_1
       (.I0(\alu0/div/rem2__0 [19]),
        .I1(\alu0/div/dso_0 [19]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_1__0
       (.I0(\alu1/div/rem2__0 [19]),
        .I1(\alu1/div/dso_0 [19]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_2
       (.I0(\alu0/div/rem2__0 [18]),
        .I1(\alu0/div/dso_0 [18]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_2__0
       (.I0(\alu1/div/rem2__0 [18]),
        .I1(\alu1/div/dso_0 [18]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_3
       (.I0(\alu0/div/rem2__0 [17]),
        .I1(\alu0/div/dso_0 [17]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_3__0
       (.I0(\alu1/div/rem2__0 [17]),
        .I1(\alu1/div/dso_0 [17]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_4
       (.I0(\alu0/div/rem2__0 [16]),
        .I1(\alu0/div/dso_0 [16]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_4__0
       (.I0(\alu1/div/rem2__0 [16]),
        .I1(\alu1/div/dso_0 [16]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__3_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_1
       (.I0(\alu0/div/rem2__0 [23]),
        .I1(\alu0/div/dso_0 [23]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_1__0
       (.I0(\alu1/div/rem2__0 [23]),
        .I1(\alu1/div/dso_0 [23]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__4_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_2
       (.I0(\alu0/div/rem2__0 [22]),
        .I1(\alu0/div/dso_0 [22]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_2__0
       (.I0(\alu1/div/rem2__0 [22]),
        .I1(\alu1/div/dso_0 [22]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__4_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_3
       (.I0(\alu0/div/rem2__0 [21]),
        .I1(\alu0/div/dso_0 [21]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_3__0
       (.I0(\alu1/div/rem2__0 [21]),
        .I1(\alu1/div/dso_0 [21]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__4_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_4
       (.I0(\alu0/div/rem2__0 [20]),
        .I1(\alu0/div/dso_0 [20]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_4__0
       (.I0(\alu1/div/rem2__0 [20]),
        .I1(\alu1/div/dso_0 [20]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__4_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_1
       (.I0(\alu0/div/rem2__0 [27]),
        .I1(\alu0/div/dso_0 [27]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_1__0
       (.I0(\alu1/div/rem2__0 [27]),
        .I1(\alu1/div/dso_0 [27]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__5_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_2
       (.I0(\alu0/div/rem2__0 [26]),
        .I1(\alu0/div/dso_0 [26]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_2__0
       (.I0(\alu1/div/rem2__0 [26]),
        .I1(\alu1/div/dso_0 [26]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__5_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_3
       (.I0(\alu0/div/rem2__0 [25]),
        .I1(\alu0/div/dso_0 [25]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_3__0
       (.I0(\alu1/div/rem2__0 [25]),
        .I1(\alu1/div/dso_0 [25]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__5_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_4
       (.I0(\alu0/div/rem2__0 [24]),
        .I1(\alu0/div/dso_0 [24]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_4__0
       (.I0(\alu1/div/rem2__0 [24]),
        .I1(\alu1/div/dso_0 [24]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__5_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_1
       (.I0(\alu0/div/rem2__0 [31]),
        .I1(\alu0/div/rem2 ),
        .I2(\alu0/div/dso_0 [31]),
        .O(rem1_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_1__0
       (.I0(\alu1/div/rem2__0 [31]),
        .I1(\alu1/div/rem2 ),
        .I2(\alu1/div/dso_0 [31]),
        .O(rem1_carry__6_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_2
       (.I0(\alu0/div/rem2__0 [30]),
        .I1(\alu0/div/dso_0 [30]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_2__0
       (.I0(\alu1/div/rem2__0 [30]),
        .I1(\alu1/div/dso_0 [30]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__6_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_3
       (.I0(\alu0/div/rem2__0 [29]),
        .I1(\alu0/div/dso_0 [29]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_3__0
       (.I0(\alu1/div/rem2__0 [29]),
        .I1(\alu1/div/dso_0 [29]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__6_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_4
       (.I0(\alu0/div/rem2__0 [28]),
        .I1(\alu0/div/dso_0 [28]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry__6_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_4__0
       (.I0(\alu1/div/rem2__0 [28]),
        .I1(\alu1/div/dso_0 [28]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry__6_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem1_carry__7_i_1
       (.I0(\alu0/div/rem2 ),
        .I1(\alu0/div/rem2__0 [32]),
        .O(rem1_carry__7_i_1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem1_carry__7_i_1__0
       (.I0(\alu1/div/rem2 ),
        .I1(\alu1/div/rem2__0 [32]),
        .O(rem1_carry__7_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem1_carry_i_1
       (.I0(\alu0/div/rem2 ),
        .O(rem1_carry_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem1_carry_i_1__0
       (.I0(\alu1/div/rem2 ),
        .O(rem1_carry_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_2
       (.I0(\alu0/div/rem2__0 [3]),
        .I1(\alu0/div/dso_0 [3]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_2__0
       (.I0(\alu1/div/rem2__0 [3]),
        .I1(\alu1/div/dso_0 [3]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_3
       (.I0(\alu0/div/rem2__0 [2]),
        .I1(\alu0/div/dso_0 [2]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_3__0
       (.I0(\alu1/div/rem2__0 [2]),
        .I1(\alu1/div/dso_0 [2]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_4
       (.I0(\alu0/div/rem2__0 [1]),
        .I1(\alu0/div/dso_0 [1]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_4__0
       (.I0(\alu1/div/rem2__0 [1]),
        .I1(\alu1/div/dso_0 [1]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_5
       (.I0(\alu0/div/den [29]),
        .I1(\alu0/div/dso_0 [0]),
        .I2(\alu0/div/rem2 ),
        .O(rem1_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_5__0
       (.I0(\alu1/div/den [29]),
        .I1(\alu1/div/dso_0 [0]),
        .I2(\alu1/div/rem2 ),
        .O(rem1_carry_i_5__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_1
       (.I0(\alu0/div/rem3__0 [7]),
        .I1(\alu0/div/dso_0 [7]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_1__0
       (.I0(\alu1/div/rem3__0 [7]),
        .I1(\alu1/div/dso_0 [7]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_2
       (.I0(\alu0/div/rem3__0 [6]),
        .I1(\alu0/div/dso_0 [6]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_2__0
       (.I0(\alu1/div/rem3__0 [6]),
        .I1(\alu1/div/dso_0 [6]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_3
       (.I0(\alu0/div/rem3__0 [5]),
        .I1(\alu0/div/dso_0 [5]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_3__0
       (.I0(\alu1/div/rem3__0 [5]),
        .I1(\alu1/div/dso_0 [5]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_4
       (.I0(\alu0/div/rem3__0 [4]),
        .I1(\alu0/div/dso_0 [4]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_4__0
       (.I0(\alu1/div/rem3__0 [4]),
        .I1(\alu1/div/dso_0 [4]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__0_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_1
       (.I0(\alu0/div/rem3__0 [11]),
        .I1(\alu0/div/dso_0 [11]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_1__0
       (.I0(\alu1/div/rem3__0 [11]),
        .I1(\alu1/div/dso_0 [11]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_2
       (.I0(\alu0/div/rem3__0 [10]),
        .I1(\alu0/div/dso_0 [10]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_2__0
       (.I0(\alu1/div/rem3__0 [10]),
        .I1(\alu1/div/dso_0 [10]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_3
       (.I0(\alu0/div/rem3__0 [9]),
        .I1(\alu0/div/dso_0 [9]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_3__0
       (.I0(\alu1/div/rem3__0 [9]),
        .I1(\alu1/div/dso_0 [9]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_4
       (.I0(\alu0/div/rem3__0 [8]),
        .I1(\alu0/div/dso_0 [8]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_4__0
       (.I0(\alu1/div/rem3__0 [8]),
        .I1(\alu1/div/dso_0 [8]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__1_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_1
       (.I0(\alu0/div/rem3__0 [15]),
        .I1(\alu0/div/rem3 ),
        .I2(\alu0/div/dso_0 [15]),
        .O(rem2_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_1__0
       (.I0(\alu1/div/rem3__0 [15]),
        .I1(\alu1/div/rem3 ),
        .I2(\alu1/div/dso_0 [15]),
        .O(rem2_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_2
       (.I0(\alu0/div/rem3__0 [14]),
        .I1(\alu0/div/dso_0 [14]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_2__0
       (.I0(\alu1/div/rem3__0 [14]),
        .I1(\alu1/div/dso_0 [14]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_3
       (.I0(\alu0/div/rem3__0 [13]),
        .I1(\alu0/div/dso_0 [13]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_3__0
       (.I0(\alu1/div/rem3__0 [13]),
        .I1(\alu1/div/dso_0 [13]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_4
       (.I0(\alu0/div/rem3__0 [12]),
        .I1(\alu0/div/dso_0 [12]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_4__0
       (.I0(\alu1/div/rem3__0 [12]),
        .I1(\alu1/div/dso_0 [12]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__2_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_1
       (.I0(\alu0/div/rem3__0 [19]),
        .I1(\alu0/div/dso_0 [19]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_1__0
       (.I0(\alu1/div/rem3__0 [19]),
        .I1(\alu1/div/dso_0 [19]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_2
       (.I0(\alu0/div/rem3__0 [18]),
        .I1(\alu0/div/dso_0 [18]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_2__0
       (.I0(\alu1/div/rem3__0 [18]),
        .I1(\alu1/div/dso_0 [18]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_3
       (.I0(\alu0/div/rem3__0 [17]),
        .I1(\alu0/div/dso_0 [17]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_3__0
       (.I0(\alu1/div/rem3__0 [17]),
        .I1(\alu1/div/dso_0 [17]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_4
       (.I0(\alu0/div/rem3__0 [16]),
        .I1(\alu0/div/dso_0 [16]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_4__0
       (.I0(\alu1/div/rem3__0 [16]),
        .I1(\alu1/div/dso_0 [16]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__3_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_1
       (.I0(\alu0/div/rem3__0 [23]),
        .I1(\alu0/div/dso_0 [23]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_1__0
       (.I0(\alu1/div/rem3__0 [23]),
        .I1(\alu1/div/dso_0 [23]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__4_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_2
       (.I0(\alu0/div/rem3__0 [22]),
        .I1(\alu0/div/dso_0 [22]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_2__0
       (.I0(\alu1/div/rem3__0 [22]),
        .I1(\alu1/div/dso_0 [22]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__4_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_3
       (.I0(\alu0/div/rem3__0 [21]),
        .I1(\alu0/div/dso_0 [21]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_3__0
       (.I0(\alu1/div/rem3__0 [21]),
        .I1(\alu1/div/dso_0 [21]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__4_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_4
       (.I0(\alu0/div/rem3__0 [20]),
        .I1(\alu0/div/dso_0 [20]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_4__0
       (.I0(\alu1/div/rem3__0 [20]),
        .I1(\alu1/div/dso_0 [20]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__4_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_1
       (.I0(\alu0/div/rem3__0 [27]),
        .I1(\alu0/div/dso_0 [27]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_1__0
       (.I0(\alu1/div/rem3__0 [27]),
        .I1(\alu1/div/dso_0 [27]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__5_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_2
       (.I0(\alu0/div/rem3__0 [26]),
        .I1(\alu0/div/dso_0 [26]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_2__0
       (.I0(\alu1/div/rem3__0 [26]),
        .I1(\alu1/div/dso_0 [26]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__5_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_3
       (.I0(\alu0/div/rem3__0 [25]),
        .I1(\alu0/div/dso_0 [25]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_3__0
       (.I0(\alu1/div/rem3__0 [25]),
        .I1(\alu1/div/dso_0 [25]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__5_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_4
       (.I0(\alu0/div/rem3__0 [24]),
        .I1(\alu0/div/dso_0 [24]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_4__0
       (.I0(\alu1/div/rem3__0 [24]),
        .I1(\alu1/div/dso_0 [24]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__5_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_1
       (.I0(\alu0/div/rem3__0 [31]),
        .I1(\alu0/div/rem3 ),
        .I2(\alu0/div/dso_0 [31]),
        .O(rem2_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_1__0
       (.I0(\alu1/div/rem3__0 [31]),
        .I1(\alu1/div/rem3 ),
        .I2(\alu1/div/dso_0 [31]),
        .O(rem2_carry__6_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_2
       (.I0(\alu0/div/rem3__0 [30]),
        .I1(\alu0/div/dso_0 [30]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_2__0
       (.I0(\alu1/div/rem3__0 [30]),
        .I1(\alu1/div/dso_0 [30]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__6_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_3
       (.I0(\alu0/div/rem3__0 [29]),
        .I1(\alu0/div/dso_0 [29]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_3__0
       (.I0(\alu1/div/rem3__0 [29]),
        .I1(\alu1/div/dso_0 [29]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__6_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_4
       (.I0(\alu0/div/rem3__0 [28]),
        .I1(\alu0/div/dso_0 [28]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry__6_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_4__0
       (.I0(\alu1/div/rem3__0 [28]),
        .I1(\alu1/div/dso_0 [28]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry__6_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem2_carry__7_i_1
       (.I0(\alu0/div/rem3 ),
        .I1(\alu0/div/rem3__0 [32]),
        .O(rem2_carry__7_i_1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem2_carry__7_i_1__0
       (.I0(\alu1/div/rem3 ),
        .I1(\alu1/div/rem3__0 [32]),
        .O(rem2_carry__7_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem2_carry_i_1
       (.I0(\alu0/div/rem3 ),
        .O(\alu0/div/fdiv/p_1_in3_in ));
  LUT1 #(
    .INIT(2'h1)) 
    rem2_carry_i_1__0
       (.I0(\alu1/div/rem3 ),
        .O(\alu1/div/fdiv/p_1_in3_in ));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_2
       (.I0(\alu0/div/rem3__0 [3]),
        .I1(\alu0/div/dso_0 [3]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_2__0
       (.I0(\alu1/div/rem3__0 [3]),
        .I1(\alu1/div/dso_0 [3]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_3
       (.I0(\alu0/div/rem3__0 [2]),
        .I1(\alu0/div/dso_0 [2]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_3__0
       (.I0(\alu1/div/rem3__0 [2]),
        .I1(\alu1/div/dso_0 [2]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_4
       (.I0(\alu0/div/rem3__0 [1]),
        .I1(\alu0/div/dso_0 [1]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_4__0
       (.I0(\alu1/div/rem3__0 [1]),
        .I1(\alu1/div/dso_0 [1]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_5
       (.I0(\alu0/div/den [30]),
        .I1(\alu0/div/dso_0 [0]),
        .I2(\alu0/div/rem3 ),
        .O(rem2_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_5__0
       (.I0(\alu1/div/den [30]),
        .I1(\alu1/div/dso_0 [0]),
        .I2(\alu1/div/rem3 ),
        .O(rem2_carry_i_5__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_1
       (.I0(\alu0/div/den [38]),
        .I1(\alu0/div/dso_0 [7]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_1__0
       (.I0(\alu1/div/den [38]),
        .I1(\alu1/div/dso_0 [7]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__0_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_2
       (.I0(\alu0/div/den [37]),
        .I1(\alu0/div/dso_0 [6]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_2__0
       (.I0(\alu1/div/den [37]),
        .I1(\alu1/div/dso_0 [6]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__0_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_3
       (.I0(\alu0/div/den [36]),
        .I1(\alu0/div/dso_0 [5]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_3__0
       (.I0(\alu1/div/den [36]),
        .I1(\alu1/div/dso_0 [5]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__0_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_4
       (.I0(\alu0/div/den [35]),
        .I1(\alu0/div/dso_0 [4]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__0_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_4__0
       (.I0(\alu1/div/den [35]),
        .I1(\alu1/div/dso_0 [4]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__0_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_1
       (.I0(\alu0/div/den [42]),
        .I1(\alu0/div/dso_0 [11]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_1__0
       (.I0(\alu1/div/den [42]),
        .I1(\alu1/div/dso_0 [11]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__1_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_2
       (.I0(\alu0/div/den [41]),
        .I1(\alu0/div/dso_0 [10]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_2__0
       (.I0(\alu1/div/den [41]),
        .I1(\alu1/div/dso_0 [10]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__1_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_3
       (.I0(\alu0/div/den [40]),
        .I1(\alu0/div/dso_0 [9]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_3__0
       (.I0(\alu1/div/den [40]),
        .I1(\alu1/div/dso_0 [9]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__1_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_4
       (.I0(\alu0/div/den [39]),
        .I1(\alu0/div/dso_0 [8]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__1_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_4__0
       (.I0(\alu1/div/den [39]),
        .I1(\alu1/div/dso_0 [8]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__1_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_1
       (.I0(\alu0/div/den [46]),
        .I1(\alu0/div/den [64]),
        .I2(\alu0/div/dso_0 [15]),
        .O(rem3_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_1__0
       (.I0(\alu1/div/den [46]),
        .I1(\alu1/div/den [64]),
        .I2(\alu1/div/dso_0 [15]),
        .O(rem3_carry__2_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_2
       (.I0(\alu0/div/den [45]),
        .I1(\alu0/div/dso_0 [14]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_2__0
       (.I0(\alu1/div/den [45]),
        .I1(\alu1/div/dso_0 [14]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__2_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_3
       (.I0(\alu0/div/den [44]),
        .I1(\alu0/div/dso_0 [13]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_3__0
       (.I0(\alu1/div/den [44]),
        .I1(\alu1/div/dso_0 [13]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__2_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_4
       (.I0(\alu0/div/den [43]),
        .I1(\alu0/div/dso_0 [12]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__2_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_4__0
       (.I0(\alu1/div/den [43]),
        .I1(\alu1/div/dso_0 [12]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__2_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_1
       (.I0(\alu0/div/den [50]),
        .I1(\alu0/div/dso_0 [19]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_1__0
       (.I0(\alu1/div/den [50]),
        .I1(\alu1/div/dso_0 [19]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__3_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_2
       (.I0(\alu0/div/den [49]),
        .I1(\alu0/div/dso_0 [18]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_2__0
       (.I0(\alu1/div/den [49]),
        .I1(\alu1/div/dso_0 [18]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__3_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_3
       (.I0(\alu0/div/den [48]),
        .I1(\alu0/div/dso_0 [17]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_3__0
       (.I0(\alu1/div/den [48]),
        .I1(\alu1/div/dso_0 [17]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__3_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_4
       (.I0(\alu0/div/den [47]),
        .I1(\alu0/div/dso_0 [16]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__3_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_4__0
       (.I0(\alu1/div/den [47]),
        .I1(\alu1/div/dso_0 [16]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__3_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_1
       (.I0(\alu0/div/den [54]),
        .I1(\alu0/div/dso_0 [23]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_1__0
       (.I0(\alu1/div/den [54]),
        .I1(\alu1/div/dso_0 [23]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__4_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_2
       (.I0(\alu0/div/den [53]),
        .I1(\alu0/div/dso_0 [22]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_2__0
       (.I0(\alu1/div/den [53]),
        .I1(\alu1/div/dso_0 [22]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__4_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_3
       (.I0(\alu0/div/den [52]),
        .I1(\alu0/div/dso_0 [21]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_3__0
       (.I0(\alu1/div/den [52]),
        .I1(\alu1/div/dso_0 [21]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__4_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_4
       (.I0(\alu0/div/den [51]),
        .I1(\alu0/div/dso_0 [20]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__4_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_4__0
       (.I0(\alu1/div/den [51]),
        .I1(\alu1/div/dso_0 [20]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__4_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_1
       (.I0(\alu0/div/den [58]),
        .I1(\alu0/div/dso_0 [27]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_1__0
       (.I0(\alu1/div/den [58]),
        .I1(\alu1/div/dso_0 [27]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__5_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_2
       (.I0(\alu0/div/den [57]),
        .I1(\alu0/div/dso_0 [26]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_2__0
       (.I0(\alu1/div/den [57]),
        .I1(\alu1/div/dso_0 [26]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__5_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_3
       (.I0(\alu0/div/den [56]),
        .I1(\alu0/div/dso_0 [25]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_3__0
       (.I0(\alu1/div/den [56]),
        .I1(\alu1/div/dso_0 [25]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__5_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_4
       (.I0(\alu0/div/den [55]),
        .I1(\alu0/div/dso_0 [24]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__5_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_4__0
       (.I0(\alu1/div/den [55]),
        .I1(\alu1/div/dso_0 [24]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__5_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_1
       (.I0(\alu0/div/den [62]),
        .I1(\alu0/div/den [64]),
        .I2(\alu0/div/dso_0 [31]),
        .O(rem3_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_1__0
       (.I0(\alu1/div/den [62]),
        .I1(\alu1/div/den [64]),
        .I2(\alu1/div/dso_0 [31]),
        .O(rem3_carry__6_i_1__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_2
       (.I0(\alu0/div/den [61]),
        .I1(\alu0/div/dso_0 [30]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_2__0
       (.I0(\alu1/div/den [61]),
        .I1(\alu1/div/dso_0 [30]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__6_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_3
       (.I0(\alu0/div/den [60]),
        .I1(\alu0/div/dso_0 [29]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_3__0
       (.I0(\alu1/div/den [60]),
        .I1(\alu1/div/dso_0 [29]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__6_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_4
       (.I0(\alu0/div/den [59]),
        .I1(\alu0/div/dso_0 [28]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry__6_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_4__0
       (.I0(\alu1/div/den [59]),
        .I1(\alu1/div/dso_0 [28]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry__6_i_4__0_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem3_carry__7_i_1
       (.I0(\alu0/div/den [63]),
        .I1(\alu0/div/den [64]),
        .O(rem3_carry__7_i_1_n_0));
  LUT2 #(
    .INIT(4'h9)) 
    rem3_carry__7_i_1__0
       (.I0(\alu1/div/den [63]),
        .I1(\alu1/div/den [64]),
        .O(rem3_carry__7_i_1__0_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem3_carry_i_1
       (.I0(\alu0/div/den [64]),
        .O(\alu0/div/fdiv/p_1_in5_in ));
  LUT1 #(
    .INIT(2'h1)) 
    rem3_carry_i_1__0
       (.I0(\alu1/div/den [64]),
        .O(\alu1/div/fdiv/p_1_in5_in ));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_2
       (.I0(\alu0/div/den [34]),
        .I1(\alu0/div/dso_0 [3]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_2__0
       (.I0(\alu1/div/den [34]),
        .I1(\alu1/div/dso_0 [3]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry_i_2__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_3
       (.I0(\alu0/div/den [33]),
        .I1(\alu0/div/dso_0 [2]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_3__0
       (.I0(\alu1/div/den [33]),
        .I1(\alu1/div/dso_0 [2]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry_i_3__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_4
       (.I0(\alu0/div/den [32]),
        .I1(\alu0/div/dso_0 [1]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry_i_4_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_4__0
       (.I0(\alu1/div/den [32]),
        .I1(\alu1/div/dso_0 [1]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry_i_4__0_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_5
       (.I0(\alu0/div/den2 ),
        .I1(\alu0/div/dso_0 [0]),
        .I2(\alu0/div/den [64]),
        .O(rem3_carry_i_5_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_5__0
       (.I0(\alu1/div/den2 ),
        .I1(\alu1/div/dso_0 [0]),
        .I2(\alu1/div/den [64]),
        .O(rem3_carry_i_5__0_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_2 
       (.I0(\alu0/div/p_0_out [11]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_2__0 
       (.I0(\alu1/div/p_0_out [11]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_3 
       (.I0(\alu0/div/p_0_out [10]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_3__0 
       (.I0(\alu1/div/p_0_out [10]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_4 
       (.I0(\alu0/div/p_0_out [9]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_4__0 
       (.I0(\alu1/div/p_0_out [9]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_5 
       (.I0(\alu0/div/p_0_out [8]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_5__0 
       (.I0(\alu1/div/p_0_out [8]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[11]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [11]),
        .I3(\alu0/div/rem [11]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [11]),
        .O(\rem[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [11]),
        .I3(\alu1/div/rem [11]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [11]),
        .O(\rem[11]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [10]),
        .I3(\alu0/div/rem [10]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [10]),
        .O(\rem[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [10]),
        .I3(\alu1/div/rem [10]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [10]),
        .O(\rem[11]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [9]),
        .I3(\alu0/div/rem [9]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [9]),
        .O(\rem[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [9]),
        .I3(\alu1/div/rem [9]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [9]),
        .O(\rem[11]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [8]),
        .I3(\alu0/div/rem [8]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [8]),
        .O(\rem[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[11]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [8]),
        .I3(\alu1/div/rem [8]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [8]),
        .O(\rem[11]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_2 
       (.I0(\alu0/div/p_0_out [15]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_2__0 
       (.I0(\alu1/div/p_0_out [15]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_3 
       (.I0(\alu0/div/p_0_out [14]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_3__0 
       (.I0(\alu1/div/p_0_out [14]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_4 
       (.I0(\alu0/div/p_0_out [13]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_4__0 
       (.I0(\alu1/div/p_0_out [13]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_5 
       (.I0(\alu0/div/p_0_out [12]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_5__0 
       (.I0(\alu1/div/p_0_out [12]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[15]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [15]),
        .I3(\alu0/div/rem [15]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [15]),
        .O(\rem[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [15]),
        .I3(\alu1/div/rem [15]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [15]),
        .O(\rem[15]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [14]),
        .I3(\alu0/div/rem [14]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [14]),
        .O(\rem[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [14]),
        .I3(\alu1/div/rem [14]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [14]),
        .O(\rem[15]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [13]),
        .I3(\alu0/div/rem [13]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [13]),
        .O(\rem[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [13]),
        .I3(\alu1/div/rem [13]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [13]),
        .O(\rem[15]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [12]),
        .I3(\alu0/div/rem [12]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [12]),
        .O(\rem[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[15]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [12]),
        .I3(\alu1/div/rem [12]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [12]),
        .O(\rem[15]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_2 
       (.I0(\alu0/div/p_0_out [19]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_2__0 
       (.I0(\alu1/div/p_0_out [19]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_3 
       (.I0(\alu0/div/p_0_out [18]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_3__0 
       (.I0(\alu1/div/p_0_out [18]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_4 
       (.I0(\alu0/div/p_0_out [17]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_4__0 
       (.I0(\alu1/div/p_0_out [17]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_5 
       (.I0(\alu0/div/p_0_out [16]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_5__0 
       (.I0(\alu1/div/p_0_out [16]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[19]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [19]),
        .I3(\alu0/div/rem [19]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [19]),
        .O(\rem[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [19]),
        .I3(\alu1/div/rem [19]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [19]),
        .O(\rem[19]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [18]),
        .I3(\alu0/div/rem [18]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [18]),
        .O(\rem[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [18]),
        .I3(\alu1/div/rem [18]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [18]),
        .O(\rem[19]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [17]),
        .I3(\alu0/div/rem [17]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [17]),
        .O(\rem[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [17]),
        .I3(\alu1/div/rem [17]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [17]),
        .O(\rem[19]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [16]),
        .I3(\alu0/div/rem [16]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [16]),
        .O(\rem[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[19]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [16]),
        .I3(\alu1/div/rem [16]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [16]),
        .O(\rem[19]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_2 
       (.I0(\alu0/div/p_0_out [23]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_2__0 
       (.I0(\alu1/div/p_0_out [23]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_3 
       (.I0(\alu0/div/p_0_out [22]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_3__0 
       (.I0(\alu1/div/p_0_out [22]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_4 
       (.I0(\alu0/div/p_0_out [21]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_4__0 
       (.I0(\alu1/div/p_0_out [21]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_5 
       (.I0(\alu0/div/p_0_out [20]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_5__0 
       (.I0(\alu1/div/p_0_out [20]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[23]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [23]),
        .I3(\alu0/div/rem [23]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [23]),
        .O(\rem[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [23]),
        .I3(\alu1/div/rem [23]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [23]),
        .O(\rem[23]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [22]),
        .I3(\alu0/div/rem [22]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [22]),
        .O(\rem[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [22]),
        .I3(\alu1/div/rem [22]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [22]),
        .O(\rem[23]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [21]),
        .I3(\alu0/div/rem [21]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [21]),
        .O(\rem[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [21]),
        .I3(\alu1/div/rem [21]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [21]),
        .O(\rem[23]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [20]),
        .I3(\alu0/div/rem [20]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [20]),
        .O(\rem[23]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[23]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [20]),
        .I3(\alu1/div/rem [20]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [20]),
        .O(\rem[23]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_2 
       (.I0(\alu0/div/p_0_out [27]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_2__0 
       (.I0(\alu1/div/p_0_out [27]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_3 
       (.I0(\alu0/div/p_0_out [26]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_3__0 
       (.I0(\alu1/div/p_0_out [26]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_4 
       (.I0(\alu0/div/p_0_out [25]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_4__0 
       (.I0(\alu1/div/p_0_out [25]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_5 
       (.I0(\alu0/div/p_0_out [24]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_5__0 
       (.I0(\alu1/div/p_0_out [24]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[27]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [27]),
        .I3(\alu0/div/rem [27]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [27]),
        .O(\rem[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [27]),
        .I3(\alu1/div/rem [27]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [27]),
        .O(\rem[27]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [26]),
        .I3(\alu0/div/rem [26]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [26]),
        .O(\rem[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [26]),
        .I3(\alu1/div/rem [26]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [26]),
        .O(\rem[27]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [25]),
        .I3(\alu0/div/rem [25]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [25]),
        .O(\rem[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [25]),
        .I3(\alu1/div/rem [25]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [25]),
        .O(\rem[27]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [24]),
        .I3(\alu0/div/rem [24]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [24]),
        .O(\rem[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[27]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [24]),
        .I3(\alu1/div/rem [24]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [24]),
        .O(\rem[27]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h0D000000FFFFFFFF)) 
    \rem[31]_i_1 
       (.I0(\alu0/div/dctl_long ),
        .I1(\alu0/div/dctl_stat [2]),
        .I2(\alu0/div/dctl_stat [3]),
        .I3(\alu0/div/dctl_stat [0]),
        .I4(\alu0/div/dctl_stat [1]),
        .I5(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_10 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [28]),
        .I3(\alu0/div/rem [28]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [28]),
        .O(\rem[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_10__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [28]),
        .I3(\alu1/div/rem [28]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [28]),
        .O(\rem[31]_i_10__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_11 
       (.I0(\alu0/div/chg_rem_sgn ),
        .I1(\alu0/div/chg_quo_sgn ),
        .O(\rem[31]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_11__0 
       (.I0(\alu1/div/chg_rem_sgn ),
        .I1(\alu1/div/chg_quo_sgn ),
        .O(\rem[31]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'h0D000000FFFFFFFF)) 
    \rem[31]_i_1__0 
       (.I0(\alu1/div/dctl_long ),
        .I1(\alu1/div/dctl_stat [2]),
        .I2(\alu1/div/dctl_stat [3]),
        .I3(\alu1/div/dctl_stat [0]),
        .I4(\alu1/div/dctl_stat [1]),
        .I5(\rem[31]_i_3__0_n_0 ),
        .O(\rem[31]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hFD77FD77FD7FFF7F)) 
    \rem[31]_i_3 
       (.I0(\alu0/div/dctl_stat [3]),
        .I1(\alu0/div/dctl_stat [1]),
        .I2(\alu0/div/dctl_stat [0]),
        .I3(\alu0/div/dctl_stat [2]),
        .I4(\alu0/div/fdiv_rem_msb_f ),
        .I5(\rem[31]_i_11_n_0 ),
        .O(\rem[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFD77FD77FD7FFF7F)) 
    \rem[31]_i_3__0 
       (.I0(\alu1/div/dctl_stat [3]),
        .I1(\alu1/div/dctl_stat [1]),
        .I2(\alu1/div/dctl_stat [0]),
        .I3(\alu1/div/dctl_stat [2]),
        .I4(\alu1/div/fdiv_rem_msb_f ),
        .I5(\rem[31]_i_11__0_n_0 ),
        .O(\rem[31]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_4 
       (.I0(\alu0/div/p_0_out [30]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_4__0 
       (.I0(\alu1/div/p_0_out [30]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[31]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_5 
       (.I0(\alu0/div/p_0_out [29]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_5__0 
       (.I0(\alu1/div/p_0_out [29]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[31]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_6 
       (.I0(\alu0/div/p_0_out [28]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_6__0 
       (.I0(\alu1/div/p_0_out [28]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[31]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [31]),
        .I3(\alu0/div/rem [31]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [31]),
        .O(\rem[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [31]),
        .I3(\alu1/div/rem [31]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [31]),
        .O(\rem[31]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [30]),
        .I3(\alu0/div/rem [30]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [30]),
        .O(\rem[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [30]),
        .I3(\alu1/div/rem [30]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [30]),
        .O(\rem[31]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [29]),
        .I3(\alu0/div/rem [29]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [29]),
        .O(\rem[31]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[31]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [29]),
        .I3(\alu1/div/rem [29]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [29]),
        .O(\rem[31]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_2 
       (.I0(\alu0/div/p_0_out [3]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_2__0 
       (.I0(\alu1/div/p_0_out [3]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_3 
       (.I0(\alu0/div/p_0_out [2]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_3__0 
       (.I0(\alu1/div/p_0_out [2]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_4 
       (.I0(\alu0/div/p_0_out [1]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_4__0 
       (.I0(\alu1/div/p_0_out [1]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_5 
       (.I0(\alu0/div/p_0_out [0]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_5__0 
       (.I0(\alu1/div/p_0_out [0]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[3]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [3]),
        .I3(\alu0/div/rem [3]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [3]),
        .O(\rem[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [3]),
        .I3(\alu1/div/rem [3]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [3]),
        .O(\rem[3]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [2]),
        .I3(\alu0/div/rem [2]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [2]),
        .O(\rem[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [2]),
        .I3(\alu1/div/rem [2]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [2]),
        .O(\rem[3]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [1]),
        .I3(\alu0/div/rem [1]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [1]),
        .O(\rem[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[3]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [1]),
        .I3(\alu1/div/rem [1]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [1]),
        .O(\rem[3]_i_8__0_n_0 ));
  LUT5 #(
    .INIT(32'hFF590059)) 
    \rem[3]_i_9 
       (.I0(\alu0/div/p_0_out [0]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\alu0/div/rem [0]),
        .I3(\rem[31]_i_3_n_0 ),
        .I4(\alu0/div/fdiv_rem [0]),
        .O(\rem[3]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFF590059)) 
    \rem[3]_i_9__0 
       (.I0(\alu1/div/p_0_out [0]),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(\alu1/div/rem [0]),
        .I3(\rem[31]_i_3__0_n_0 ),
        .I4(\alu1/div/fdiv_rem [0]),
        .O(\rem[3]_i_9__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_2 
       (.I0(\alu0/div/p_0_out [7]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_2__0 
       (.I0(\alu1/div/p_0_out [7]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_3 
       (.I0(\alu0/div/p_0_out [6]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_3__0 
       (.I0(\alu1/div/p_0_out [6]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_3__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_4 
       (.I0(\alu0/div/p_0_out [5]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_4__0 
       (.I0(\alu1/div/p_0_out [5]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_4__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_5 
       (.I0(\alu0/div/p_0_out [4]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_5__0 
       (.I0(\alu1/div/p_0_out [4]),
        .I1(\rem[31]_i_3__0_n_0 ),
        .O(\rem[7]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_6 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [7]),
        .I3(\alu0/div/rem [7]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [7]),
        .O(\rem[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_6__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [7]),
        .I3(\alu1/div/rem [7]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [7]),
        .O(\rem[7]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_7 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [6]),
        .I3(\alu0/div/rem [6]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [6]),
        .O(\rem[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_7__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [6]),
        .I3(\alu1/div/rem [6]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [6]),
        .O(\rem[7]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_8 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [5]),
        .I3(\alu0/div/rem [5]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [5]),
        .O(\rem[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_8__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [5]),
        .I3(\alu1/div/rem [5]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [5]),
        .O(\rem[7]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_9 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\alu0/div/p_0_out [4]),
        .I3(\alu0/div/rem [4]),
        .I4(\dso[31]_i_4_n_0 ),
        .I5(\alu0/div/fdiv_rem [4]),
        .O(\rem[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hDEFCFCFC12303030)) 
    \rem[7]_i_9__0 
       (.I0(\dso[31]_i_3__0_n_0 ),
        .I1(\rem[31]_i_3__0_n_0 ),
        .I2(\alu1/div/p_0_out [4]),
        .I3(\alu1/div/rem [4]),
        .I4(\dso[31]_i_4__0_n_0 ),
        .I5(\alu1/div/fdiv_rem [4]),
        .O(\rem[7]_i_9__0_n_0 ));
  CARRY4 \rem_reg[11]_i_1 
       (.CI(\rem_reg[7]_i_1_n_0 ),
        .CO({\rem_reg[11]_i_1_n_0 ,\rem_reg[11]_i_1_n_1 ,\rem_reg[11]_i_1_n_2 ,\rem_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[11]_i_2_n_0 ,\rem[11]_i_3_n_0 ,\rem[11]_i_4_n_0 ,\rem[11]_i_5_n_0 }),
        .O({\rem_reg[11]_i_1_n_4 ,\rem_reg[11]_i_1_n_5 ,\rem_reg[11]_i_1_n_6 ,\rem_reg[11]_i_1_n_7 }),
        .S({\rem[11]_i_6_n_0 ,\rem[11]_i_7_n_0 ,\rem[11]_i_8_n_0 ,\rem[11]_i_9_n_0 }));
  CARRY4 \rem_reg[11]_i_1__0 
       (.CI(\rem_reg[7]_i_1__0_n_0 ),
        .CO({\rem_reg[11]_i_1__0_n_0 ,\rem_reg[11]_i_1__0_n_1 ,\rem_reg[11]_i_1__0_n_2 ,\rem_reg[11]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[11]_i_2__0_n_0 ,\rem[11]_i_3__0_n_0 ,\rem[11]_i_4__0_n_0 ,\rem[11]_i_5__0_n_0 }),
        .O({\rem_reg[11]_i_1__0_n_4 ,\rem_reg[11]_i_1__0_n_5 ,\rem_reg[11]_i_1__0_n_6 ,\rem_reg[11]_i_1__0_n_7 }),
        .S({\rem[11]_i_6__0_n_0 ,\rem[11]_i_7__0_n_0 ,\rem[11]_i_8__0_n_0 ,\rem[11]_i_9__0_n_0 }));
  CARRY4 \rem_reg[15]_i_1 
       (.CI(\rem_reg[11]_i_1_n_0 ),
        .CO({\rem_reg[15]_i_1_n_0 ,\rem_reg[15]_i_1_n_1 ,\rem_reg[15]_i_1_n_2 ,\rem_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[15]_i_2_n_0 ,\rem[15]_i_3_n_0 ,\rem[15]_i_4_n_0 ,\rem[15]_i_5_n_0 }),
        .O({\rem_reg[15]_i_1_n_4 ,\rem_reg[15]_i_1_n_5 ,\rem_reg[15]_i_1_n_6 ,\rem_reg[15]_i_1_n_7 }),
        .S({\rem[15]_i_6_n_0 ,\rem[15]_i_7_n_0 ,\rem[15]_i_8_n_0 ,\rem[15]_i_9_n_0 }));
  CARRY4 \rem_reg[15]_i_1__0 
       (.CI(\rem_reg[11]_i_1__0_n_0 ),
        .CO({\rem_reg[15]_i_1__0_n_0 ,\rem_reg[15]_i_1__0_n_1 ,\rem_reg[15]_i_1__0_n_2 ,\rem_reg[15]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[15]_i_2__0_n_0 ,\rem[15]_i_3__0_n_0 ,\rem[15]_i_4__0_n_0 ,\rem[15]_i_5__0_n_0 }),
        .O({\rem_reg[15]_i_1__0_n_4 ,\rem_reg[15]_i_1__0_n_5 ,\rem_reg[15]_i_1__0_n_6 ,\rem_reg[15]_i_1__0_n_7 }),
        .S({\rem[15]_i_6__0_n_0 ,\rem[15]_i_7__0_n_0 ,\rem[15]_i_8__0_n_0 ,\rem[15]_i_9__0_n_0 }));
  CARRY4 \rem_reg[19]_i_1 
       (.CI(\rem_reg[15]_i_1_n_0 ),
        .CO({\rem_reg[19]_i_1_n_0 ,\rem_reg[19]_i_1_n_1 ,\rem_reg[19]_i_1_n_2 ,\rem_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[19]_i_2_n_0 ,\rem[19]_i_3_n_0 ,\rem[19]_i_4_n_0 ,\rem[19]_i_5_n_0 }),
        .O({\rem_reg[19]_i_1_n_4 ,\rem_reg[19]_i_1_n_5 ,\rem_reg[19]_i_1_n_6 ,\rem_reg[19]_i_1_n_7 }),
        .S({\rem[19]_i_6_n_0 ,\rem[19]_i_7_n_0 ,\rem[19]_i_8_n_0 ,\rem[19]_i_9_n_0 }));
  CARRY4 \rem_reg[19]_i_1__0 
       (.CI(\rem_reg[15]_i_1__0_n_0 ),
        .CO({\rem_reg[19]_i_1__0_n_0 ,\rem_reg[19]_i_1__0_n_1 ,\rem_reg[19]_i_1__0_n_2 ,\rem_reg[19]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[19]_i_2__0_n_0 ,\rem[19]_i_3__0_n_0 ,\rem[19]_i_4__0_n_0 ,\rem[19]_i_5__0_n_0 }),
        .O({\rem_reg[19]_i_1__0_n_4 ,\rem_reg[19]_i_1__0_n_5 ,\rem_reg[19]_i_1__0_n_6 ,\rem_reg[19]_i_1__0_n_7 }),
        .S({\rem[19]_i_6__0_n_0 ,\rem[19]_i_7__0_n_0 ,\rem[19]_i_8__0_n_0 ,\rem[19]_i_9__0_n_0 }));
  CARRY4 \rem_reg[23]_i_1 
       (.CI(\rem_reg[19]_i_1_n_0 ),
        .CO({\rem_reg[23]_i_1_n_0 ,\rem_reg[23]_i_1_n_1 ,\rem_reg[23]_i_1_n_2 ,\rem_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[23]_i_2_n_0 ,\rem[23]_i_3_n_0 ,\rem[23]_i_4_n_0 ,\rem[23]_i_5_n_0 }),
        .O({\rem_reg[23]_i_1_n_4 ,\rem_reg[23]_i_1_n_5 ,\rem_reg[23]_i_1_n_6 ,\rem_reg[23]_i_1_n_7 }),
        .S({\rem[23]_i_6_n_0 ,\rem[23]_i_7_n_0 ,\rem[23]_i_8_n_0 ,\rem[23]_i_9_n_0 }));
  CARRY4 \rem_reg[23]_i_1__0 
       (.CI(\rem_reg[19]_i_1__0_n_0 ),
        .CO({\rem_reg[23]_i_1__0_n_0 ,\rem_reg[23]_i_1__0_n_1 ,\rem_reg[23]_i_1__0_n_2 ,\rem_reg[23]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[23]_i_2__0_n_0 ,\rem[23]_i_3__0_n_0 ,\rem[23]_i_4__0_n_0 ,\rem[23]_i_5__0_n_0 }),
        .O({\rem_reg[23]_i_1__0_n_4 ,\rem_reg[23]_i_1__0_n_5 ,\rem_reg[23]_i_1__0_n_6 ,\rem_reg[23]_i_1__0_n_7 }),
        .S({\rem[23]_i_6__0_n_0 ,\rem[23]_i_7__0_n_0 ,\rem[23]_i_8__0_n_0 ,\rem[23]_i_9__0_n_0 }));
  CARRY4 \rem_reg[27]_i_1 
       (.CI(\rem_reg[23]_i_1_n_0 ),
        .CO({\rem_reg[27]_i_1_n_0 ,\rem_reg[27]_i_1_n_1 ,\rem_reg[27]_i_1_n_2 ,\rem_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[27]_i_2_n_0 ,\rem[27]_i_3_n_0 ,\rem[27]_i_4_n_0 ,\rem[27]_i_5_n_0 }),
        .O({\rem_reg[27]_i_1_n_4 ,\rem_reg[27]_i_1_n_5 ,\rem_reg[27]_i_1_n_6 ,\rem_reg[27]_i_1_n_7 }),
        .S({\rem[27]_i_6_n_0 ,\rem[27]_i_7_n_0 ,\rem[27]_i_8_n_0 ,\rem[27]_i_9_n_0 }));
  CARRY4 \rem_reg[27]_i_1__0 
       (.CI(\rem_reg[23]_i_1__0_n_0 ),
        .CO({\rem_reg[27]_i_1__0_n_0 ,\rem_reg[27]_i_1__0_n_1 ,\rem_reg[27]_i_1__0_n_2 ,\rem_reg[27]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[27]_i_2__0_n_0 ,\rem[27]_i_3__0_n_0 ,\rem[27]_i_4__0_n_0 ,\rem[27]_i_5__0_n_0 }),
        .O({\rem_reg[27]_i_1__0_n_4 ,\rem_reg[27]_i_1__0_n_5 ,\rem_reg[27]_i_1__0_n_6 ,\rem_reg[27]_i_1__0_n_7 }),
        .S({\rem[27]_i_6__0_n_0 ,\rem[27]_i_7__0_n_0 ,\rem[27]_i_8__0_n_0 ,\rem[27]_i_9__0_n_0 }));
  CARRY4 \rem_reg[31]_i_2 
       (.CI(\rem_reg[27]_i_1_n_0 ),
        .CO({\rem_reg[31]_i_2_n_1 ,\rem_reg[31]_i_2_n_2 ,\rem_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rem[31]_i_4_n_0 ,\rem[31]_i_5_n_0 ,\rem[31]_i_6_n_0 }),
        .O({\rem_reg[31]_i_2_n_4 ,\rem_reg[31]_i_2_n_5 ,\rem_reg[31]_i_2_n_6 ,\rem_reg[31]_i_2_n_7 }),
        .S({\rem[31]_i_7_n_0 ,\rem[31]_i_8_n_0 ,\rem[31]_i_9_n_0 ,\rem[31]_i_10_n_0 }));
  CARRY4 \rem_reg[31]_i_2__0 
       (.CI(\rem_reg[27]_i_1__0_n_0 ),
        .CO({\rem_reg[31]_i_2__0_n_1 ,\rem_reg[31]_i_2__0_n_2 ,\rem_reg[31]_i_2__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rem[31]_i_4__0_n_0 ,\rem[31]_i_5__0_n_0 ,\rem[31]_i_6__0_n_0 }),
        .O({\rem_reg[31]_i_2__0_n_4 ,\rem_reg[31]_i_2__0_n_5 ,\rem_reg[31]_i_2__0_n_6 ,\rem_reg[31]_i_2__0_n_7 }),
        .S({\rem[31]_i_7__0_n_0 ,\rem[31]_i_8__0_n_0 ,\rem[31]_i_9__0_n_0 ,\rem[31]_i_10__0_n_0 }));
  CARRY4 \rem_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\rem_reg[3]_i_1_n_0 ,\rem_reg[3]_i_1_n_1 ,\rem_reg[3]_i_1_n_2 ,\rem_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[3]_i_2_n_0 ,\rem[3]_i_3_n_0 ,\rem[3]_i_4_n_0 ,\rem[3]_i_5_n_0 }),
        .O({\rem_reg[3]_i_1_n_4 ,\rem_reg[3]_i_1_n_5 ,\rem_reg[3]_i_1_n_6 ,\rem_reg[3]_i_1_n_7 }),
        .S({\rem[3]_i_6_n_0 ,\rem[3]_i_7_n_0 ,\rem[3]_i_8_n_0 ,\rem[3]_i_9_n_0 }));
  CARRY4 \rem_reg[3]_i_1__0 
       (.CI(\<const0> ),
        .CO({\rem_reg[3]_i_1__0_n_0 ,\rem_reg[3]_i_1__0_n_1 ,\rem_reg[3]_i_1__0_n_2 ,\rem_reg[3]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[3]_i_2__0_n_0 ,\rem[3]_i_3__0_n_0 ,\rem[3]_i_4__0_n_0 ,\rem[3]_i_5__0_n_0 }),
        .O({\rem_reg[3]_i_1__0_n_4 ,\rem_reg[3]_i_1__0_n_5 ,\rem_reg[3]_i_1__0_n_6 ,\rem_reg[3]_i_1__0_n_7 }),
        .S({\rem[3]_i_6__0_n_0 ,\rem[3]_i_7__0_n_0 ,\rem[3]_i_8__0_n_0 ,\rem[3]_i_9__0_n_0 }));
  CARRY4 \rem_reg[7]_i_1 
       (.CI(\rem_reg[3]_i_1_n_0 ),
        .CO({\rem_reg[7]_i_1_n_0 ,\rem_reg[7]_i_1_n_1 ,\rem_reg[7]_i_1_n_2 ,\rem_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[7]_i_2_n_0 ,\rem[7]_i_3_n_0 ,\rem[7]_i_4_n_0 ,\rem[7]_i_5_n_0 }),
        .O({\rem_reg[7]_i_1_n_4 ,\rem_reg[7]_i_1_n_5 ,\rem_reg[7]_i_1_n_6 ,\rem_reg[7]_i_1_n_7 }),
        .S({\rem[7]_i_6_n_0 ,\rem[7]_i_7_n_0 ,\rem[7]_i_8_n_0 ,\rem[7]_i_9_n_0 }));
  CARRY4 \rem_reg[7]_i_1__0 
       (.CI(\rem_reg[3]_i_1__0_n_0 ),
        .CO({\rem_reg[7]_i_1__0_n_0 ,\rem_reg[7]_i_1__0_n_1 ,\rem_reg[7]_i_1__0_n_2 ,\rem_reg[7]_i_1__0_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[7]_i_2__0_n_0 ,\rem[7]_i_3__0_n_0 ,\rem[7]_i_4__0_n_0 ,\rem[7]_i_5__0_n_0 }),
        .O({\rem_reg[7]_i_1__0_n_4 ,\rem_reg[7]_i_1__0_n_5 ,\rem_reg[7]_i_1__0_n_6 ,\rem_reg[7]_i_1__0_n_7 }),
        .S({\rem[7]_i_6__0_n_0 ,\rem[7]_i_7__0_n_0 ,\rem[7]_i_8__0_n_0 ,\rem[7]_i_9__0_n_0 }));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[0]_i_1 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/add_out [0]),
        .I3(\remden[64]_i_1_n_0 ),
        .I4(a0bus_0[0]),
        .O(\remden[0]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[0]_i_1__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/add_out [0]),
        .I3(\remden[64]_i_1__0_n_0 ),
        .I4(a1bus_0[0]),
        .O(\remden[0]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[10]_i_1 
       (.I0(\alu0/div/add_out [10]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [6]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[10]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[10]_i_1__0 
       (.I0(\alu1/div/add_out [10]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[10]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [6]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[10]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[11]_i_1 
       (.I0(\alu0/div/add_out [11]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [7]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[11]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[11]_i_1__0 
       (.I0(\alu1/div/add_out [11]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[11]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [7]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[11]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[12]_i_1 
       (.I0(\alu0/div/add_out [12]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [8]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[12]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[12]_i_1__0 
       (.I0(\alu1/div/add_out [12]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[12]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [8]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[12]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[13]_i_1 
       (.I0(\alu0/div/add_out [13]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[13]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [9]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[13]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[13]_i_1__0 
       (.I0(\alu1/div/add_out [13]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[13]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [9]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[13]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[14]_i_1 
       (.I0(\alu0/div/add_out [14]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[14]),
        .I4(\alu0/div/den [10]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[14]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[14]_i_1__0 
       (.I0(\alu1/div/add_out [14]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[14]),
        .I4(\alu1/div/den [10]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[14]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[15]_i_1 
       (.I0(\alu0/div/add_out [15]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [11]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[15]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[15]_i_1__0 
       (.I0(\alu1/div/add_out [15]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [11]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[15]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[16]_i_1 
       (.I0(\alu0/div/add_out [16]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[16]_i_2_n_0 ),
        .O(\remden[16]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[16]_i_1__0 
       (.I0(\alu1/div/add_out [16]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[16]_i_2__0_n_0 ),
        .O(\remden[16]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[16]_i_2 
       (.I0(a0bus_0[16]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[0]),
        .I4(\alu0/div/den [12]),
        .O(\remden[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[16]_i_2__0 
       (.I0(a1bus_0[16]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[0]),
        .I4(\alu1/div/den [12]),
        .O(\remden[16]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[17]_i_1 
       (.I0(\alu0/div/add_out [17]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[17]_i_2_n_0 ),
        .O(\remden[17]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[17]_i_1__0 
       (.I0(\alu1/div/add_out [17]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[17]_i_2__0_n_0 ),
        .O(\remden[17]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[17]_i_2 
       (.I0(a0bus_0[17]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[1]),
        .I4(\alu0/div/den [13]),
        .O(\remden[17]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[17]_i_2__0 
       (.I0(a1bus_0[17]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[1]),
        .I4(\alu1/div/den [13]),
        .O(\remden[17]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[18]_i_1 
       (.I0(\alu0/div/add_out [18]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[18]_i_2_n_0 ),
        .O(\remden[18]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[18]_i_1__0 
       (.I0(\alu1/div/add_out [18]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[18]_i_2__0_n_0 ),
        .O(\remden[18]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[18]_i_2 
       (.I0(a0bus_0[18]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[2]),
        .I4(\alu0/div/den [14]),
        .O(\remden[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[18]_i_2__0 
       (.I0(a1bus_0[18]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[2]),
        .I4(\alu1/div/den [14]),
        .O(\remden[18]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[19]_i_1 
       (.I0(\alu0/div/add_out [19]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[19]_i_2_n_0 ),
        .O(\remden[19]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[19]_i_1__0 
       (.I0(\alu1/div/add_out [19]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[19]_i_2__0_n_0 ),
        .O(\remden[19]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[19]_i_2 
       (.I0(a0bus_0[19]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[3]),
        .I4(\alu0/div/den [15]),
        .O(\remden[19]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[19]_i_2__0 
       (.I0(a1bus_0[19]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[3]),
        .I4(\alu1/div/den [15]),
        .O(\remden[19]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[1]_i_1 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/add_out [1]),
        .I3(\remden[64]_i_1_n_0 ),
        .I4(a0bus_0[1]),
        .O(\remden[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[1]_i_1__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/add_out [1]),
        .I3(\remden[64]_i_1__0_n_0 ),
        .I4(a1bus_0[1]),
        .O(\remden[1]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[20]_i_1 
       (.I0(\alu0/div/add_out [20]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[20]_i_2_n_0 ),
        .O(\remden[20]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[20]_i_1__0 
       (.I0(\alu1/div/add_out [20]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[20]_i_2__0_n_0 ),
        .O(\remden[20]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[20]_i_2 
       (.I0(a0bus_0[20]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[4]),
        .I4(\alu0/div/den [16]),
        .O(\remden[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[20]_i_2__0 
       (.I0(a1bus_0[20]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[4]),
        .I4(\alu1/div/den [16]),
        .O(\remden[20]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[21]_i_1 
       (.I0(\alu0/div/add_out [21]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[21]_i_2_n_0 ),
        .O(\remden[21]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[21]_i_1__0 
       (.I0(\alu1/div/add_out [21]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[21]_i_2__0_n_0 ),
        .O(\remden[21]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[21]_i_2 
       (.I0(\alu0/div/den [17]),
        .I1(\alu0/mul_a_i [21]),
        .I2(\dso[31]_i_5_n_0 ),
        .I3(a0bus_0[5]),
        .I4(\rgf/sreg/sr [8]),
        .O(\remden[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[21]_i_2__0 
       (.I0(\alu1/div/den [17]),
        .I1(\alu1/mul_a_i [21]),
        .I2(\dso[31]_i_5__0_n_0 ),
        .I3(a1bus_0[5]),
        .I4(\rgf/sreg/sr [8]),
        .O(\remden[21]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[22]_i_1 
       (.I0(\alu0/div/add_out [22]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[22]_i_2_n_0 ),
        .O(\remden[22]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[22]_i_1__0 
       (.I0(\alu1/div/add_out [22]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[22]_i_2__0_n_0 ),
        .O(\remden[22]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[22]_i_2 
       (.I0(a0bus_0[22]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[6]),
        .I4(\alu0/div/den [18]),
        .O(\remden[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[22]_i_2__0 
       (.I0(a1bus_0[22]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[6]),
        .I4(\alu1/div/den [18]),
        .O(\remden[22]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[23]_i_1 
       (.I0(\alu0/div/add_out [23]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[23]_i_2_n_0 ),
        .O(\remden[23]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[23]_i_1__0 
       (.I0(\alu1/div/add_out [23]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[23]_i_2__0_n_0 ),
        .O(\remden[23]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[23]_i_2 
       (.I0(a0bus_0[23]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[7]),
        .I4(\alu0/div/den [19]),
        .O(\remden[23]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[23]_i_2__0 
       (.I0(a1bus_0[23]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[7]),
        .I4(\alu1/div/den [19]),
        .O(\remden[23]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[24]_i_1 
       (.I0(\alu0/div/add_out [24]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[24]_i_2_n_0 ),
        .O(\remden[24]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[24]_i_1__0 
       (.I0(\alu1/div/add_out [24]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[24]_i_2__0_n_0 ),
        .O(\remden[24]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[24]_i_2 
       (.I0(a0bus_0[24]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[8]),
        .I4(\alu0/div/den [20]),
        .O(\remden[24]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[24]_i_2__0 
       (.I0(a1bus_0[24]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[8]),
        .I4(\alu1/div/den [20]),
        .O(\remden[24]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[25]_i_1 
       (.I0(\alu0/div/add_out [25]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[25]_i_2_n_0 ),
        .O(\remden[25]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[25]_i_1__0 
       (.I0(\alu1/div/add_out [25]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[25]_i_2__0_n_0 ),
        .O(\remden[25]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[25]_i_2 
       (.I0(a0bus_0[25]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[9]),
        .I4(\alu0/div/den [21]),
        .O(\remden[25]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[25]_i_2__0 
       (.I0(a1bus_0[25]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[9]),
        .I4(\alu1/div/den [21]),
        .O(\remden[25]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[26]_i_1 
       (.I0(\alu0/div/add_out [26]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[26]_i_2_n_0 ),
        .O(\remden[26]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[26]_i_1__0 
       (.I0(\alu1/div/add_out [26]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[26]_i_2__0_n_0 ),
        .O(\remden[26]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[26]_i_2 
       (.I0(\alu0/div/den [22]),
        .I1(\alu0/mul_a_i [26]),
        .I2(\dso[31]_i_5_n_0 ),
        .I3(a0bus_0[10]),
        .I4(\rgf/sreg/sr [8]),
        .O(\remden[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hCACAFACA)) 
    \remden[26]_i_2__0 
       (.I0(\alu1/div/den [22]),
        .I1(\alu1/mul_a_i [26]),
        .I2(\dso[31]_i_5__0_n_0 ),
        .I3(a1bus_0[10]),
        .I4(\rgf/sreg/sr [8]),
        .O(\remden[26]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[27]_i_1 
       (.I0(\alu0/div/add_out [27]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[27]_i_2_n_0 ),
        .O(\remden[27]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[27]_i_1__0 
       (.I0(\alu1/div/add_out [27]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[27]_i_2__0_n_0 ),
        .O(\remden[27]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[27]_i_2 
       (.I0(a0bus_0[27]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[11]),
        .I4(\alu0/div/den [23]),
        .O(\remden[27]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[27]_i_2__0 
       (.I0(a1bus_0[27]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[11]),
        .I4(\alu1/div/den [23]),
        .O(\remden[27]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[28]_i_1 
       (.I0(\alu0/div/add_out [28]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[28]_i_2_n_0 ),
        .O(\remden[28]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[28]_i_1__0 
       (.I0(\alu1/div/add_out [28]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[28]_i_2__0_n_0 ),
        .O(\remden[28]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[28]_i_2 
       (.I0(a0bus_0[28]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[12]),
        .I4(\alu0/div/den [24]),
        .O(\remden[28]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[28]_i_2__0 
       (.I0(a1bus_0[28]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[12]),
        .I4(\alu1/div/den [24]),
        .O(\remden[28]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[29]_i_1 
       (.I0(\alu0/div/add_out [29]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[29]_i_2_n_0 ),
        .O(\remden[29]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[29]_i_1__0 
       (.I0(\alu1/div/add_out [29]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[29]_i_2__0_n_0 ),
        .O(\remden[29]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[29]_i_2 
       (.I0(a0bus_0[29]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[13]),
        .I4(\alu0/div/den [25]),
        .O(\remden[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[29]_i_2__0 
       (.I0(a1bus_0[29]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[13]),
        .I4(\alu1/div/den [25]),
        .O(\remden[29]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[2]_i_1 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/add_out [2]),
        .I3(\remden[64]_i_1_n_0 ),
        .I4(a0bus_0[2]),
        .O(\remden[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[2]_i_1__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/add_out [2]),
        .I3(\remden[64]_i_1__0_n_0 ),
        .I4(a1bus_0[2]),
        .O(\remden[2]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[30]_i_1 
       (.I0(\alu0/div/add_out [30]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\remden[30]_i_2_n_0 ),
        .O(\remden[30]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \remden[30]_i_1__0 
       (.I0(\alu1/div/add_out [30]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\remden[30]_i_2__0_n_0 ),
        .O(\remden[30]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[30]_i_2 
       (.I0(a0bus_0[30]),
        .I1(\dso[31]_i_5_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[14]),
        .I4(\alu0/div/den [26]),
        .O(\remden[30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[30]_i_2__0 
       (.I0(a1bus_0[30]),
        .I1(\dso[31]_i_5__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[14]),
        .I4(\alu1/div/den [26]),
        .O(\remden[30]_i_2__0_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFF1)) 
    \remden[31]_i_1 
       (.I0(\remden[64]_i_4_n_0 ),
        .I1(\alu0/div/dctl_stat [1]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[64]_i_1_n_0 ),
        .I4(rst_n),
        .O(\remden[31]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFF1)) 
    \remden[31]_i_1__0 
       (.I0(\remden[64]_i_4__0_n_0 ),
        .I1(\alu1/div/dctl_stat [1]),
        .I2(\remden[64]_i_5__0_n_0 ),
        .I3(\remden[64]_i_1__0_n_0 ),
        .I4(rst_n),
        .O(\remden[31]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hBB88B8B8)) 
    \remden[31]_i_2 
       (.I0(\alu0/div/add_out [31]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\alu0/div/den [27]),
        .I3(\remden[31]_i_3_n_0 ),
        .I4(\dso[31]_i_5_n_0 ),
        .O(\remden[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB88B8B8B8B8)) 
    \remden[31]_i_2__0 
       (.I0(\alu1/div/add_out [31]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\alu1/div/den [27]),
        .I3(\alu1/mul_a_i [31]),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[31]_i_2__0_n_0 ));
  LUT3 #(
    .INIT(8'hD8)) 
    \remden[31]_i_3 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(a0bus_0[15]),
        .O(\remden[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[32]_i_1 
       (.I0(\alu0/div/fdiv_rem [0]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[32]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[32]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [0]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[32]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[33]_i_1 
       (.I0(\alu0/div/fdiv_rem [1]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[33]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[33]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [1]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[33]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[34]_i_1 
       (.I0(\alu0/div/fdiv_rem [2]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[34]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[34]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [2]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[34]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[35]_i_1 
       (.I0(\alu0/div/fdiv_rem [3]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[35]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[35]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [3]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[35]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[36]_i_1 
       (.I0(\alu0/div/fdiv_rem [4]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[36]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[36]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [4]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[36]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[37]_i_1 
       (.I0(\alu0/div/fdiv_rem [5]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[37]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[37]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [5]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[37]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[38]_i_1 
       (.I0(\alu0/div/fdiv_rem [6]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[38]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[38]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [6]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[38]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[39]_i_1 
       (.I0(\alu0/div/fdiv_rem [7]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[39]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[39]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [7]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[39]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[3]_i_1 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu0/div/add_out [3]),
        .I3(\remden[64]_i_1_n_0 ),
        .I4(a0bus_0[3]),
        .O(\remden[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hF088F000)) 
    \remden[3]_i_1__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\alu1/div/add_out [3]),
        .I3(\remden[64]_i_1__0_n_0 ),
        .I4(a1bus_0[3]),
        .O(\remden[3]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[40]_i_1 
       (.I0(\alu0/div/fdiv_rem [8]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[40]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[40]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [8]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[40]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[41]_i_1 
       (.I0(\alu0/div/fdiv_rem [9]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[41]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[41]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [9]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[41]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[42]_i_1 
       (.I0(\alu0/div/fdiv_rem [10]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[42]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[42]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [10]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[42]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[43]_i_1 
       (.I0(\alu0/div/fdiv_rem [11]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[43]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[43]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [11]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[43]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[44]_i_1 
       (.I0(\alu0/div/fdiv_rem [12]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[44]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[44]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [12]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[44]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[45]_i_1 
       (.I0(\alu0/div/fdiv_rem [13]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[45]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[45]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [13]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[45]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[46]_i_1 
       (.I0(\alu0/div/fdiv_rem [14]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[46]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[46]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [14]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[46]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[47]_i_1 
       (.I0(\alu0/div/fdiv_rem [15]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[47]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[47]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [15]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[47]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[48]_i_1 
       (.I0(\alu0/div/fdiv_rem [16]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[48]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[48]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [16]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[48]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[49]_i_1 
       (.I0(\alu0/div/fdiv_rem [17]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[49]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[49]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [17]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[49]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[4]_i_1 
       (.I0(\alu0/div/add_out [4]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [0]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[4]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[4]_i_1__0 
       (.I0(\alu1/div/add_out [4]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[4]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [0]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[4]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[50]_i_1 
       (.I0(\alu0/div/fdiv_rem [18]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[50]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[50]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [18]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[50]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[51]_i_1 
       (.I0(\alu0/div/fdiv_rem [19]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[51]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[51]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [19]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[51]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[52]_i_1 
       (.I0(\alu0/div/fdiv_rem [20]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[52]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[52]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [20]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[52]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[53]_i_1 
       (.I0(\alu0/div/fdiv_rem [21]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[53]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[53]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [21]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[53]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[54]_i_1 
       (.I0(\alu0/div/fdiv_rem [22]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[54]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[54]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [22]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[54]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[55]_i_1 
       (.I0(\alu0/div/fdiv_rem [23]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[55]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[55]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [23]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[55]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[56]_i_1 
       (.I0(\alu0/div/fdiv_rem [24]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[56]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[56]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [24]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[56]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[57]_i_1 
       (.I0(\alu0/div/fdiv_rem [25]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[57]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[57]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [25]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[57]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[58]_i_1 
       (.I0(\alu0/div/fdiv_rem [26]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[58]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[58]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [26]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[58]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[59]_i_1 
       (.I0(\alu0/div/fdiv_rem [27]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[59]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[59]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [27]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[59]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[5]_i_1 
       (.I0(\alu0/div/add_out [5]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [1]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[5]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[5]_i_1__0 
       (.I0(\alu1/div/add_out [5]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[5]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [1]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[5]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[60]_i_1 
       (.I0(\alu0/div/fdiv_rem [28]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[60]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[60]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [28]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[60]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[61]_i_1 
       (.I0(\alu0/div/fdiv_rem [29]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[61]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[61]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [29]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[61]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[62]_i_1 
       (.I0(\alu0/div/fdiv_rem [30]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[62]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[62]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [30]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[62]_i_1__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[63]_i_1 
       (.I0(\alu0/div/fdiv_rem [31]),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[63]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[63]_i_1__0 
       (.I0(\alu1/div/fdiv_rem [31]),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[63]_i_1__0_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \remden[64]_i_1 
       (.I0(\dso[31]_i_4_n_0 ),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\rem[31]_i_3_n_0 ),
        .O(\remden[64]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \remden[64]_i_1__0 
       (.I0(\dso[31]_i_4__0_n_0 ),
        .I1(\dso[31]_i_3__0_n_0 ),
        .I2(\rem[31]_i_3__0_n_0 ),
        .O(\remden[64]_i_1__0_n_0 ));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \remden[64]_i_2 
       (.I0(\remden[64]_i_4_n_0 ),
        .I1(\alu0/div/dctl_stat [1]),
        .I2(\remden[64]_i_5_n_0 ),
        .I3(\remden[64]_i_1_n_0 ),
        .O(\remden[64]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \remden[64]_i_2__0 
       (.I0(\remden[64]_i_4__0_n_0 ),
        .I1(\alu1/div/dctl_stat [1]),
        .I2(\remden[64]_i_5__0_n_0 ),
        .I3(\remden[64]_i_1__0_n_0 ),
        .O(\remden[64]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[64]_i_3 
       (.I0(\alu0/div/p_0_in0 ),
        .I1(\remden[64]_i_6_n_0 ),
        .O(\remden[64]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[64]_i_3__0 
       (.I0(\alu1/div/p_0_in0 ),
        .I1(\remden[64]_i_6__0_n_0 ),
        .O(\remden[64]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hD5000055DD550055)) 
    \remden[64]_i_4 
       (.I0(\alu0/div/dctl_stat [0]),
        .I1(\alu0/div/dctl/dctl_sign ),
        .I2(\alu0/div/den2 ),
        .I3(\alu0/div/dctl_stat [2]),
        .I4(\alu0/div/dctl_stat [3]),
        .I5(chg_quo_sgn_i_2_n_0),
        .O(\remden[64]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hD5000055DD550055)) 
    \remden[64]_i_4__0 
       (.I0(\alu1/div/dctl_stat [0]),
        .I1(\alu1/div/dctl/dctl_sign ),
        .I2(\alu1/div/den2 ),
        .I3(\alu1/div/dctl_stat [2]),
        .I4(\alu1/div/dctl_stat [3]),
        .I5(chg_quo_sgn_i_2__0_n_0),
        .O(\remden[64]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAFEAABAAABA)) 
    \remden[64]_i_5 
       (.I0(\remden[64]_i_6_n_0 ),
        .I1(\alu0/div/dctl_stat [0]),
        .I2(\alu0/div/dctl_stat [1]),
        .I3(\alu0/div/dctl_stat [3]),
        .I4(\alu0/div/dctl_stat [2]),
        .I5(\alu0/div/dctl_long ),
        .O(\remden[64]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAFEAABAAABA)) 
    \remden[64]_i_5__0 
       (.I0(\remden[64]_i_6__0_n_0 ),
        .I1(\alu1/div/dctl_stat [0]),
        .I2(\alu1/div/dctl_stat [1]),
        .I3(\alu1/div/dctl_stat [3]),
        .I4(\alu1/div/dctl_stat [2]),
        .I5(\alu1/div/dctl_long ),
        .O(\remden[64]_i_5__0_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_6 
       (.I0(\dso[31]_i_5_n_0 ),
        .I1(rst_n),
        .O(\remden[64]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_6__0 
       (.I0(\dso[31]_i_5__0_n_0 ),
        .I1(rst_n),
        .O(\remden[64]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[6]_i_1 
       (.I0(\alu0/div/add_out [6]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [2]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[6]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[6]_i_1__0 
       (.I0(\alu1/div/add_out [6]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[6]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [2]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[6]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[7]_i_1 
       (.I0(\alu0/div/add_out [7]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [3]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[7]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[7]_i_1__0 
       (.I0(\alu1/div/add_out [7]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[7]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [3]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[7]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[8]_i_1 
       (.I0(\alu0/div/add_out [8]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu0/div/den [4]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[8]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[8]_i_1__0 
       (.I0(\alu1/div/add_out [8]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(a1bus_0[8]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/div/den [4]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[8]_i_1__0_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[9]_i_1 
       (.I0(\alu0/div/add_out [9]),
        .I1(\remden[64]_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a0bus_0[9]),
        .I4(\alu0/div/den [5]),
        .I5(\dso[31]_i_5_n_0 ),
        .O(\remden[9]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[9]_i_1__0 
       (.I0(\alu1/div/add_out [9]),
        .I1(\remden[64]_i_1__0_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(a1bus_0[9]),
        .I4(\alu1/div/den [5]),
        .I5(\dso[31]_i_5__0_n_0 ),
        .O(\remden[9]_i_1__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \rgf/a0bus_out/badr[0]_INST_0_i_12 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/sp [0]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(fch_pc0[0]),
        .I4(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[0]_INST_0_i_2 
       (.I0(\badr[0]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/p_1_in [0]),
        .I2(\rgf/bank02/p_0_in [0]),
        .I3(\rgf/a0bus_sr [0]),
        .I4(\rgf/a0bus_b13 [0]),
        .I5(\rgf/a0bus_out/badr[0]_INST_0_i_12_n_0 ),
        .O(a0bus_0[0]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[10]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc0[10]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[10]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[10]_INST_0_i_2 
       (.I0(\badr[10]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [10]),
        .I2(\rgf/bank02/p_0_in [10]),
        .I3(\rgf/a0bus_sr [10]),
        .I4(\rgf/a0bus_b13 [10]),
        .I5(\rgf/a0bus_out/badr[10]_INST_0_i_14_n_0 ),
        .O(a0bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[11]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc0[11]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[11]_INST_0_i_2 
       (.I0(\badr[11]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [11]),
        .I2(\rgf/bank02/p_0_in [11]),
        .I3(\rgf/a0bus_sr [11]),
        .I4(\rgf/a0bus_b13 [11]),
        .I5(\rgf/a0bus_out/badr[11]_INST_0_i_14_n_0 ),
        .O(a0bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[12]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc0[12]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[12]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[12]_INST_0_i_2 
       (.I0(\badr[12]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [12]),
        .I2(\rgf/bank02/p_0_in [12]),
        .I3(\rgf/a0bus_sr [12]),
        .I4(\rgf/a0bus_b13 [12]),
        .I5(\rgf/a0bus_out/badr[12]_INST_0_i_14_n_0 ),
        .O(a0bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[13]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc0[13]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[13]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[13]_INST_0_i_2 
       (.I0(\badr[13]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [13]),
        .I2(\rgf/bank02/p_0_in [13]),
        .I3(\rgf/a0bus_sr [13]),
        .I4(\rgf/a0bus_b13 [13]),
        .I5(\rgf/a0bus_out/badr[13]_INST_0_i_14_n_0 ),
        .O(a0bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[14]_INST_0_i_12 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc0[14]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[14]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[14]_INST_0_i_2 
       (.I0(\badr[14]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/p_1_in [14]),
        .I2(\rgf/bank02/p_0_in [14]),
        .I3(\rgf/a0bus_sr [14]),
        .I4(\rgf/a0bus_b13 [14]),
        .I5(\rgf/a0bus_out/badr[14]_INST_0_i_12_n_0 ),
        .O(a0bus_0[14]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[15]_INST_0_i_13 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc0[15]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[15]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[15]_INST_0_i_2 
       (.I0(\badr[15]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank02/p_1_in [15]),
        .I2(\rgf/bank02/p_0_in [15]),
        .I3(\rgf/a0bus_sr [15]),
        .I4(\rgf/a0bus_b13 [15]),
        .I5(\rgf/a0bus_out/badr[15]_INST_0_i_13_n_0 ),
        .O(a0bus_0[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[16]_INST_0_i_2 
       (.I0(\badr[16]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [16]),
        .O(a0bus_0[16]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[17]_INST_0_i_2 
       (.I0(\badr[17]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [17]),
        .O(a0bus_0[17]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[18]_INST_0_i_2 
       (.I0(\badr[18]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [18]),
        .O(a0bus_0[18]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[19]_INST_0_i_2 
       (.I0(\badr[19]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [19]),
        .O(a0bus_0[19]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[1]_INST_0_i_12 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc0[1]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[1]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[1]_INST_0_i_2 
       (.I0(\badr[1]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/p_1_in [1]),
        .I2(\rgf/bank02/p_0_in [1]),
        .I3(\rgf/a0bus_sr [1]),
        .I4(\rgf/a0bus_b13 [1]),
        .I5(\rgf/a0bus_out/badr[1]_INST_0_i_12_n_0 ),
        .O(a0bus_0[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[20]_INST_0_i_2 
       (.I0(\badr[20]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [20]),
        .O(a0bus_0[20]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[21]_INST_0_i_2 
       (.I0(\badr[21]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [21]),
        .O(a0bus_0[21]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[22]_INST_0_i_2 
       (.I0(\badr[22]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [22]),
        .O(a0bus_0[22]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[23]_INST_0_i_2 
       (.I0(\badr[23]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [23]),
        .O(a0bus_0[23]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[24]_INST_0_i_2 
       (.I0(\badr[24]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [24]),
        .O(a0bus_0[24]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[25]_INST_0_i_2 
       (.I0(\badr[25]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [25]),
        .O(a0bus_0[25]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[26]_INST_0_i_2 
       (.I0(\badr[26]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [26]),
        .O(a0bus_0[26]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[27]_INST_0_i_2 
       (.I0(\badr[27]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [27]),
        .O(a0bus_0[27]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[28]_INST_0_i_2 
       (.I0(\badr[28]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [28]),
        .O(a0bus_0[28]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[29]_INST_0_i_2 
       (.I0(\badr[29]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [29]),
        .O(a0bus_0[29]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[2]_INST_0_i_12 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc0[2]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[2]_INST_0_i_2 
       (.I0(\badr[2]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/p_1_in [2]),
        .I2(\rgf/bank02/p_0_in [2]),
        .I3(\rgf/a0bus_sr [2]),
        .I4(\rgf/a0bus_b13 [2]),
        .I5(\rgf/a0bus_out/badr[2]_INST_0_i_12_n_0 ),
        .O(a0bus_0[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[30]_INST_0_i_2 
       (.I0(\badr[30]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_12_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_13_n_0 ),
        .I5(\rgf/a0bus_sp [30]),
        .O(a0bus_0[30]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[31]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_12_n_0 ),
        .I2(\rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_13_n_0 ),
        .I3(\rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_15_n_0 ),
        .I5(\rgf/a0bus_sp [31]),
        .O(a0bus_0[31]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[3]_INST_0_i_12 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc0[3]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[3]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[3]_INST_0_i_2 
       (.I0(\badr[3]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/p_1_in [3]),
        .I2(\rgf/bank02/p_0_in [3]),
        .I3(\rgf/a0bus_sr [3]),
        .I4(\rgf/a0bus_b13 [3]),
        .I5(\rgf/a0bus_out/badr[3]_INST_0_i_12_n_0 ),
        .O(a0bus_0[3]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[4]_INST_0_i_12 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc0[4]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[4]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[4]_INST_0_i_2 
       (.I0(\badr[4]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/p_1_in [4]),
        .I2(\rgf/bank02/p_0_in [4]),
        .I3(\rgf/a0bus_sr [4]),
        .I4(\rgf/a0bus_b13 [4]),
        .I5(\rgf/a0bus_out/badr[4]_INST_0_i_12_n_0 ),
        .O(a0bus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[5]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc0[5]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[5]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[5]_INST_0_i_2 
       (.I0(\badr[5]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [5]),
        .I2(\rgf/bank02/p_0_in [5]),
        .I3(\rgf/a0bus_sr [5]),
        .I4(\rgf/a0bus_b13 [5]),
        .I5(\rgf/a0bus_out/badr[5]_INST_0_i_14_n_0 ),
        .O(a0bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[6]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc0[6]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[6]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[6]_INST_0_i_2 
       (.I0(\badr[6]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [6]),
        .I2(\rgf/bank02/p_0_in [6]),
        .I3(\rgf/a0bus_sr [6]),
        .I4(\rgf/a0bus_b13 [6]),
        .I5(\rgf/a0bus_out/badr[6]_INST_0_i_14_n_0 ),
        .O(a0bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[7]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc0[7]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[7]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[7]_INST_0_i_2 
       (.I0(\badr[7]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [7]),
        .I2(\rgf/bank02/p_0_in [7]),
        .I3(\rgf/a0bus_sr [7]),
        .I4(\rgf/a0bus_b13 [7]),
        .I5(\rgf/a0bus_out/badr[7]_INST_0_i_14_n_0 ),
        .O(a0bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[8]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc0[8]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[8]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[8]_INST_0_i_2 
       (.I0(\badr[8]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [8]),
        .I2(\rgf/bank02/p_0_in [8]),
        .I3(\rgf/a0bus_sr [8]),
        .I4(\rgf/a0bus_b13 [8]),
        .I5(\rgf/a0bus_out/badr[8]_INST_0_i_14_n_0 ),
        .O(a0bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a0bus_out/badr[9]_INST_0_i_14 
       (.I0(\rgf/a0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/a0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc0[9]),
        .I5(\rgf/a0bus_sel_cr [1]),
        .O(\rgf/a0bus_out/badr[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a0bus_out/badr[9]_INST_0_i_2 
       (.I0(\badr[9]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/p_1_in [9]),
        .I2(\rgf/bank02/p_0_in [9]),
        .I3(\rgf/a0bus_sr [9]),
        .I4(\rgf/a0bus_b13 [9]),
        .I5(\rgf/a0bus_out/badr[9]_INST_0_i_14_n_0 ),
        .O(a0bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/a1bus_out/badr[0]_INST_0_i_1 
       (.I0(\badr[0]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [0]),
        .I2(\rgf/a1bus_sel_cr [0]),
        .I3(\rgf/sreg/sr [0]),
        .I4(\rgf/a1bus_b13 [0]),
        .I5(\rgf/a1bus_out/badr[0]_INST_0_i_6_n_0 ),
        .O(a1bus_0[0]));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \rgf/a1bus_out/badr[0]_INST_0_i_6 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/sp [0]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(fch_pc1[0]),
        .I4(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[10]_INST_0_i_1 
       (.I0(\badr[10]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [10]),
        .I2(\rgf/bank02/p_0_in0_in [10]),
        .I3(\rgf/a1bus_sr [10]),
        .I4(\rgf/a1bus_b13 [10]),
        .I5(\rgf/a1bus_out/badr[10]_INST_0_i_8_n_0 ),
        .O(a1bus_0[10]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[10]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc1[10]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[11]_INST_0_i_1 
       (.I0(\badr[11]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [11]),
        .I2(\rgf/bank02/p_0_in0_in [11]),
        .I3(\rgf/a1bus_sr [11]),
        .I4(\rgf/a1bus_b13 [11]),
        .I5(\rgf/a1bus_out/badr[11]_INST_0_i_8_n_0 ),
        .O(a1bus_0[11]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[11]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc1[11]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[11]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[12]_INST_0_i_1 
       (.I0(\badr[12]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [12]),
        .I2(\rgf/bank02/p_0_in0_in [12]),
        .I3(\rgf/a1bus_sr [12]),
        .I4(\rgf/a1bus_b13 [12]),
        .I5(\rgf/a1bus_out/badr[12]_INST_0_i_8_n_0 ),
        .O(a1bus_0[12]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[12]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc1[12]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[12]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[13]_INST_0_i_1 
       (.I0(\badr[13]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [13]),
        .I2(\rgf/bank02/p_0_in0_in [13]),
        .I3(\rgf/a1bus_sr [13]),
        .I4(\rgf/a1bus_b13 [13]),
        .I5(\rgf/a1bus_out/badr[13]_INST_0_i_8_n_0 ),
        .O(a1bus_0[13]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[13]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc1[13]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[13]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/a1bus_out/badr[14]_INST_0_i_1 
       (.I0(\rgf/a1bus_out/badr[14]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [14]),
        .I2(\rgf/a1bus_sel_cr [0]),
        .I3(\rgf/sreg/sr [14]),
        .I4(\rgf/a1bus_b13 [14]),
        .I5(\rgf/a1bus_out/badr[14]_INST_0_i_6_n_0 ),
        .O(a1bus_0[14]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \rgf/a1bus_out/badr[14]_INST_0_i_3 
       (.I0(\rgf/treg/tr [14]),
        .I1(\rgf/ivec/iv [14]),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .I5(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_out/badr[14]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[14]_INST_0_i_6 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc1[14]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[14]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/a1bus_out/badr[15]_INST_0_i_1 
       (.I0(\rgf/a1bus_out/badr[15]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [15]),
        .I2(\rgf/a1bus_sel_cr [0]),
        .I3(\rgf/sreg/sr [15]),
        .I4(\rgf/a1bus_b13 [15]),
        .I5(\rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ),
        .O(a1bus_0[15]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \rgf/a1bus_out/badr[15]_INST_0_i_3 
       (.I0(\rgf/treg/tr [15]),
        .I1(\rgf/ivec/iv [15]),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .I5(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_out/badr[15]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[15]_INST_0_i_7 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc1[15]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[16]_INST_0_i_1 
       (.I0(\badr[16]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [16]),
        .O(a1bus_0[16]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[17]_INST_0_i_1 
       (.I0(\badr[17]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [17]),
        .O(a1bus_0[17]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[18]_INST_0_i_1 
       (.I0(\badr[18]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [18]),
        .O(a1bus_0[18]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[19]_INST_0_i_1 
       (.I0(\badr[19]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [19]),
        .O(a1bus_0[19]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/a1bus_out/badr[1]_INST_0_i_1 
       (.I0(\rgf/a1bus_out/badr[1]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [1]),
        .I2(\rgf/a1bus_sel_cr [0]),
        .I3(\rgf/sreg/sr [1]),
        .I4(\rgf/a1bus_b13 [1]),
        .I5(\rgf/a1bus_out/badr[1]_INST_0_i_6_n_0 ),
        .O(a1bus_0[1]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \rgf/a1bus_out/badr[1]_INST_0_i_3 
       (.I0(\rgf/treg/tr [1]),
        .I1(\rgf/ivec/iv [1]),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .I5(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_out/badr[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[1]_INST_0_i_6 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc1[1]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[20]_INST_0_i_1 
       (.I0(\badr[20]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [20]),
        .O(a1bus_0[20]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[21]_INST_0_i_1 
       (.I0(\badr[21]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [21]),
        .O(a1bus_0[21]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[22]_INST_0_i_1 
       (.I0(\badr[22]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [22]),
        .O(a1bus_0[22]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[23]_INST_0_i_1 
       (.I0(\badr[23]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [23]),
        .O(a1bus_0[23]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[24]_INST_0_i_1 
       (.I0(\badr[24]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [24]),
        .O(a1bus_0[24]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[25]_INST_0_i_1 
       (.I0(\badr[25]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [25]),
        .O(a1bus_0[25]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[26]_INST_0_i_1 
       (.I0(\badr[26]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [26]),
        .O(a1bus_0[26]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[27]_INST_0_i_1 
       (.I0(\badr[27]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [27]),
        .O(a1bus_0[27]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[28]_INST_0_i_1 
       (.I0(\badr[28]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [28]),
        .O(a1bus_0[28]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[29]_INST_0_i_1 
       (.I0(\badr[29]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [29]),
        .O(a1bus_0[29]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/a1bus_out/badr[2]_INST_0_i_1 
       (.I0(\rgf/a1bus_out/badr[2]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [2]),
        .I2(\rgf/a1bus_sel_cr [0]),
        .I3(\rgf/sreg/sr [2]),
        .I4(\rgf/a1bus_b13 [2]),
        .I5(\rgf/a1bus_out/badr[2]_INST_0_i_6_n_0 ),
        .O(a1bus_0[2]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \rgf/a1bus_out/badr[2]_INST_0_i_3 
       (.I0(\rgf/treg/tr [2]),
        .I1(\rgf/ivec/iv [2]),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .I5(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_out/badr[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[2]_INST_0_i_6 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc1[2]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[30]_INST_0_i_1 
       (.I0(\badr[30]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_4_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_5_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_6_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_7_n_0 ),
        .I5(\rgf/a1bus_sp [30]),
        .O(a1bus_0[30]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[31]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_5_n_0 ),
        .I1(\rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_6_n_0 ),
        .I2(\rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_7_n_0 ),
        .I3(\rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_8_n_0 ),
        .I4(\rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_9_n_0 ),
        .I5(\rgf/a1bus_sp [31]),
        .O(a1bus_0[31]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/a1bus_out/badr[3]_INST_0_i_1 
       (.I0(\rgf/a1bus_out/badr[3]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [3]),
        .I2(\rgf/a1bus_sel_cr [0]),
        .I3(\rgf/sreg/sr [3]),
        .I4(\rgf/a1bus_b13 [3]),
        .I5(\rgf/a1bus_out/badr[3]_INST_0_i_6_n_0 ),
        .O(a1bus_0[3]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \rgf/a1bus_out/badr[3]_INST_0_i_3 
       (.I0(\rgf/treg/tr [3]),
        .I1(\rgf/ivec/iv [3]),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .I5(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_out/badr[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[3]_INST_0_i_6 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc1[3]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/a1bus_out/badr[4]_INST_0_i_1 
       (.I0(\rgf/a1bus_out/badr[4]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [4]),
        .I2(\rgf/a1bus_sel_cr [0]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\rgf/a1bus_b13 [4]),
        .I5(\rgf/a1bus_out/badr[4]_INST_0_i_6_n_0 ),
        .O(a1bus_0[4]));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \rgf/a1bus_out/badr[4]_INST_0_i_3 
       (.I0(\rgf/treg/tr [4]),
        .I1(\rgf/ivec/iv [4]),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .I5(\badr[31]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_out/badr[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[4]_INST_0_i_6 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc1[4]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[4]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[5]_INST_0_i_1 
       (.I0(\badr[5]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [5]),
        .I2(\rgf/bank02/p_0_in0_in [5]),
        .I3(\rgf/a1bus_sr [5]),
        .I4(\rgf/a1bus_b13 [5]),
        .I5(\rgf/a1bus_out/badr[5]_INST_0_i_8_n_0 ),
        .O(a1bus_0[5]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[5]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc1[5]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[5]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[6]_INST_0_i_1 
       (.I0(\badr[6]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [6]),
        .I2(\rgf/bank02/p_0_in0_in [6]),
        .I3(\rgf/a1bus_sr [6]),
        .I4(\rgf/a1bus_b13 [6]),
        .I5(\rgf/a1bus_out/badr[6]_INST_0_i_8_n_0 ),
        .O(a1bus_0[6]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[6]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc1[6]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[7]_INST_0_i_1 
       (.I0(\badr[7]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [7]),
        .I2(\rgf/bank02/p_0_in0_in [7]),
        .I3(\rgf/a1bus_sr [7]),
        .I4(\rgf/a1bus_b13 [7]),
        .I5(\rgf/a1bus_out/badr[7]_INST_0_i_8_n_0 ),
        .O(a1bus_0[7]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[7]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc1[7]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[8]_INST_0_i_1 
       (.I0(\badr[8]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [8]),
        .I2(\rgf/bank02/p_0_in0_in [8]),
        .I3(\rgf/a1bus_sr [8]),
        .I4(\rgf/a1bus_b13 [8]),
        .I5(\rgf/a1bus_out/badr[8]_INST_0_i_8_n_0 ),
        .O(a1bus_0[8]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[8]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc1[8]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/badr[9]_INST_0_i_1 
       (.I0(\badr[9]_INST_0_i_3_n_0 ),
        .I1(\rgf/bank02/p_1_in1_in [9]),
        .I2(\rgf/bank02/p_0_in0_in [9]),
        .I3(\rgf/a1bus_sr [9]),
        .I4(\rgf/a1bus_b13 [9]),
        .I5(\rgf/a1bus_out/badr[9]_INST_0_i_8_n_0 ),
        .O(a1bus_0[9]));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/a1bus_out/badr[9]_INST_0_i_8 
       (.I0(\rgf/a1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/a1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc1[9]),
        .I5(\rgf/a1bus_sel_cr [1]),
        .O(\rgf/a1bus_out/badr[9]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[10]_i_32 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[10]_i_34_n_0 ),
        .I4(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_13_n_0 ),
        .I5(\rgf/a1bus_out/badr[14]_INST_0_i_3_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[10]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[10]_i_33 
       (.I0(\rgf/a1bus_sr [14]),
        .I1(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_23_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_36_n_0 ),
        .I5(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_19_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[10]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[19]_i_39 
       (.I0(\rgf/a1bus_sr [15]),
        .I1(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_27_n_0 ),
        .I2(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_26_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_25_n_0 ),
        .I4(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[19]_i_43_n_0 ),
        .I5(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_22_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[19]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_43 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_19_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_53_n_0 ),
        .I4(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_16_n_0 ),
        .I5(\rgf/a1bus_out/badr[15]_INST_0_i_3_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_44 
       (.I0(\rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_22_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[19]_i_43_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_25_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_54_n_0 ),
        .I5(\rgf/a1bus_sr [15]),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_45 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_55_n_0 ),
        .I4(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_13_n_0 ),
        .I5(\rgf/a1bus_out/badr[2]_INST_0_i_3_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_46 
       (.I0(\rgf/a1bus_sr [2]),
        .I1(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_23_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_57_n_0 ),
        .I5(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_19_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_47 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_58_n_0 ),
        .I4(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_13_n_0 ),
        .I5(\rgf/a1bus_out/badr[1]_INST_0_i_3_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_48 
       (.I0(\rgf/a1bus_out/badr[1]_INST_0_i_6_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_19_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_59_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_60_n_0 ),
        .I5(\rgf/a1bus_sr [1]),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_49 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_62_n_0 ),
        .I4(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_13_n_0 ),
        .I5(\rgf/a1bus_out/badr[4]_INST_0_i_3_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_50 
       (.I0(\rgf/a1bus_sr [4]),
        .I1(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_23_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_64_n_0 ),
        .I5(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_19_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_51 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_65_n_0 ),
        .I4(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_13_n_0 ),
        .I5(\rgf/a1bus_out/badr[3]_INST_0_i_3_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[28]_i_52 
       (.I0(\rgf/a1bus_out/badr[3]_INST_0_i_6_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_19_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_66_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_67_n_0 ),
        .I5(\rgf/a1bus_sr [3]),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/a1bus_out/rgf_c1bus_wb[4]_i_28 
       (.I0(\rgf/a1bus_sr [0]),
        .I1(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_23_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[4]_i_29_n_0 ),
        .I5(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_19_n_0 ),
        .O(\rgf/a1bus_out/rgf_c1bus_wb[4]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \rgf/b0bus_out/bbus_o[0]_INST_0_i_17 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/sp [0]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(fch_pc0[0]),
        .I4(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[0]_INST_0_i_3 
       (.I0(\rgf/treg/tr [0]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [0]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[0]_INST_0_i_6 
       (.I0(\rgf/b0bus_out/bbus_o[0]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18_n_0 ),
        .I2(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_20_n_0 ),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_21_n_0 ),
        .I5(\rgf/b0bus_sr ),
        .O(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[1]_INST_0_i_11 
       (.I0(\rgf/treg/tr [1]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [1]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[1]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[1]_INST_0_i_3 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_8_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9_n_0 ),
        .I3(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[1]_INST_0_i_11_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/b0bus_out/bbus_o[1]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [1]),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_14_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_15_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[1]_INST_0_i_5 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc0[1]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[1]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[2]_INST_0_i_11 
       (.I0(\rgf/treg/tr [2]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [2]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[2]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[2]_INST_0_i_3 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_8_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9_n_0 ),
        .I3(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[2]_INST_0_i_11_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/b0bus_out/bbus_o[2]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [2]),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_14_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_15_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[2]_INST_0_i_5 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc0[2]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[2]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[3]_INST_0_i_12 
       (.I0(\rgf/treg/tr [3]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [3]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[3]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[3]_INST_0_i_3 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_9_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10_n_0 ),
        .I3(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[3]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/b0bus_out/bbus_o[3]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [3]),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_13_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_15_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_16_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[3]_INST_0_i_5 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc0[3]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[3]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[4]_INST_0_i_11 
       (.I0(\rgf/treg/tr [4]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [4]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[4]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[4]_INST_0_i_3 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_7_n_0 ),
        .I1(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_8_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9_n_0 ),
        .I3(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[4]_INST_0_i_11_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[4]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/b0bus_out/bbus_o[4]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_14_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_15_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[4]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[4]_INST_0_i_5 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc0[4]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[4]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b0bus_out/bbus_o[5]_INST_0_i_18 
       (.I0(\rgf/treg/tr [5]),
        .I1(\rgf/b0bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [5]),
        .I3(\rgf/b0bus_sel_cr [3]),
        .O(\rgf/b0bus_out/bbus_o[5]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/b0bus_out/bbus_o[5]_INST_0_i_4 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_15_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_17_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[5]_INST_0_i_18_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[5]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf/b0bus_out/bbus_o[5]_INST_0_i_5 
       (.I0(\rgf/b0bus_sel_cr [0]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_19_n_0 ),
        .I3(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_20_n_0 ),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22_n_0 ),
        .O(\rgf/b0bus_out/bbus_o[5]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[5]_INST_0_i_6 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc0[5]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[5]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bbus_o[6]_INST_0_i_3 
       (.I0(\rgf/bank02/p_0_in2_in [6]),
        .I1(\rgf/bank02/p_1_in3_in [6]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [6]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [6]),
        .O(\rgf/b0bus_out/bbus_o[6]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bbus_o[6]_INST_0_i_4 
       (.I0(\rgf/b0bus_out/bbus_o[6]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [6]),
        .I2(\rgf/bank13/p_0_in2_in [6]),
        .I3(\rgf/sreg/sr [6]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bbus_o[6]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[6]_INST_0_i_8 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc0[6]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bbus_o[7]_INST_0_i_3 
       (.I0(\rgf/bank02/p_0_in2_in [7]),
        .I1(\rgf/bank02/p_1_in3_in [7]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [7]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [7]),
        .O(\rgf/b0bus_out/bbus_o[7]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bbus_o[7]_INST_0_i_4 
       (.I0(\rgf/b0bus_out/bbus_o[7]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [7]),
        .I2(\rgf/bank13/p_0_in2_in [7]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bbus_o[7]_INST_0_i_8 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc0[7]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bbus_o[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[10]_INST_0_i_10 
       (.I0(\rgf/bank02/p_0_in2_in [10]),
        .I1(\rgf/bank02/p_1_in3_in [10]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [10]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [10]),
        .O(\rgf/b0bus_out/bdatw[10]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[10]_INST_0_i_11 
       (.I0(\rgf/b0bus_out/bdatw[10]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [10]),
        .I2(\rgf/bank13/p_0_in2_in [10]),
        .I3(\rgf/sreg/sr [10]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[10]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[10]_INST_0_i_22 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc0[10]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[10]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[11]_INST_0_i_10 
       (.I0(\rgf/bank02/p_0_in2_in [11]),
        .I1(\rgf/bank02/p_1_in3_in [11]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [11]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [11]),
        .O(\rgf/b0bus_out/bdatw[11]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[11]_INST_0_i_11 
       (.I0(\rgf/b0bus_out/bdatw[11]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [11]),
        .I2(\rgf/bank13/p_0_in2_in [11]),
        .I3(\rgf/sreg/sr [11]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[11]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[11]_INST_0_i_22 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc0[11]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[11]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[12]_INST_0_i_10 
       (.I0(\rgf/b0bus_out/bdatw[12]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [12]),
        .I2(\rgf/bank13/p_0_in2_in [12]),
        .I3(\rgf/sreg/sr [12]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[12]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[12]_INST_0_i_26 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc0[12]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[12]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[12]_INST_0_i_9 
       (.I0(\rgf/bank02/p_0_in2_in [12]),
        .I1(\rgf/bank02/p_1_in3_in [12]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [12]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [12]),
        .O(\rgf/b0bus_out/bdatw[12]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[13]_INST_0_i_17 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc0[13]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[13]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[13]_INST_0_i_8 
       (.I0(\rgf/bank02/p_0_in2_in [13]),
        .I1(\rgf/bank02/p_1_in3_in [13]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [13]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [13]),
        .O(\rgf/b0bus_out/bdatw[13]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[13]_INST_0_i_9 
       (.I0(\rgf/b0bus_out/bdatw[13]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [13]),
        .I2(\rgf/bank13/p_0_in2_in [13]),
        .I3(\rgf/sreg/sr [13]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[13]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[14]_INST_0_i_10 
       (.I0(\rgf/b0bus_out/bdatw[14]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [14]),
        .I2(\rgf/bank13/p_0_in2_in [14]),
        .I3(\rgf/sreg/sr [14]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[14]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[14]_INST_0_i_18 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc0[14]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[14]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[14]_INST_0_i_9 
       (.I0(\rgf/bank02/p_0_in2_in [14]),
        .I1(\rgf/bank02/p_1_in3_in [14]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [14]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [14]),
        .O(\rgf/b0bus_out/bdatw[14]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[15]_INST_0_i_12 
       (.I0(\rgf/bank02/p_0_in2_in [15]),
        .I1(\rgf/bank02/p_1_in3_in [15]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [15]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [15]),
        .O(\rgf/b0bus_out/bdatw[15]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[15]_INST_0_i_13 
       (.I0(\rgf/b0bus_out/bdatw[15]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [15]),
        .I2(\rgf/bank13/p_0_in2_in [15]),
        .I3(\rgf/sreg/sr [15]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[15]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[15]_INST_0_i_26 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc0[15]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[15]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[16]_INST_0_i_3 
       (.I0(\bdatw[16]_INST_0_i_7_n_0 ),
        .I1(\bdatw[16]_INST_0_i_8_n_0 ),
        .I2(\bdatw[16]_INST_0_i_9_n_0 ),
        .I3(\bdatw[16]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [16]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[16]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[16]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [16]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [16]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[16]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[17]_INST_0_i_3 
       (.I0(\bdatw[17]_INST_0_i_7_n_0 ),
        .I1(\bdatw[17]_INST_0_i_8_n_0 ),
        .I2(\bdatw[17]_INST_0_i_9_n_0 ),
        .I3(\bdatw[17]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [17]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[17]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[17]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [17]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [17]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[17]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[18]_INST_0_i_3 
       (.I0(\bdatw[18]_INST_0_i_7_n_0 ),
        .I1(\bdatw[18]_INST_0_i_8_n_0 ),
        .I2(\bdatw[18]_INST_0_i_9_n_0 ),
        .I3(\bdatw[18]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [18]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[18]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[18]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [18]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [18]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[18]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[19]_INST_0_i_3 
       (.I0(\bdatw[19]_INST_0_i_7_n_0 ),
        .I1(\bdatw[19]_INST_0_i_8_n_0 ),
        .I2(\bdatw[19]_INST_0_i_9_n_0 ),
        .I3(\bdatw[19]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [19]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[19]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[19]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [19]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [19]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[19]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[20]_INST_0_i_3 
       (.I0(\bdatw[20]_INST_0_i_7_n_0 ),
        .I1(\bdatw[20]_INST_0_i_8_n_0 ),
        .I2(\bdatw[20]_INST_0_i_9_n_0 ),
        .I3(\bdatw[20]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [20]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[20]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[20]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [20]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [20]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[20]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[21]_INST_0_i_3 
       (.I0(\bdatw[21]_INST_0_i_7_n_0 ),
        .I1(\bdatw[21]_INST_0_i_8_n_0 ),
        .I2(\bdatw[21]_INST_0_i_9_n_0 ),
        .I3(\bdatw[21]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [21]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[21]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[21]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [21]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [21]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[21]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[22]_INST_0_i_3 
       (.I0(\bdatw[22]_INST_0_i_7_n_0 ),
        .I1(\bdatw[22]_INST_0_i_8_n_0 ),
        .I2(\bdatw[22]_INST_0_i_9_n_0 ),
        .I3(\bdatw[22]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [22]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[22]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[22]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [22]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [22]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[22]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[23]_INST_0_i_3 
       (.I0(\bdatw[23]_INST_0_i_7_n_0 ),
        .I1(\bdatw[23]_INST_0_i_8_n_0 ),
        .I2(\bdatw[23]_INST_0_i_9_n_0 ),
        .I3(\bdatw[23]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [23]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[23]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[23]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [23]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [23]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[23]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[24]_INST_0_i_3 
       (.I0(\bdatw[24]_INST_0_i_7_n_0 ),
        .I1(\bdatw[24]_INST_0_i_8_n_0 ),
        .I2(\bdatw[24]_INST_0_i_9_n_0 ),
        .I3(\bdatw[24]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [24]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[24]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[24]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [24]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [24]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[24]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[25]_INST_0_i_3 
       (.I0(\bdatw[25]_INST_0_i_7_n_0 ),
        .I1(\bdatw[25]_INST_0_i_8_n_0 ),
        .I2(\bdatw[25]_INST_0_i_9_n_0 ),
        .I3(\bdatw[25]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [25]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[25]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[25]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [25]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [25]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[25]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[26]_INST_0_i_3 
       (.I0(\bdatw[26]_INST_0_i_7_n_0 ),
        .I1(\bdatw[26]_INST_0_i_8_n_0 ),
        .I2(\bdatw[26]_INST_0_i_9_n_0 ),
        .I3(\bdatw[26]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [26]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[26]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[26]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [26]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [26]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[26]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[27]_INST_0_i_3 
       (.I0(\bdatw[27]_INST_0_i_7_n_0 ),
        .I1(\bdatw[27]_INST_0_i_8_n_0 ),
        .I2(\bdatw[27]_INST_0_i_9_n_0 ),
        .I3(\bdatw[27]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [27]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[27]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[27]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [27]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [27]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[27]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[28]_INST_0_i_3 
       (.I0(\bdatw[28]_INST_0_i_7_n_0 ),
        .I1(\bdatw[28]_INST_0_i_8_n_0 ),
        .I2(\bdatw[28]_INST_0_i_9_n_0 ),
        .I3(\bdatw[28]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [28]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[28]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[28]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [28]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [28]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[28]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[29]_INST_0_i_3 
       (.I0(\bdatw[29]_INST_0_i_7_n_0 ),
        .I1(\bdatw[29]_INST_0_i_8_n_0 ),
        .I2(\bdatw[29]_INST_0_i_9_n_0 ),
        .I3(\bdatw[29]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [29]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[29]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[29]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [29]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [29]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[29]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[30]_INST_0_i_3 
       (.I0(\bdatw[30]_INST_0_i_7_n_0 ),
        .I1(\bdatw[30]_INST_0_i_8_n_0 ),
        .I2(\bdatw[30]_INST_0_i_9_n_0 ),
        .I3(\bdatw[30]_INST_0_i_10_n_0 ),
        .I4(\rgf/treg/tr [30]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[30]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[30]_INST_0_i_4 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [30]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [30]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_12_n_0 ),
        .O(\rgf/b0bus_out/bdatw[30]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b0bus_out/bdatw[31]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_14_n_0 ),
        .I1(\bdatw[31]_INST_0_i_15_n_0 ),
        .I2(\bdatw[31]_INST_0_i_16_n_0 ),
        .I3(\bdatw[31]_INST_0_i_17_n_0 ),
        .I4(\rgf/treg/tr [31]),
        .I5(\rgf/b0bus_sel_cr [4]),
        .O(\rgf/b0bus_out/bdatw[31]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b0bus_out/bdatw[31]_INST_0_i_5 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [31]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [31]),
        .I4(\rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_22_n_0 ),
        .O(\rgf/b0bus_out/bdatw[31]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[8]_INST_0_i_18 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc0[8]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[8]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[8]_INST_0_i_7 
       (.I0(\rgf/bank02/p_0_in2_in [8]),
        .I1(\rgf/bank02/p_1_in3_in [8]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [8]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [8]),
        .O(\rgf/b0bus_out/bdatw[8]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[8]_INST_0_i_8 
       (.I0(\rgf/b0bus_out/bdatw[8]_INST_0_i_18_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [8]),
        .I2(\rgf/bank13/p_0_in2_in [8]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[8]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b0bus_out/bdatw[9]_INST_0_i_20 
       (.I0(\rgf/b0bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/b0bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc0[9]),
        .I5(\rgf/b0bus_sel_cr [1]),
        .O(\rgf/b0bus_out/bdatw[9]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b0bus_out/bdatw[9]_INST_0_i_8 
       (.I0(\rgf/bank02/p_0_in2_in [9]),
        .I1(\rgf/bank02/p_1_in3_in [9]),
        .I2(\rgf/b0bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [9]),
        .I4(\rgf/b0bus_sel_cr [4]),
        .I5(\rgf/treg/tr [9]),
        .O(\rgf/b0bus_out/bdatw[9]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b0bus_out/bdatw[9]_INST_0_i_9 
       (.I0(\rgf/b0bus_out/bdatw[9]_INST_0_i_20_n_0 ),
        .I1(\rgf/bank13/p_1_in3_in [9]),
        .I2(\rgf/bank13/p_0_in2_in [9]),
        .I3(\rgf/sreg/sr [9]),
        .I4(\rgf/b0bus_sel_cr [0]),
        .O(\rgf/b0bus_out/bdatw[9]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf/b0bus_out/rgf_c0bus_wb[31]_i_77 
       (.I0(\rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_80_n_0 ),
        .I1(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_81_n_0 ),
        .I3(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_12_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[0]_INST_0_i_3_n_0 ),
        .O(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_14 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [10]),
        .I4(fch_pc1[10]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_7 
       (.I0(\rgf/b1bus_out/bdatw[10]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_15_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_16_n_0 ),
        .I3(\rgf/sreg/sr [10]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[10]_INST_0_i_8 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_18_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [10]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [10]),
        .O(\rgf/b1bus_out/bdatw[10]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_13 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [11]),
        .I4(fch_pc1[11]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_7 
       (.I0(\rgf/b1bus_out/bdatw[11]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_15_n_0 ),
        .I3(\rgf/sreg/sr [11]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[11]_INST_0_i_8 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_16_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_17_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [11]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [11]),
        .O(\rgf/b1bus_out/bdatw[11]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_12 
       (.I0(\rgf/treg/tr [4]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [4]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_15 
       (.I0(\rgf/b1bus_out/bdatw[12]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_42_n_0 ),
        .I5(\rgf/b1bus_sr [4]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_19 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [12]),
        .I4(fch_pc1[12]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_38 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [4]),
        .I4(fch_pc1[4]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_6 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_18_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [12]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [12]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[12]_INST_0_i_7 
       (.I0(\rgf/b1bus_out/bdatw[12]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_21_n_0 ),
        .I3(\rgf/sreg/sr [12]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[12]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_12 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [13]),
        .I4(fch_pc1[13]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_5 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_10_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_11_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [13]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [13]),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[13]_INST_0_i_6 
       (.I0(\rgf/b1bus_out/bdatw[13]_INST_0_i_12_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_13_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_14_n_0 ),
        .I3(\rgf/sreg/sr [13]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[13]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_11 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [14]),
        .I4(fch_pc1[14]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_6 
       (.I0(\rgf/b1bus_out/bdatw[14]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_12_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_13_n_0 ),
        .I3(\rgf/sreg/sr [14]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[14]_INST_0_i_7 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_15_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [14]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [14]),
        .O(\rgf/b1bus_out/bdatw[14]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_10 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_20_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [15]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [15]),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_15 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [15]),
        .I4(fch_pc1[15]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[15]_INST_0_i_9 
       (.I0(\rgf/b1bus_out/bdatw[15]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_17_n_0 ),
        .I3(\rgf/sreg/sr [15]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[15]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[16]_INST_0_i_5 
       (.I0(\bdatw[16]_INST_0_i_13_n_0 ),
        .I1(\bdatw[16]_INST_0_i_14_n_0 ),
        .I2(\bdatw[16]_INST_0_i_15_n_0 ),
        .I3(\bdatw[16]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [16]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[16]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[16]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [16]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [16]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[16]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[17]_INST_0_i_5 
       (.I0(\bdatw[17]_INST_0_i_13_n_0 ),
        .I1(\bdatw[17]_INST_0_i_14_n_0 ),
        .I2(\bdatw[17]_INST_0_i_15_n_0 ),
        .I3(\bdatw[17]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [17]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[17]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[17]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [17]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [17]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[17]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[18]_INST_0_i_5 
       (.I0(\bdatw[18]_INST_0_i_13_n_0 ),
        .I1(\bdatw[18]_INST_0_i_14_n_0 ),
        .I2(\bdatw[18]_INST_0_i_15_n_0 ),
        .I3(\bdatw[18]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [18]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[18]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[18]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [18]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [18]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[18]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[19]_INST_0_i_5 
       (.I0(\bdatw[19]_INST_0_i_13_n_0 ),
        .I1(\bdatw[19]_INST_0_i_14_n_0 ),
        .I2(\bdatw[19]_INST_0_i_15_n_0 ),
        .I3(\bdatw[19]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [19]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[19]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[19]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [19]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [19]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[19]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[20]_INST_0_i_5 
       (.I0(\bdatw[20]_INST_0_i_13_n_0 ),
        .I1(\bdatw[20]_INST_0_i_14_n_0 ),
        .I2(\bdatw[20]_INST_0_i_15_n_0 ),
        .I3(\bdatw[20]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [20]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[20]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[20]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [20]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [20]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[20]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[21]_INST_0_i_5 
       (.I0(\bdatw[21]_INST_0_i_13_n_0 ),
        .I1(\bdatw[21]_INST_0_i_14_n_0 ),
        .I2(\bdatw[21]_INST_0_i_15_n_0 ),
        .I3(\bdatw[21]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [21]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[21]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[21]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [21]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [21]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[21]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[22]_INST_0_i_5 
       (.I0(\bdatw[22]_INST_0_i_13_n_0 ),
        .I1(\bdatw[22]_INST_0_i_14_n_0 ),
        .I2(\bdatw[22]_INST_0_i_15_n_0 ),
        .I3(\bdatw[22]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [22]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[22]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[22]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [22]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [22]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[22]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[23]_INST_0_i_5 
       (.I0(\bdatw[23]_INST_0_i_13_n_0 ),
        .I1(\bdatw[23]_INST_0_i_14_n_0 ),
        .I2(\bdatw[23]_INST_0_i_15_n_0 ),
        .I3(\bdatw[23]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [23]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[23]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[23]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [23]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [23]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[23]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[24]_INST_0_i_5 
       (.I0(\bdatw[24]_INST_0_i_13_n_0 ),
        .I1(\bdatw[24]_INST_0_i_14_n_0 ),
        .I2(\bdatw[24]_INST_0_i_15_n_0 ),
        .I3(\bdatw[24]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [24]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[24]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[24]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [24]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [24]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[24]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[25]_INST_0_i_5 
       (.I0(\bdatw[25]_INST_0_i_13_n_0 ),
        .I1(\bdatw[25]_INST_0_i_14_n_0 ),
        .I2(\bdatw[25]_INST_0_i_15_n_0 ),
        .I3(\bdatw[25]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [25]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[25]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[25]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [25]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [25]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[25]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[26]_INST_0_i_5 
       (.I0(\bdatw[26]_INST_0_i_13_n_0 ),
        .I1(\bdatw[26]_INST_0_i_14_n_0 ),
        .I2(\bdatw[26]_INST_0_i_15_n_0 ),
        .I3(\bdatw[26]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [26]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[26]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[26]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [26]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [26]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[26]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[27]_INST_0_i_5 
       (.I0(\bdatw[27]_INST_0_i_13_n_0 ),
        .I1(\bdatw[27]_INST_0_i_14_n_0 ),
        .I2(\bdatw[27]_INST_0_i_15_n_0 ),
        .I3(\bdatw[27]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [27]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[27]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[27]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [27]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [27]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[27]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[28]_INST_0_i_5 
       (.I0(\bdatw[28]_INST_0_i_13_n_0 ),
        .I1(\bdatw[28]_INST_0_i_14_n_0 ),
        .I2(\bdatw[28]_INST_0_i_15_n_0 ),
        .I3(\bdatw[28]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [28]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[28]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[28]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [28]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [28]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[28]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[29]_INST_0_i_5 
       (.I0(\bdatw[29]_INST_0_i_13_n_0 ),
        .I1(\bdatw[29]_INST_0_i_14_n_0 ),
        .I2(\bdatw[29]_INST_0_i_15_n_0 ),
        .I3(\bdatw[29]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [29]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[29]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[29]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [29]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [29]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[29]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[30]_INST_0_i_5 
       (.I0(\bdatw[30]_INST_0_i_13_n_0 ),
        .I1(\bdatw[30]_INST_0_i_14_n_0 ),
        .I2(\bdatw[30]_INST_0_i_15_n_0 ),
        .I3(\bdatw[30]_INST_0_i_16_n_0 ),
        .I4(\rgf/treg/tr [30]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[30]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[30]_INST_0_i_6 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [30]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [30]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_18_n_0 ),
        .O(\rgf/b1bus_out/bdatw[30]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/b1bus_out/bdatw[31]_INST_0_i_10 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [31]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [31]),
        .I4(\rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_38_n_0 ),
        .I5(\rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_39_n_0 ),
        .O(\rgf/b1bus_out/bdatw[31]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \rgf/b1bus_out/bdatw[31]_INST_0_i_9 
       (.I0(\bdatw[31]_INST_0_i_31_n_0 ),
        .I1(\bdatw[31]_INST_0_i_32_n_0 ),
        .I2(\bdatw[31]_INST_0_i_33_n_0 ),
        .I3(\bdatw[31]_INST_0_i_34_n_0 ),
        .I4(\rgf/treg/tr [31]),
        .I5(\rgf/b1bus_sel_cr [4]),
        .O(\rgf/b1bus_out/bdatw[31]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_13 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [8]),
        .I4(fch_pc1[8]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_5 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_12_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [8]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [8]),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[8]_INST_0_i_6 
       (.I0(\rgf/b1bus_out/bdatw[8]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_15_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[8]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_14 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [9]),
        .I4(fch_pc1[9]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_5 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_12_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_13_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [9]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [9]),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/bdatw[9]_INST_0_i_6 
       (.I0(\rgf/b1bus_out/bdatw[9]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_15_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_16_n_0 ),
        .I3(\rgf/sreg/sr [9]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/bdatw[9]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_17 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/sp [0]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(fch_pc1[0]),
        .I4(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_3 
       (.I0(\rgf/treg/tr [0]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [0]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_6 
       (.I0(\rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_18_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_19_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_20_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_21_n_0 ),
        .I5(\rgf/b1bus_sr [0]),
        .O(\rgf/b1bus_out/niss_dsp_b1[0]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_17 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [1]),
        .I4(fch_pc1[1]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_3 
       (.I0(\rgf/treg/tr [1]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [1]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_6 
       (.I0(\rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_18_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_19_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_20_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_21_n_0 ),
        .I5(\rgf/b1bus_sr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_19 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [2]),
        .I4(fch_pc1[2]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_3 
       (.I0(\rgf/treg/tr [2]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [2]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_6 
       (.I0(\rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_23_n_0 ),
        .I5(\rgf/b1bus_sr [2]),
        .O(\rgf/b1bus_out/niss_dsp_b1[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_5 
       (.I0(\rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_9_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_10_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_11_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_12_n_0 ),
        .I5(\rgf/b1bus_sr [3]),
        .O(\rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_7 
       (.I0(\rgf/treg/tr [3]),
        .I1(\rgf/b1bus_sel_cr [4]),
        .I2(\rgf/ivec/iv [3]),
        .I3(\rgf/b1bus_sel_cr [3]),
        .O(\rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_8 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [3]),
        .I4(fch_pc1[3]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_10 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [5]),
        .I4(fch_pc1[5]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_5 
       (.I0(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_10_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_11_n_0 ),
        .I2(\rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_12_n_0 ),
        .I3(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_13_n_0 ),
        .I4(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_14_n_0 ),
        .I5(\rgf/b1bus_sr [5]),
        .O(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000AC000)) 
    \rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_7 
       (.I0(\rgf/treg/tr [5]),
        .I1(\rgf/ivec/iv [5]),
        .I2(ctl_selb1_rn[1]),
        .I3(ctl_selb1_rn[0]),
        .I4(ctl_selb1_rn[2]),
        .I5(\niss_dsp_b1[5]_INST_0_i_25_n_0 ),
        .O(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_3 
       (.I0(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_6_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_7_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [6]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [6]),
        .O(\rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_4 
       (.I0(\rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_9_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_10_n_0 ),
        .I3(\rgf/sreg/sr [6]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_8 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [6]),
        .I4(fch_pc1[6]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[6]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_3 
       (.I0(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_6_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_7_n_0 ),
        .I2(\rgf/b1bus_sel_cr [3]),
        .I3(\rgf/ivec/iv [7]),
        .I4(\rgf/b1bus_sel_cr [4]),
        .I5(\rgf/treg/tr [7]),
        .O(\rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_4 
       (.I0(\rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_8_n_0 ),
        .I1(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_9_n_0 ),
        .I2(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_10_n_0 ),
        .I3(\rgf/sreg/sr [7]),
        .I4(\rgf/b1bus_sel_cr [0]),
        .O(\rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_8 
       (.I0(\rgf/b1bus_sel_cr [5]),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/b1bus_sel_cr [2]),
        .I3(\rgf/sptr/sp [7]),
        .I4(fch_pc1[7]),
        .I5(\rgf/b1bus_sel_cr [1]),
        .O(\rgf/b1bus_out/niss_dsp_b1[7]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/b1bus_out/rgf_c1bus_wb[31]_i_68 
       (.I0(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_79_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_18_n_0 ),
        .I3(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_17_n_0 ),
        .I4(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_16_n_0 ),
        .I5(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_7_n_0 ),
        .O(\rgf/b1bus_out/rgf_c1bus_wb[31]_i_68_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_26 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_27 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_28 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_29 
       (.I0(\rgf/bank02/gr04 [0]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [0]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[0]_INST_0_i_8 
       (.I0(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_27_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_28_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[0]_INST_0_i_29_n_0 ),
        .O(\rgf/bank02/p_1_in [0]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [10]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [10]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[10]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [10]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [10]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[10]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [11]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [11]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[11]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [11]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [11]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[11]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_1_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [12]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [12]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[12]_INST_0_i_33 
       (.I0(\rgf/bank02/gr04 [12]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [12]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[12]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_32_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_33_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_34_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_35_n_0 ),
        .O(\rgf/bank02/p_1_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_32 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_33 
       (.I0(\rgf/bank02/gr00 [13]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [13]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_34 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[13]_INST_0_i_35 
       (.I0(\rgf/bank02/gr04 [13]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [13]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[13]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_25 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_26 
       (.I0(\rgf/bank02/gr00 [14]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [14]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_27 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_28 
       (.I0(\rgf/bank02/gr04 [14]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [14]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[14]_INST_0_i_8 
       (.I0(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_27_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[14]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/p_1_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [15]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [15]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_33 
       (.I0(\rgf/bank02/gr04 [15]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [15]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_81 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso/gr6_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_82 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso/gr5_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_83 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_84 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[15]_INST_0_i_129_n_0 ),
        .I4(\badr[31]_INST_0_i_81_n_0 ),
        .O(\bank02/a0buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_85 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso/gr2_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_86 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso/gr1_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_87 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_81_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso/gr4_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_88 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[15]_INST_0_i_9 
       (.I0(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[15]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_1_in [15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_25 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_26 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_27 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_28 
       (.I0(\rgf/bank02/gr04 [1]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [1]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[1]_INST_0_i_8 
       (.I0(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_27_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[1]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/p_1_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_25 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_26 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_27 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_28 
       (.I0(\rgf/bank02/gr04 [2]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [2]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[2]_INST_0_i_8 
       (.I0(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_27_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[2]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/p_1_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_25 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_26 
       (.I0(\rgf/bank02/gr00 [3]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [3]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_27 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_28 
       (.I0(\rgf/bank02/gr04 [3]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [3]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[3]_INST_0_i_8 
       (.I0(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_27_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[3]_INST_0_i_28_n_0 ),
        .O(\rgf/bank02/p_1_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_26 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_27 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_28 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_29 
       (.I0(\rgf/bank02/gr04 [4]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [4]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[4]_INST_0_i_8 
       (.I0(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_27_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_28_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[4]_INST_0_i_29_n_0 ),
        .O(\rgf/bank02/p_1_in [4]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [5]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [5]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[5]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [5]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [5]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[5]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [6]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [6]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[6]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [6]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [6]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[6]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [7]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [7]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[7]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [7]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [7]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[7]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_1_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [8]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [8]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[8]_INST_0_i_33 
       (.I0(\rgf/bank02/gr04 [8]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [8]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_29 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/a0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/a0buso/gr5_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_30 
       (.I0(\rgf/bank02/gr00 [9]),
        .I1(\bank02/a0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [9]),
        .I3(\bank02/a0buso/gr7_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_31 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/a0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/a0buso/gr1_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso/i_/badr[9]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [9]),
        .I1(\bank02/a0buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [9]),
        .I3(\bank02/a0buso/gr3_bus1 ),
        .O(\rgf/bank02/a0buso/i_/badr[9]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [0]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [0]),
        .I4(\badr[16]_INST_0_i_22_n_0 ),
        .I5(\badr[16]_INST_0_i_23_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [0]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [0]),
        .I4(\badr[16]_INST_0_i_24_n_0 ),
        .I5(\badr[16]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[16]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [1]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [1]),
        .I4(\badr[17]_INST_0_i_21_n_0 ),
        .I5(\badr[17]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [1]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [1]),
        .I4(\badr[17]_INST_0_i_23_n_0 ),
        .I5(\badr[17]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[17]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [2]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [2]),
        .I4(\badr[18]_INST_0_i_21_n_0 ),
        .I5(\badr[18]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [2]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [2]),
        .I4(\badr[18]_INST_0_i_23_n_0 ),
        .I5(\badr[18]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[18]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [3]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [3]),
        .I4(\badr[19]_INST_0_i_21_n_0 ),
        .I5(\badr[19]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [3]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [3]),
        .I4(\badr[19]_INST_0_i_23_n_0 ),
        .I5(\badr[19]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[19]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [4]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [4]),
        .I4(\badr[20]_INST_0_i_22_n_0 ),
        .I5(\badr[20]_INST_0_i_23_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [4]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [4]),
        .I4(\badr[20]_INST_0_i_24_n_0 ),
        .I5(\badr[20]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[20]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [5]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [5]),
        .I4(\badr[21]_INST_0_i_21_n_0 ),
        .I5(\badr[21]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [5]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [5]),
        .I4(\badr[21]_INST_0_i_23_n_0 ),
        .I5(\badr[21]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[21]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [6]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [6]),
        .I4(\badr[22]_INST_0_i_21_n_0 ),
        .I5(\badr[22]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [6]),
        .I4(\badr[22]_INST_0_i_23_n_0 ),
        .I5(\badr[22]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[22]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [7]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [7]),
        .I4(\badr[23]_INST_0_i_21_n_0 ),
        .I5(\badr[23]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [7]),
        .I4(\badr[23]_INST_0_i_23_n_0 ),
        .I5(\badr[23]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[23]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [8]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [8]),
        .I4(\badr[24]_INST_0_i_22_n_0 ),
        .I5(\badr[24]_INST_0_i_23_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [8]),
        .I4(\badr[24]_INST_0_i_24_n_0 ),
        .I5(\badr[24]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[24]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [9]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [9]),
        .I4(\badr[25]_INST_0_i_21_n_0 ),
        .I5(\badr[25]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [9]),
        .I4(\badr[25]_INST_0_i_23_n_0 ),
        .I5(\badr[25]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[25]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [10]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [10]),
        .I4(\badr[26]_INST_0_i_21_n_0 ),
        .I5(\badr[26]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [10]),
        .I4(\badr[26]_INST_0_i_23_n_0 ),
        .I5(\badr[26]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[26]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [11]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [11]),
        .I4(\badr[27]_INST_0_i_21_n_0 ),
        .I5(\badr[27]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [11]),
        .I4(\badr[27]_INST_0_i_23_n_0 ),
        .I5(\badr[27]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[27]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [12]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [12]),
        .I4(\badr[28]_INST_0_i_22_n_0 ),
        .I5(\badr[28]_INST_0_i_23_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [12]),
        .I4(\badr[28]_INST_0_i_24_n_0 ),
        .I5(\badr[28]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[28]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [13]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [13]),
        .I4(\badr[29]_INST_0_i_21_n_0 ),
        .I5(\badr[29]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [13]),
        .I4(\badr[29]_INST_0_i_23_n_0 ),
        .I5(\badr[29]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[29]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_10 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [14]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [14]),
        .I4(\badr[30]_INST_0_i_21_n_0 ),
        .I5(\badr[30]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_11 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\badr[30]_INST_0_i_23_n_0 ),
        .I5(\badr[30]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[30]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_12 
       (.I0(\bank02/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [15]),
        .I2(\bank02/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [15]),
        .I4(\badr[31]_INST_0_i_43_n_0 ),
        .I5(\badr[31]_INST_0_i_44_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_13 
       (.I0(\bank02/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\badr[31]_INST_0_i_47_n_0 ),
        .I5(\badr[31]_INST_0_i_48_n_0 ),
        .O(\rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_41 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_80_n_0 ),
        .I4(\badr[31]_INST_0_i_39_n_0 ),
        .O(\bank02/a0buso2h/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_42 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[31]_INST_0_i_80_n_0 ),
        .O(\bank02/a0buso2h/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_45 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_39_n_0 ),
        .I4(\badr[31]_INST_0_i_80_n_0 ),
        .O(\bank02/a0buso2h/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a0buso2h/i_/badr[31]_INST_0_i_46 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_39_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_80_n_0 ),
        .O(\bank02/a0buso2h/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_30 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_31 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_32 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_33 
       (.I0(\rgf/bank02/gr24 [0]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [0]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_9 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[0]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_0_in [0]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [10]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [10]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [10]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [10]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [11]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [11]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [11]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [11]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/p_0_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_34 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [12]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [12]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [12]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [12]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[12]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_36_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_37_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_38_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/p_0_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_36 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_37 
       (.I0(\rgf/bank02/gr20 [13]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [13]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_38 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_39 
       (.I0(\rgf/bank02/gr24 [13]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [13]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[13]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_30 
       (.I0(\rgf/bank02/gr20 [14]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [14]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_31 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_32 
       (.I0(\rgf/bank02/gr24 [14]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [14]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_9 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[14]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_0_in [14]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_10 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/p_0_in [15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_34 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [15]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [15]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [15]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [15]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_89 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso2l/gr6_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_90 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_81_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_58_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso2l/gr5_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_91 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso2l/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_92 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[15]_INST_0_i_129_n_0 ),
        .I4(\badr[31]_INST_0_i_81_n_0 ),
        .O(\bank02/a0buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_93 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_57_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso2l/gr2_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_94 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso2l/gr1_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_95 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_81_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso2l/gr4_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a0buso2l/i_/badr[15]_INST_0_i_96 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[15]_INST_0_i_129_n_0 ),
        .O(\bank02/a0buso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_30 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_31 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_32 
       (.I0(\rgf/bank02/gr24 [1]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [1]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_9 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[1]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_0_in [1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_30 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_31 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_32 
       (.I0(\rgf/bank02/gr24 [2]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [2]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_9 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[2]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_0_in [2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_30 
       (.I0(\rgf/bank02/gr20 [3]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [3]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_31 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_32 
       (.I0(\rgf/bank02/gr24 [3]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [3]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_9 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_30_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_31_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[3]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_0_in [3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_30 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_31 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_32 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_33 
       (.I0(\rgf/bank02/gr24 [4]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [4]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_9 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[4]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/p_0_in [4]));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [5]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [5]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [5]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [5]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[5]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [6]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [6]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [6]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [6]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[6]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [7]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [7]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [7]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [7]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[7]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/p_0_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_34 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [8]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [8]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [8]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [8]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[8]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_11 
       (.I0(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_0_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_34 
       (.I0(\rgf/bank02/gr20 [9]),
        .I1(\bank02/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [9]),
        .I3(\bank02/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_35 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\bank02/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\bank02/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_36 
       (.I0(\rgf/bank02/gr24 [9]),
        .I1(\bank02/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [9]),
        .I3(\bank02/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a0buso2l/i_/badr[9]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_13 
       (.I0(\bank02/a1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [0]),
        .I2(\bank02/a1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [0]),
        .I4(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_14 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso/i_/badr[0]_INST_0_i_40 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\rgf/bank02/gr01 [0]),
        .I2(\rgf/bank_sel [0]),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [10]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [10]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [10]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [10]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[10]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [10]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[10]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[10]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [11]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [11]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [11]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [11]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[11]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [11]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[11]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[11]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [12]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [12]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [12]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [12]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[12]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [12]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[12]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[12]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_16 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_17 
       (.I0(\rgf/bank02/gr00 [13]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [13]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_18 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso/gr2_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_20 
       (.I0(\rgf/bank02/gr04 [13]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [13]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[13]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_16_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/gr02 [13]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[13]_INST_0_i_19_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[13]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_13 
       (.I0(\bank02/a1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [14]),
        .I2(\bank02/a1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [14]),
        .I4(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_14 
       (.I0(\rgf/bank02/gr00 [14]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [14]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso/i_/badr[14]_INST_0_i_39 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\rgf/bank02/gr01 [14]),
        .I2(\rgf/bank_sel [0]),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_16 
       (.I0(\bank02/a1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [15]),
        .I2(\bank02/a1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [15]),
        .I4(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_55_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_17 
       (.I0(\rgf/bank02/gr00 [15]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [15]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_18 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_53 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_54 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[31]_INST_0_i_19_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_55 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\rgf/bank02/gr01 [15]),
        .I2(\rgf/bank_sel [0]),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_55_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_56 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_57 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_67_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .O(\bank02/a1buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_58 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso/gr6_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a1buso/i_/badr[15]_INST_0_i_59 
       (.I0(\rgf/bank_sel [0]),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso/gr5_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_13 
       (.I0(\bank02/a1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [1]),
        .I2(\bank02/a1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [1]),
        .I4(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_14 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso/i_/badr[1]_INST_0_i_39 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\rgf/bank02/gr01 [1]),
        .I2(\rgf/bank_sel [0]),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_13 
       (.I0(\bank02/a1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [2]),
        .I2(\bank02/a1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [2]),
        .I4(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_14 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso/i_/badr[2]_INST_0_i_39 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\rgf/bank02/gr01 [2]),
        .I2(\rgf/bank_sel [0]),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_13 
       (.I0(\bank02/a1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [3]),
        .I2(\bank02/a1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [3]),
        .I4(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_14 
       (.I0(\rgf/bank02/gr00 [3]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [3]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso/i_/badr[3]_INST_0_i_39 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\rgf/bank02/gr01 [3]),
        .I2(\rgf/bank_sel [0]),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_13 
       (.I0(\bank02/a1buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [4]),
        .I2(\bank02/a1buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [4]),
        .I4(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_14 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso/i_/badr[4]_INST_0_i_40 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\rgf/bank02/gr01 [4]),
        .I2(\rgf/bank_sel [0]),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [5]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [5]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [5]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [5]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[5]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [5]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[5]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[5]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [6]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [6]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [6]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [6]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[6]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [6]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[6]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[6]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [7]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [7]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [7]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [7]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[7]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [7]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[7]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[7]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [8]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [8]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [8]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [8]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[8]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [8]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[8]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[8]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_15 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/a1buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/a1buso/gr5_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_16 
       (.I0(\rgf/bank02/gr00 [9]),
        .I1(\bank02/a1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [9]),
        .I3(\bank02/a1buso/gr7_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_18 
       (.I0(\rgf/bank02/gr04 [9]),
        .I1(\bank02/a1buso/gr4_bus1 ),
        .I2(\rgf/bank02/gr03 [9]),
        .I3(\bank02/a1buso/gr3_bus1 ),
        .O(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso/i_/badr[9]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_16_n_0 ),
        .I2(\rgf/bank02/gr02 [9]),
        .I3(\bank02/a1buso/gr2_bus1 ),
        .I4(\badr[9]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso/i_/badr[9]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/p_1_in1_in [9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso/i_/rgf_c1bus_wb[10]_i_34 
       (.I0(\bank02/a1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [14]),
        .I2(\bank02/a1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [14]),
        .I4(\rgf_c1bus_wb[10]_i_37_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_38_n_0 ),
        .O(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[10]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_53 
       (.I0(\bank02/a1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [15]),
        .I2(\bank02/a1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [15]),
        .I4(\rgf_c1bus_wb[28]_i_69_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_70_n_0 ),
        .O(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_55 
       (.I0(\bank02/a1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [2]),
        .I2(\bank02/a1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [2]),
        .I4(\rgf_c1bus_wb[28]_i_73_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_74_n_0 ),
        .O(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_58 
       (.I0(\bank02/a1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [1]),
        .I2(\bank02/a1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [1]),
        .I4(\rgf_c1bus_wb[28]_i_77_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_78_n_0 ),
        .O(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_62 
       (.I0(\bank02/a1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [4]),
        .I2(\bank02/a1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [4]),
        .I4(\rgf_c1bus_wb[28]_i_83_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_84_n_0 ),
        .O(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_65 
       (.I0(\bank02/a1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [3]),
        .I2(\bank02/a1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [3]),
        .I4(\rgf_c1bus_wb[28]_i_87_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_88_n_0 ),
        .O(\rgf/bank02/a1buso/i_/rgf_c1bus_wb[28]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\rgf/bank02/gr21 [0]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [0]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [0]),
        .I4(\badr[16]_INST_0_i_15_n_0 ),
        .I5(\badr[16]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [0]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [0]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[16]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\rgf/bank02/gr21 [1]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [1]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [1]),
        .I4(\badr[17]_INST_0_i_15_n_0 ),
        .I5(\badr[17]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [1]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [1]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[17]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\rgf/bank02/gr21 [2]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [2]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [2]),
        .I4(\badr[18]_INST_0_i_15_n_0 ),
        .I5(\badr[18]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [2]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [2]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[18]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\rgf/bank02/gr21 [3]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [3]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [3]),
        .I4(\badr[19]_INST_0_i_15_n_0 ),
        .I5(\badr[19]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [3]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [3]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[19]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\rgf/bank02/gr21 [4]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [4]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [4]),
        .I4(\badr[20]_INST_0_i_15_n_0 ),
        .I5(\badr[20]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [4]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [4]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[20]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\rgf/bank02/gr21 [5]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [5]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [5]),
        .I4(\badr[21]_INST_0_i_15_n_0 ),
        .I5(\badr[21]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [5]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [5]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[21]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\rgf/bank02/gr21 [6]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [6]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [6]),
        .I4(\badr[22]_INST_0_i_15_n_0 ),
        .I5(\badr[22]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [6]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[22]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\rgf/bank02/gr21 [7]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [7]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [7]),
        .I4(\badr[23]_INST_0_i_15_n_0 ),
        .I5(\badr[23]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [7]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[23]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\rgf/bank02/gr21 [8]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [8]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [8]),
        .I4(\badr[24]_INST_0_i_15_n_0 ),
        .I5(\badr[24]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [8]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[24]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\rgf/bank02/gr21 [9]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [9]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [9]),
        .I4(\badr[25]_INST_0_i_15_n_0 ),
        .I5(\badr[25]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [9]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[25]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\rgf/bank02/gr21 [10]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [10]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [10]),
        .I4(\badr[26]_INST_0_i_15_n_0 ),
        .I5(\badr[26]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [10]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[26]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\rgf/bank02/gr21 [11]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [11]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [11]),
        .I4(\badr[27]_INST_0_i_15_n_0 ),
        .I5(\badr[27]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [11]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[27]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\rgf/bank02/gr21 [12]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [12]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [12]),
        .I4(\badr[28]_INST_0_i_15_n_0 ),
        .I5(\badr[28]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [12]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[28]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\rgf/bank02/gr21 [13]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [13]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [13]),
        .I4(\badr[29]_INST_0_i_15_n_0 ),
        .I5(\badr[29]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [13]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[29]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\rgf/bank02/gr21 [14]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_4 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [14]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [14]),
        .I4(\badr[30]_INST_0_i_15_n_0 ),
        .I5(\badr[30]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_5 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[30]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_21 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_67_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .O(\bank02/a1buso2h/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_22 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2h/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_25 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2h/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_26 
       (.I0(\rgf/bank02/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[31]_INST_0_i_19_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2h/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_27 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\rgf/bank02/gr21 [15]),
        .I2(\rgf/bank02/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_6 
       (.I0(\bank02/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [15]),
        .I2(\bank02/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [15]),
        .I4(\badr[31]_INST_0_i_23_n_0 ),
        .I5(\badr[31]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_7 
       (.I0(\bank02/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_27_n_0 ),
        .O(\rgf/bank02/a1buso2h/i_/badr[31]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_16 
       (.I0(\bank02/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [0]),
        .I2(\bank02/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [0]),
        .I4(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_17 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_18 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_41 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\rgf/bank02/gr21 [0]),
        .I2(\badr[13]_INST_0_i_46_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [10]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [10]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [10]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [10]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [10]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[10]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[10]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [11]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [11]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [11]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [11]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [11]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[11]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[11]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [12]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [12]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [12]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [12]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [12]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[12]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[12]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_21 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_22 
       (.I0(\rgf/bank02/gr20 [13]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [13]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_23 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2l/gr2_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_25 
       (.I0(\rgf/bank02/gr24 [13]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [13]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_22_n_0 ),
        .I2(\rgf/bank02/gr22 [13]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[13]_INST_0_i_24_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[13]_INST_0_i_25_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [13]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_16 
       (.I0(\bank02/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_17 
       (.I0(\rgf/bank02/gr20 [14]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [14]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_18 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_40 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\rgf/bank02/gr21 [14]),
        .I2(\badr[13]_INST_0_i_46_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_19 
       (.I0(\bank02/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_62_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [15]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [15]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_21 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_60 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2l/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_61 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[31]_INST_0_i_19_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_62 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\rgf/bank02/gr21 [15]),
        .I2(\badr[13]_INST_0_i_46_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_62_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_63 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2l/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_64 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_67_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .O(\bank02/a1buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_65 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2l/gr6_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_66 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank02/a1buso2l/gr5_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_16 
       (.I0(\bank02/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [1]),
        .I2(\bank02/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [1]),
        .I4(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_17 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_18 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_40 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\rgf/bank02/gr21 [1]),
        .I2(\badr[13]_INST_0_i_46_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_16 
       (.I0(\bank02/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [2]),
        .I2(\bank02/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [2]),
        .I4(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_17 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_18 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_40 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\rgf/bank02/gr21 [2]),
        .I2(\badr[13]_INST_0_i_46_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_16 
       (.I0(\bank02/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [3]),
        .I2(\bank02/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [3]),
        .I4(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_17 
       (.I0(\rgf/bank02/gr20 [3]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [3]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_18 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_40 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\rgf/bank02/gr21 [3]),
        .I2(\badr[13]_INST_0_i_46_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_16 
       (.I0(\bank02/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [4]),
        .I2(\bank02/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [4]),
        .I4(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_17 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_18 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_41 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\rgf/bank02/gr21 [4]),
        .I2(\badr[13]_INST_0_i_46_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [5]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [5]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [5]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [5]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [5]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[5]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[5]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [6]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [6]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [6]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [6]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [6]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[6]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[6]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [7]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [7]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [7]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [7]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [7]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[7]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[7]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [8]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [8]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [8]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [8]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [8]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[8]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[8]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_19 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_20 
       (.I0(\rgf/bank02/gr20 [9]),
        .I1(\bank02/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [9]),
        .I3(\bank02/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_22 
       (.I0(\rgf/bank02/gr24 [9]),
        .I1(\bank02/a1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr23 [9]),
        .I3(\bank02/a1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEEE)) 
    \rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_5 
       (.I0(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank02/gr22 [9]),
        .I3(\bank02/a1buso2l/gr2_bus1 ),
        .I4(\badr[9]_INST_0_i_21_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[9]_INST_0_i_22_n_0 ),
        .O(\rgf/bank02/p_0_in0_in [9]));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_10 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [5]),
        .O(\bank02/b0buso/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/b0buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/b0buso/gr7_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_12 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_23_n_0 ),
        .I1(\bank02/b0buso/gr1_bus1 ),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\bank02/b0buso/gr2_bus1 ),
        .I4(\rgf/bank02/gr02 [0]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_23 
       (.I0(\rgf/bank02/gr04 [0]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr03 [0]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_4 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_11_n_0 ),
        .I5(\rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [0]));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bbus_o[0]_INST_0_i_9 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .O(\bank02/b0buso/gr6_bus1 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_19_n_0 ),
        .I1(\bank02/b0buso/gr1_bus1 ),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\bank02/b0buso/gr2_bus1 ),
        .I4(\rgf/bank02/gr02 [1]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_18 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr05 [1]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_19 
       (.I0(\rgf/bank02/gr04 [1]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr03 [1]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9 
       (.I0(\bank02/b0buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [1]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [1]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[1]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_19_n_0 ),
        .I1(\bank02/b0buso/gr1_bus1 ),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\bank02/b0buso/gr2_bus1 ),
        .I4(\rgf/bank02/gr02 [2]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_18 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr05 [2]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_19 
       (.I0(\rgf/bank02/gr04 [2]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr03 [2]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9 
       (.I0(\bank02/b0buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [2]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [2]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[2]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10 
       (.I0(\bank02/b0buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [3]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [3]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_20_n_0 ),
        .I1(\bank02/b0buso/gr1_bus1 ),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\bank02/b0buso/gr2_bus1 ),
        .I4(\rgf/bank02/gr02 [3]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_19 
       (.I0(\rgf/bank02/gr06 [3]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr05 [3]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_20 
       (.I0(\rgf/bank02/gr04 [3]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr03 [3]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[3]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_19_n_0 ),
        .I1(\bank02/b0buso/gr1_bus1 ),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\bank02/b0buso/gr2_bus1 ),
        .I4(\rgf/bank02/gr02 [4]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_18 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr05 [4]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_19 
       (.I0(\rgf/bank02/gr04 [4]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr03 [4]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9 
       (.I0(\bank02/b0buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [4]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [4]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[4]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_16 
       (.I0(\bank02/b0buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [5]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [5]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_31_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_17 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_32_n_0 ),
        .I1(\bank02/b0buso/gr1_bus1 ),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\bank02/b0buso/gr2_bus1 ),
        .I4(\rgf/bank02/gr02 [5]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_31 
       (.I0(\rgf/bank02/gr06 [5]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr05 [5]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_32 
       (.I0(\rgf/bank02/gr04 [5]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr03 [5]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_33 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [1]),
        .O(\bank02/b0buso/gr1_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bbus_o[5]_INST_0_i_34 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .O(\bank02/b0buso/gr2_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_13 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [6]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_14 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [6]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [6]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_20 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_7 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/gr00 [6]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [6]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bbus_o[6]_INST_0_i_14_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_13 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [7]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_14 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [7]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [7]),
        .I4(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_20 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_7 
       (.I0(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/gr00 [7]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [7]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bbus_o[7]_INST_0_i_14_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_21 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank02/gr00 [10]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [10]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_35 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [10]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_36 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [10]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [10]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_46 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[10]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_21 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank02/gr00 [11]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [11]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_35 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [11]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_36 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [11]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [11]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_46_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_46 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[11]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_25 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_54_n_0 ),
        .I1(\rgf/bank02/gr00 [12]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [12]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_55_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_54 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [12]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_54_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_55 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [12]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [12]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_73_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_73 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[12]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_16 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/gr00 [13]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [13]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_31_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [13]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_31 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [13]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [13]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_41 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[13]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_17 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/gr00 [14]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [14]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_31 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [14]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_32 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [14]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [14]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_42_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_42 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[14]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_24 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_50_n_0 ),
        .I1(\rgf/bank02/gr00 [15]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [15]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_53_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_50 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [15]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_51 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .O(\bank02/b0buso/gr0_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_52 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [7]),
        .O(\bank02/b0buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_53 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [15]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [15]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_79_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_77 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [3]),
        .O(\bank02/b0buso/gr3_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_78 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .O(\bank02/b0buso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_79 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[15]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_17 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/gr00 [8]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [8]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_34_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_33 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [8]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_34 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [8]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [8]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_44_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_44 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[8]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_19 
       (.I0(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/gr00 [9]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr07 [9]),
        .I4(\bank02/b0buso/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_34_n_0 ),
        .O(\rgf/bank02/p_1_in3_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_33 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\bank02/b0buso/gr6_bus1 ),
        .I2(\rgf/bank02/gr05 [9]),
        .I3(\bank02/b0buso/gr5_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_34 
       (.I0(\bank02/b0buso/gr3_bus1 ),
        .I1(\rgf/bank02/gr03 [9]),
        .I2(\bank02/b0buso/gr4_bus1 ),
        .I3(\rgf/bank02/gr04 [9]),
        .I4(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_44_n_0 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_44 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/b0buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/b0buso/gr1_bus1 ),
        .O(\rgf/bank02/b0buso/i_/bdatw[9]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_81 
       (.I0(\bank02/b0buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [0]),
        .I2(\bank02/b0buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [0]),
        .I4(\rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_84_n_0 ),
        .O(\rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_81_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_84 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr05 [0]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso/i_/rgf_c0bus_wb[31]_i_84_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_13 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .O(\bank02/b0buso2l/gr6_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_14 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [5]),
        .O(\bank02/b0buso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_15 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/b0buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/b0buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_16 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_24_n_0 ),
        .I1(\bank02/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\bank02/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank02/gr22 [0]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_24 
       (.I0(\rgf/bank02/gr24 [0]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr23 [0]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_5 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_15_n_0 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[0]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [0]));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_16 
       (.I0(\rgf/bank02/gr26 [1]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr25 [1]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_17 
       (.I0(\rgf/bank02/gr24 [1]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr23 [1]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_7 
       (.I0(\bank02/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [1]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [1]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_8 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_17_n_0 ),
        .I1(\bank02/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\bank02/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank02/gr22 [1]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[1]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_16 
       (.I0(\rgf/bank02/gr26 [2]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr25 [2]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_17 
       (.I0(\rgf/bank02/gr24 [2]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr23 [2]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_7 
       (.I0(\bank02/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [2]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [2]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_8 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_17_n_0 ),
        .I1(\bank02/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\bank02/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank02/gr22 [2]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[2]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_17 
       (.I0(\rgf/bank02/gr26 [3]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr25 [3]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_18 
       (.I0(\rgf/bank02/gr24 [3]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr23 [3]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_8 
       (.I0(\bank02/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [3]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [3]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_17_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_9 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_18_n_0 ),
        .I1(\bank02/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\bank02/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank02/gr22 [3]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[3]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_16 
       (.I0(\rgf/bank02/gr26 [4]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr25 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_17 
       (.I0(\rgf/bank02/gr24 [4]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr23 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_7 
       (.I0(\bank02/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [4]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [4]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_8 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_17_n_0 ),
        .I1(\bank02/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\bank02/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank02/gr22 [4]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[4]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_14 
       (.I0(\bank02/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [5]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [5]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_27_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_15 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_28_n_0 ),
        .I1(\bank02/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\bank02/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank02/gr22 [5]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_27 
       (.I0(\rgf/bank02/gr26 [5]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr25 [5]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_28 
       (.I0(\rgf/bank02/gr24 [5]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank02/gr23 [5]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_29 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [1]),
        .O(\bank02/b0buso2l/gr1_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[5]_INST_0_i_30 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .O(\bank02/b0buso2l/gr2_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [6]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [6]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_19 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_6 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/gr20 [6]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [6]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[6]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [7]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [7]),
        .I4(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_19 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_6 
       (.I0(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/gr20 [7]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [7]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bbus_o[7]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_20 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/gr20 [10]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [10]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_34_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [10]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_34 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [10]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_45 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[10]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_20 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank02/gr20 [11]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [11]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_34_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_33 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [11]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_34 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [11]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_45 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[11]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_24 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_52_n_0 ),
        .I1(\rgf/bank02/gr20 [12]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [12]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_53_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_52 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [12]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_53 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [12]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_72_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_53_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_72 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[12]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_15 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_28_n_0 ),
        .I1(\rgf/bank02/gr20 [13]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [13]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_29_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_28 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [13]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_29 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [13]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_40 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[13]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_16 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/gr20 [14]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [14]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_30_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [14]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_30 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [14]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_41_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_41 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[14]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_23 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_46_n_0 ),
        .I1(\rgf/bank02/gr20 [15]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [15]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_49_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_46 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [15]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_47 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .O(\bank02/b0buso2l/gr0_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_48 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [7]),
        .O(\bank02/b0buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_49 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [15]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_76_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_74 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [3]),
        .O(\bank02/b0buso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_75 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .O(\bank02/b0buso2l/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_76 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[15]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_16 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/gr20 [8]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [8]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_31 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [8]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_32 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [8]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_43_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_43 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[8]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_18 
       (.I0(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/gr20 [9]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [9]),
        .I4(\bank02/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_32_n_0 ),
        .O(\rgf/bank02/p_0_in2_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_31 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\bank02/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank02/gr25 [9]),
        .I3(\bank02/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_32 
       (.I0(\bank02/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\bank02/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank02/gr24 [9]),
        .I4(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_43_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_43 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\bank02/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\bank02/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank02/b0buso2l/i_/bdatw[9]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_80 
       (.I0(\bank02/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank02/gr27 [0]),
        .I2(\bank02/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr20 [0]),
        .I4(\rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_83_n_0 ),
        .O(\rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_80_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_83 
       (.I0(\rgf/bank02/gr26 [0]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank02/gr25 [0]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank02/b0buso2l/i_/rgf_c0bus_wb[31]_i_83_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_18 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_32_n_0 ),
        .I2(\rgf/bank02/gr04 [10]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [10]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_31 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [10]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [10]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_44_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [10]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [10]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_44 
       (.I0(\rgf/bank02/gr06 [10]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [10]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[10]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_17 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_32_n_0 ),
        .I2(\rgf/bank02/gr04 [11]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [11]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_31 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [11]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [11]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_44_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [11]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [11]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_44 
       (.I0(\rgf/bank02/gr06 [11]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [11]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[11]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_30_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_31_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_32_n_0 ),
        .I3(\rgf/bank02/gr04 [4]),
        .I4(\bank02/b1buso/gr4_bus1 ),
        .I5(\bdatw[12]_INST_0_i_33_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_18 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_46_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_47_n_0 ),
        .I2(\rgf/bank02/gr04 [12]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [12]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_30 
       (.I0(\rgf/bank02/gr06 [4]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [4]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_31 
       (.I0(\rgf/bank02/gr00 [4]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [4]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_32 
       (.I0(\rgf/bank02/gr02 [4]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [4]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_46 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [12]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [12]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_69_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_47 
       (.I0(\rgf/bank02/gr02 [12]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [12]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_69 
       (.I0(\rgf/bank02/gr06 [12]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [12]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_11 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_23_n_0 ),
        .I2(\rgf/bank02/gr04 [13]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [13]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_22 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [13]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [13]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_23 
       (.I0(\rgf/bank02/gr02 [13]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [13]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_37 
       (.I0(\rgf/bank02/gr06 [13]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [13]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[13]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_15 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_27_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_28_n_0 ),
        .I2(\rgf/bank02/gr04 [14]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [14]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_27 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [14]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [14]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_28 
       (.I0(\rgf/bank02/gr02 [14]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [14]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_40 
       (.I0(\rgf/bank02/gr06 [14]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [14]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[14]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_20 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_43_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_44_n_0 ),
        .I2(\rgf/bank02/gr04 [15]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [15]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_43 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [15]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [15]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_71_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_44 
       (.I0(\rgf/bank02/gr02 [15]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [15]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_45 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso/gr3_bus1 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_71 
       (.I0(\rgf/bank02/gr06 [15]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [15]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_71_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_72 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b1bus_sel_0 [2]),
        .O(\bank02/b1buso/gr2_bus1 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b1buso/i_/bdatw[15]_INST_0_i_73 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b1bus_sel_0 [1]),
        .O(\bank02/b1buso/gr1_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_12 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank02/gr04 [8]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [8]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [8]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [8]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26 
       (.I0(\rgf/bank02/gr02 [8]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [8]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_40 
       (.I0(\rgf/bank02/gr06 [8]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [8]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[8]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_13 
       (.I0(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_26_n_0 ),
        .I2(\rgf/bank02/gr04 [9]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [9]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_25 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [9]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [9]),
        .I4(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_40_n_0 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_26 
       (.I0(\rgf/bank02/gr02 [9]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [9]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_40 
       (.I0(\rgf/bank02/gr06 [9]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [9]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/bdatw[9]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [0]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [0]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_11 
       (.I0(\rgf/bank02/gr02 [0]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [0]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_4 
       (.I0(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank02/gr04 [0]),
        .I4(\bank02/b1buso/gr4_bus1 ),
        .I5(\niss_dsp_b1[0]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_9 
       (.I0(\rgf/bank02/gr06 [0]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [0]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[0]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [1]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [1]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_11 
       (.I0(\rgf/bank02/gr02 [1]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [1]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_4 
       (.I0(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank02/gr04 [1]),
        .I4(\bank02/b1buso/gr4_bus1 ),
        .I5(\niss_dsp_b1[1]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_9 
       (.I0(\rgf/bank02/gr06 [1]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [1]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[1]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_10 
       (.I0(\rgf/bank02/gr00 [2]),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr07 [2]),
        .I3(\bank02/b1buso/gr7_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_11 
       (.I0(\rgf/bank02/gr02 [2]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [2]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_12 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b1bus_sel_0 [4]),
        .O(\bank02/b1buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_25 
       (.I0(\rgf/bank_sel [0]),
        .I1(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_26 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_0[1]),
        .I4(ctl_selb1_0[2]),
        .I5(ctl_selb1_rn[2]),
        .O(\bank02/b1buso/gr7_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFEFE)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_4 
       (.I0(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_9_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_10_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_11_n_0 ),
        .I3(\rgf/bank02/gr04 [2]),
        .I4(\bank02/b1buso/gr4_bus1 ),
        .I5(\niss_dsp_b1[2]_INST_0_i_13_n_0 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_9 
       (.I0(\rgf/bank02/gr06 [2]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [2]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[2]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_14 
       (.I0(\rgf/bank02/gr04 [3]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr03 [3]),
        .I4(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_15 
       (.I0(\rgf/bank02/gr02 [3]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [3]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_16 
       (.I0(\niss_dsp_b1[3]_INST_0_i_28_n_0 ),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr00 [3]),
        .I3(\niss_dsp_b1[3]_INST_0_i_29_n_0 ),
        .I4(\bank02/b1buso/gr6_bus1 ),
        .I5(\rgf/bank02/gr06 [3]),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_16 
       (.I0(\rgf/bank02/gr04 [5]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr03 [5]),
        .I4(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_17 
       (.I0(\rgf/bank02/gr02 [5]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr01 [5]),
        .I3(\rgf/bank_sel [0]),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_18 
       (.I0(\niss_dsp_b1[5]_INST_0_i_40_n_0 ),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr00 [5]),
        .I3(\niss_dsp_b1[5]_INST_0_i_42_n_0 ),
        .I4(\bank02/b1buso/gr6_bus1 ),
        .I5(\rgf/bank02/gr06 [5]),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_41 
       (.I0(\rgf/bank_sel [0]),
        .I1(\bdatw[15]_INST_0_i_63_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_43 
       (.I0(\rgf/bank_sel [0]),
        .I1(\niss_dsp_b1[5]_INST_0_i_62_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso/gr6_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_13 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [6]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [6]),
        .I4(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_14 
       (.I0(\rgf/bank02/gr02 [6]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [6]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_20 
       (.I0(\rgf/bank02/gr06 [6]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [6]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_7 
       (.I0(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/gr04 [6]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [6]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[6]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_13 
       (.I0(\bank02/b1buso/gr7_bus1 ),
        .I1(\rgf/bank02/gr07 [7]),
        .I2(\bank02/b1buso/gr0_bus1 ),
        .I3(\rgf/bank02/gr00 [7]),
        .I4(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_20_n_0 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_14 
       (.I0(\rgf/bank02/gr02 [7]),
        .I1(\bank02/b1buso/gr2_bus1 ),
        .I2(\rgf/bank02/gr01 [7]),
        .I3(\bank02/b1buso/gr1_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_20 
       (.I0(\rgf/bank02/gr06 [7]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr05 [7]),
        .I4(\bank02/b1buso/gr5_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_7 
       (.I0(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/gr04 [7]),
        .I3(\bank02/b1buso/gr4_bus1 ),
        .I4(\rgf/bank02/gr03 [7]),
        .I5(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/niss_dsp_b1[7]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_80 
       (.I0(\rgf/bank02/gr04 [4]),
        .I1(\rgf/bank_sel [0]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr03 [4]),
        .I4(\bank02/b1buso/gr3_bus1 ),
        .O(\rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_81 
       (.I0(\rgf_c1bus_wb[31]_i_87_n_0 ),
        .I1(\bank02/b1buso/gr0_bus1 ),
        .I2(\rgf/bank02/gr00 [4]),
        .I3(\rgf_c1bus_wb[31]_i_88_n_0 ),
        .I4(\bank02/b1buso/gr6_bus1 ),
        .I5(\rgf/bank02/gr06 [4]),
        .O(\rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_17 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/gr20 [10]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [10]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_30_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [10]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [10]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_30 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [10]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [10]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_43_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_43 
       (.I0(\rgf/bank02/gr22 [10]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [10]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[10]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_16 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank02/gr20 [11]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [11]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_30_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_29 
       (.I0(\rgf/bank02/gr26 [11]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [11]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_30 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [11]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [11]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43 
       (.I0(\rgf/bank02/gr22 [11]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [11]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[11]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14 
       (.I0(\bdatw[12]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank02/gr25 [4]),
        .I2(\bank02/b1buso2l/gr5_bus1 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_35_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_36_n_0 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_37_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_17 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_44_n_0 ),
        .I1(\rgf/bank02/gr20 [12]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [12]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_45_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_35 
       (.I0(\rgf/bank02/gr20 [4]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [4]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [4]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_37 
       (.I0(\rgf/bank02/gr24 [4]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr23 [4]),
        .I4(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_44 
       (.I0(\rgf/bank02/gr26 [12]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [12]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_45 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [12]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [12]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_68_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_68 
       (.I0(\rgf/bank02/gr22 [12]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [12]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_10 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_20_n_0 ),
        .I1(\rgf/bank02/gr20 [13]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [13]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_21_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_20 
       (.I0(\rgf/bank02/gr26 [13]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [13]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_21 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [13]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [13]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_36_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_36 
       (.I0(\rgf/bank02/gr22 [13]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [13]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[13]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank02/gr20 [14]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [14]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_26_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_25 
       (.I0(\rgf/bank02/gr26 [14]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [14]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_26 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [14]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [14]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_39 
       (.I0(\rgf/bank02/gr22 [14]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [14]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[14]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_19 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank02/gr20 [15]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [15]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_42_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_39 
       (.I0(\rgf/bank02/gr26 [15]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [15]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_40 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\bdatw[15]_INST_0_i_63_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_41 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_0[1]),
        .I4(ctl_selb1_0[2]),
        .I5(ctl_selb1_rn[2]),
        .O(\bank02/b1buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_42 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [15]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [15]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_70_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_70 
       (.I0(\rgf/bank02/gr22 [15]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [15]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_11 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank02/gr20 [8]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [8]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_23 
       (.I0(\rgf/bank02/gr26 [8]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [8]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_24 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [8]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [8]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39 
       (.I0(\rgf/bank02/gr22 [8]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [8]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[8]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_12 
       (.I0(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank02/gr20 [9]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [9]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23 
       (.I0(\rgf/bank02/gr26 [9]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [9]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [9]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [9]),
        .I5(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_39_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_39 
       (.I0(\rgf/bank02/gr22 [9]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [9]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/bdatw[9]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_14 
       (.I0(\rgf/bank02/gr20 [0]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [0]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_15 
       (.I0(\rgf/bank02/gr22 [0]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [0]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_16 
       (.I0(\rgf/bank02/gr24 [0]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr23 [0]),
        .I4(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_5 
       (.I0(\niss_dsp_b1[0]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/gr25 [0]),
        .I2(\bank02/b1buso2l/gr5_bus1 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_15_n_0 ),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_14 
       (.I0(\rgf/bank02/gr20 [1]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [1]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_15 
       (.I0(\rgf/bank02/gr22 [1]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [1]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_16 
       (.I0(\rgf/bank02/gr24 [1]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr23 [1]),
        .I4(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_5 
       (.I0(\niss_dsp_b1[1]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/gr25 [1]),
        .I2(\bank02/b1buso2l/gr5_bus1 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_14_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_15_n_0 ),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_16_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_15 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_16 
       (.I0(\rgf/bank02/gr20 [2]),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr27 [2]),
        .I3(\bank02/b1buso2l/gr7_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_17 
       (.I0(\rgf/bank02/gr22 [2]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [2]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_18 
       (.I0(\rgf/bank02/gr24 [2]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr23 [2]),
        .I4(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_5 
       (.I0(\niss_dsp_b1[2]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank02/gr25 [2]),
        .I2(\bank02/b1buso2l/gr5_bus1 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_18_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_17 
       (.I0(\rgf/bank02/gr24 [3]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr23 [3]),
        .I4(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_18 
       (.I0(\rgf/bank02/gr22 [3]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [3]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_19 
       (.I0(\niss_dsp_b1[3]_INST_0_i_30_n_0 ),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr20 [3]),
        .I3(\niss_dsp_b1[3]_INST_0_i_31_n_0 ),
        .I4(\bank02/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank02/gr26 [3]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_19 
       (.I0(\rgf/bank02/gr24 [5]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\rgf/bank02/gr23 [5]),
        .I4(\bank02/b1buso2l/gr3_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_20 
       (.I0(\rgf/bank02/gr22 [5]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [5]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_21 
       (.I0(\niss_dsp_b1[5]_INST_0_i_45_n_0 ),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr20 [5]),
        .I3(\niss_dsp_b1[5]_INST_0_i_46_n_0 ),
        .I4(\bank02/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank02/gr26 [5]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_44 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso2l/gr3_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_47 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_62_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso2l/gr6_bus1 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_11 
       (.I0(\rgf/bank02/gr26 [6]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [6]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_12 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [6]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [6]),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_19 
       (.I0(\rgf/bank02/gr22 [6]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [6]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_6 
       (.I0(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/gr20 [6]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [6]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_11 
       (.I0(\rgf/bank02/gr26 [7]),
        .I1(\badr[13]_INST_0_i_46_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank02/gr25 [7]),
        .I4(\bank02/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_12 
       (.I0(\bank02/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank02/gr23 [7]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/bank02/gr24 [7]),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_19_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_19 
       (.I0(\rgf/bank02/gr22 [7]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank02/gr21 [7]),
        .I3(\badr[13]_INST_0_i_46_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_6 
       (.I0(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_11_n_0 ),
        .I1(\rgf/bank02/gr20 [7]),
        .I2(\bank02/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank02/gr27 [7]),
        .I4(\bank02/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_12_n_0 ),
        .O(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_79 
       (.I0(\rgf_c1bus_wb[31]_i_83_n_0 ),
        .I1(\bank02/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank02/gr24 [5]),
        .I3(\rgf_c1bus_wb[31]_i_85_n_0 ),
        .I4(\bank02/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank02/gr22 [5]),
        .O(\rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_82 
       (.I0(\rgf_c1bus_wb[31]_i_89_n_0 ),
        .I1(\bank02/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank02/gr20 [4]),
        .I3(\rgf_c1bus_wb[31]_i_90_n_0 ),
        .I4(\bank02/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank02/gr26 [4]),
        .O(\rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_84 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_59_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_86 
       (.I0(\badr[13]_INST_0_i_46_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_61_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank02/b1buso2l/gr2_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/badr[0]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[0]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[0]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_b02 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/badr[14]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[14]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[14]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_b02 [14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/badr[15]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_16_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[15]_INST_0_i_18_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_20_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[15]_INST_0_i_21_n_0 ),
        .O(\rgf/a1bus_b02 [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/badr[1]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[1]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[1]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_b02 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/badr[2]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[2]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[2]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_b02 [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/badr[3]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[3]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[3]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_b02 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/badr[4]_INST_0_i_4 
       (.I0(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_13_n_0 ),
        .I1(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_14_n_0 ),
        .I2(\rgf/bank02/a1buso/i_/badr[4]_INST_0_i_15_n_0 ),
        .I3(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_16_n_0 ),
        .I4(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_17_n_0 ),
        .I5(\rgf/bank02/a1buso2l/i_/badr[4]_INST_0_i_18_n_0 ),
        .O(\rgf/a1bus_b02 [4]));
  FDRE \rgf/bank02/grn00/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [0]),
        .Q(\rgf/bank02/gr00 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [10]),
        .Q(\rgf/bank02/gr00 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [11]),
        .Q(\rgf/bank02/gr00 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [12]),
        .Q(\rgf/bank02/gr00 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [13]),
        .Q(\rgf/bank02/gr00 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [14]),
        .Q(\rgf/bank02/gr00 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [15]),
        .Q(\rgf/bank02/gr00 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [1]),
        .Q(\rgf/bank02/gr00 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [2]),
        .Q(\rgf/bank02/gr00 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [3]),
        .Q(\rgf/bank02/gr00 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [4]),
        .Q(\rgf/bank02/gr00 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [5]),
        .Q(\rgf/bank02/gr00 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [6]),
        .Q(\rgf/bank02/gr00 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [7]),
        .Q(\rgf/bank02/gr00 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [8]),
        .Q(\rgf/bank02/gr00 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn00/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__30_n_0 ),
        .D(\rgf/p_2_in [9]),
        .Q(\rgf/bank02/gr00 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[0]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[10]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[11]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[12]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[13]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[14]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[15]_i_2__0_n_0 ),
        .Q(\rgf/bank02/gr01 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[1]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[2]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[3]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[4]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[5]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[6]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[7]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[8]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn01/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__4_n_0 ),
        .D(\grn[9]_i_1__0_n_0 ),
        .Q(\rgf/bank02/gr01 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[0]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[10]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[11]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[12]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[13]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[14]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[15]_i_2__1_n_0 ),
        .Q(\rgf/bank02/gr02 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[1]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[2]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[3]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[4]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[5]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[6]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[7]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[8]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn02/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__3_n_0 ),
        .D(\grn[9]_i_1__1_n_0 ),
        .Q(\rgf/bank02/gr02 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[0]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[10]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[11]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[12]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[13]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[14]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[15]_i_2__2_n_0 ),
        .Q(\rgf/bank02/gr03 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[1]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[2]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[3]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[4]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[5]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[6]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[7]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[8]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn03/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__26_n_0 ),
        .D(\grn[9]_i_1__2_n_0 ),
        .Q(\rgf/bank02/gr03 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[0]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[10]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[11]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[12]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[13]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[14]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[15]_i_2__3_n_0 ),
        .Q(\rgf/bank02/gr04 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[1]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[2]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[3]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[4]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[5]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[6]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[7]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[8]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn04/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__2_n_0 ),
        .D(\grn[9]_i_1__3_n_0 ),
        .Q(\rgf/bank02/gr04 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[0]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[10]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[11]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[12]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[13]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[14]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[15]_i_2__4_n_0 ),
        .Q(\rgf/bank02/gr05 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[1]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[2]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[3]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[4]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[5]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[6]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[7]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[8]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn05/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__1_n_0 ),
        .D(\grn[9]_i_1__4_n_0 ),
        .Q(\rgf/bank02/gr05 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[0]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[10]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[11]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[12]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[13]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[14]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[15]_i_2__5_n_0 ),
        .Q(\rgf/bank02/gr06 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[1]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[2]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[3]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[4]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[5]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[6]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[7]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[8]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn06/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__0_n_0 ),
        .D(\grn[9]_i_1__5_n_0 ),
        .Q(\rgf/bank02/gr06 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[0]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[10]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[11]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[12]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[13]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[14]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[15]_i_2__6_n_0 ),
        .Q(\rgf/bank02/gr07 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[1]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[2]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[3]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[4]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[5]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[6]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[7]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[8]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn07/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1_n_0 ),
        .D(\grn[9]_i_1__6_n_0 ),
        .Q(\rgf/bank02/gr07 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[0]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[10]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[11]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[12]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[13]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[14]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[15]_i_2__15_n_0 ),
        .Q(\rgf/bank02/gr20 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[1]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[2]_i_1__30_n_0 ),
        .Q(\rgf/bank02/gr20 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[3]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[4]_i_1__30_n_0 ),
        .Q(\rgf/bank02/gr20 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[5]_i_1__30_n_0 ),
        .Q(\rgf/bank02/gr20 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[6]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[7]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[8]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn20/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__28_n_0 ),
        .D(\grn[9]_i_1__15_n_0 ),
        .Q(\rgf/bank02/gr20 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[0]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[10]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[11]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[12]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[13]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[14]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[15]_i_2__16_n_0 ),
        .Q(\rgf/bank02/gr21 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[1]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[2]_i_1__29_n_0 ),
        .Q(\rgf/bank02/gr21 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[3]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[4]_i_1__29_n_0 ),
        .Q(\rgf/bank02/gr21 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[5]_i_1__29_n_0 ),
        .Q(\rgf/bank02/gr21 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[6]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[7]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[8]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn21/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__16_n_0 ),
        .D(\grn[9]_i_1__16_n_0 ),
        .Q(\rgf/bank02/gr21 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[0]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[10]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[11]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[12]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[13]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[14]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[15]_i_2__17_n_0 ),
        .Q(\rgf/bank02/gr22 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[1]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[2]_i_1__28_n_0 ),
        .Q(\rgf/bank02/gr22 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[3]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[4]_i_1__28_n_0 ),
        .Q(\rgf/bank02/gr22 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[5]_i_1__28_n_0 ),
        .Q(\rgf/bank02/gr22 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[6]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[7]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[8]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn22/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__15_n_0 ),
        .D(\grn[9]_i_1__17_n_0 ),
        .Q(\rgf/bank02/gr22 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[0]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[10]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[11]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[12]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[13]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[14]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[15]_i_2__18_n_0 ),
        .Q(\rgf/bank02/gr23 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[1]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[2]_i_1__27_n_0 ),
        .Q(\rgf/bank02/gr23 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[3]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[4]_i_1__27_n_0 ),
        .Q(\rgf/bank02/gr23 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[5]_i_1__27_n_0 ),
        .Q(\rgf/bank02/gr23 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[6]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[7]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[8]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn23/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__24_n_0 ),
        .D(\grn[9]_i_1__18_n_0 ),
        .Q(\rgf/bank02/gr23 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[0]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[10]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[11]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[12]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[13]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[14]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[15]_i_2__19_n_0 ),
        .Q(\rgf/bank02/gr24 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[1]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[2]_i_1__26_n_0 ),
        .Q(\rgf/bank02/gr24 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[3]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[4]_i_1__26_n_0 ),
        .Q(\rgf/bank02/gr24 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[5]_i_1__26_n_0 ),
        .Q(\rgf/bank02/gr24 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[6]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[7]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[8]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn24/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__14_n_0 ),
        .D(\grn[9]_i_1__19_n_0 ),
        .Q(\rgf/bank02/gr24 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[0]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[10]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[11]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[12]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[13]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[14]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[15]_i_2__20_n_0 ),
        .Q(\rgf/bank02/gr25 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[1]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[2]_i_1__25_n_0 ),
        .Q(\rgf/bank02/gr25 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[3]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[4]_i_1__25_n_0 ),
        .Q(\rgf/bank02/gr25 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[5]_i_1__25_n_0 ),
        .Q(\rgf/bank02/gr25 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[6]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[7]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[8]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn25/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__13_n_0 ),
        .D(\grn[9]_i_1__20_n_0 ),
        .Q(\rgf/bank02/gr25 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[0]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[10]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[11]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[12]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[13]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[14]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[15]_i_2__21_n_0 ),
        .Q(\rgf/bank02/gr26 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[1]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[2]_i_1__24_n_0 ),
        .Q(\rgf/bank02/gr26 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[3]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[4]_i_1__24_n_0 ),
        .Q(\rgf/bank02/gr26 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[5]_i_1__24_n_0 ),
        .Q(\rgf/bank02/gr26 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[6]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[7]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[8]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn26/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__12_n_0 ),
        .D(\grn[9]_i_1__21_n_0 ),
        .Q(\rgf/bank02/gr26 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[0]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[10]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[11]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[12]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[13]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[14]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[15]_i_2__22_n_0 ),
        .Q(\rgf/bank02/gr27 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[1]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[2]_i_1__23_n_0 ),
        .Q(\rgf/bank02/gr27 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[3]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[4]_i_1__23_n_0 ),
        .Q(\rgf/bank02/gr27 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[5]_i_1__23_n_0 ),
        .Q(\rgf/bank02/gr27 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[6]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[7]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[8]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank02/grn27/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__11_n_0 ),
        .D(\grn[9]_i_1__22_n_0 ),
        .Q(\rgf/bank02/gr27 [9]),
        .R(\alu1/div/p_0_in__0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/niss_dsp_b1[3]_INST_0_i_6 
       (.I0(\rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_14_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_15_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[3]_INST_0_i_16_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_17_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_18_n_0 ),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_19_n_0 ),
        .O(\rgf/b1bus_b02 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/niss_dsp_b1[5]_INST_0_i_6 
       (.I0(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_16_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_17_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/niss_dsp_b1[5]_INST_0_i_18_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_20_n_0 ),
        .I5(\rgf/bank02/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_21_n_0 ),
        .O(\rgf/b1bus_b02 [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank02/rgf_c1bus_wb[31]_i_69 
       (.I0(\rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_80_n_0 ),
        .I1(\rgf/bank02/b1buso/i_/bdatw[12]_INST_0_i_32_n_0 ),
        .I2(\rgf/bank02/b1buso/i_/rgf_c1bus_wb[31]_i_81_n_0 ),
        .I3(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_37_n_0 ),
        .I4(\rgf/bank02/b1buso2l/i_/bdatw[12]_INST_0_i_36_n_0 ),
        .I5(\rgf/bank02/b1buso2l/i_/rgf_c1bus_wb[31]_i_82_n_0 ),
        .O(\rgf/b1bus_b02 [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_34 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [0]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [0]),
        .I4(\badr[0]_INST_0_i_44_n_0 ),
        .I5(\badr[0]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[0]_INST_0_i_35 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [0]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [0]),
        .I4(\badr[0]_INST_0_i_46_n_0 ),
        .I5(\badr[0]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_37 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [10]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [10]),
        .I4(\badr[10]_INST_0_i_45_n_0 ),
        .I5(\badr[10]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[10]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [10]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [10]),
        .I4(\badr[10]_INST_0_i_47_n_0 ),
        .I5(\badr[10]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_37 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [11]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [11]),
        .I4(\badr[11]_INST_0_i_45_n_0 ),
        .I5(\badr[11]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[11]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [11]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [11]),
        .I4(\badr[11]_INST_0_i_47_n_0 ),
        .I5(\badr[11]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [12]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [12]),
        .I4(\badr[12]_INST_0_i_50_n_0 ),
        .I5(\badr[12]_INST_0_i_51_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[12]_INST_0_i_39 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [12]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [12]),
        .I4(\badr[12]_INST_0_i_52_n_0 ),
        .I5(\badr[12]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_40 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [13]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [13]),
        .I4(\badr[13]_INST_0_i_49_n_0 ),
        .I5(\badr[13]_INST_0_i_50_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[13]_INST_0_i_41 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [13]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [13]),
        .I4(\badr[13]_INST_0_i_51_n_0 ),
        .I5(\badr[13]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_33 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [14]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [14]),
        .I4(\badr[14]_INST_0_i_43_n_0 ),
        .I5(\badr[14]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[14]_INST_0_i_34 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [14]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [14]),
        .I4(\badr[14]_INST_0_i_45_n_0 ),
        .I5(\badr[14]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_101 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[15]_INST_0_i_132_n_0 ),
        .I4(\badr[0]_INST_0_i_25_n_0 ),
        .O(\bank13/a0buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_102 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\badr[15]_INST_0_i_99_n_0 ),
        .I5(\badr[15]_INST_0_i_100_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_39 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\badr[15]_INST_0_i_103_n_0 ),
        .I5(\badr[15]_INST_0_i_104_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_97 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a0buso/i_/badr[15]_INST_0_i_98 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[0]_INST_0_i_25_n_0 ),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_33 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [1]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [1]),
        .I4(\badr[1]_INST_0_i_43_n_0 ),
        .I5(\badr[1]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[1]_INST_0_i_34 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [1]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [1]),
        .I4(\badr[1]_INST_0_i_45_n_0 ),
        .I5(\badr[1]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_33 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [2]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [2]),
        .I4(\badr[2]_INST_0_i_43_n_0 ),
        .I5(\badr[2]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[2]_INST_0_i_34 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [2]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [2]),
        .I4(\badr[2]_INST_0_i_45_n_0 ),
        .I5(\badr[2]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_33 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [3]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [3]),
        .I4(\badr[3]_INST_0_i_43_n_0 ),
        .I5(\badr[3]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[3]_INST_0_i_34 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [3]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [3]),
        .I4(\badr[3]_INST_0_i_45_n_0 ),
        .I5(\badr[3]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_34 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [4]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [4]),
        .I4(\badr[4]_INST_0_i_50_n_0 ),
        .I5(\badr[4]_INST_0_i_51_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[4]_INST_0_i_35 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [4]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [4]),
        .I4(\badr[4]_INST_0_i_52_n_0 ),
        .I5(\badr[4]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_37 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [5]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [5]),
        .I4(\badr[5]_INST_0_i_45_n_0 ),
        .I5(\badr[5]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[5]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [5]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [5]),
        .I4(\badr[5]_INST_0_i_47_n_0 ),
        .I5(\badr[5]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_37 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [6]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [6]),
        .I4(\badr[6]_INST_0_i_45_n_0 ),
        .I5(\badr[6]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[6]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [6]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [6]),
        .I4(\badr[6]_INST_0_i_47_n_0 ),
        .I5(\badr[6]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_37 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [7]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [7]),
        .I4(\badr[7]_INST_0_i_45_n_0 ),
        .I5(\badr[7]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[7]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [7]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [7]),
        .I4(\badr[7]_INST_0_i_47_n_0 ),
        .I5(\badr[7]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [8]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [8]),
        .I4(\badr[8]_INST_0_i_50_n_0 ),
        .I5(\badr[8]_INST_0_i_51_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[8]_INST_0_i_39 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [8]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [8]),
        .I4(\badr[8]_INST_0_i_52_n_0 ),
        .I5(\badr[8]_INST_0_i_53_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_37 
       (.I0(\bank13/a0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [9]),
        .I2(\bank13/a0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [9]),
        .I4(\badr[9]_INST_0_i_45_n_0 ),
        .I5(\badr[9]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso/i_/badr[9]_INST_0_i_38 
       (.I0(\bank13/a0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [9]),
        .I2(\bank13/a0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [9]),
        .I4(\badr[9]_INST_0_i_47_n_0 ),
        .I5(\badr[9]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\badr[16]_INST_0_i_26_n_0 ),
        .I5(\badr[16]_INST_0_i_27_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\badr[16]_INST_0_i_28_n_0 ),
        .I5(\badr[16]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[16]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\badr[17]_INST_0_i_25_n_0 ),
        .I5(\badr[17]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\badr[17]_INST_0_i_27_n_0 ),
        .I5(\badr[17]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[17]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\badr[18]_INST_0_i_25_n_0 ),
        .I5(\badr[18]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\badr[18]_INST_0_i_27_n_0 ),
        .I5(\badr[18]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[18]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\badr[19]_INST_0_i_25_n_0 ),
        .I5(\badr[19]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\badr[19]_INST_0_i_27_n_0 ),
        .I5(\badr[19]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[19]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\badr[20]_INST_0_i_26_n_0 ),
        .I5(\badr[20]_INST_0_i_27_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\badr[20]_INST_0_i_28_n_0 ),
        .I5(\badr[20]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[20]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\badr[21]_INST_0_i_25_n_0 ),
        .I5(\badr[21]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\badr[21]_INST_0_i_27_n_0 ),
        .I5(\badr[21]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[21]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\badr[22]_INST_0_i_25_n_0 ),
        .I5(\badr[22]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\badr[22]_INST_0_i_27_n_0 ),
        .I5(\badr[22]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[22]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\badr[23]_INST_0_i_25_n_0 ),
        .I5(\badr[23]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\badr[23]_INST_0_i_27_n_0 ),
        .I5(\badr[23]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[23]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\badr[24]_INST_0_i_26_n_0 ),
        .I5(\badr[24]_INST_0_i_27_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\badr[24]_INST_0_i_28_n_0 ),
        .I5(\badr[24]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[24]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\badr[25]_INST_0_i_25_n_0 ),
        .I5(\badr[25]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\badr[25]_INST_0_i_27_n_0 ),
        .I5(\badr[25]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[25]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\badr[26]_INST_0_i_25_n_0 ),
        .I5(\badr[26]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\badr[26]_INST_0_i_27_n_0 ),
        .I5(\badr[26]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[26]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\badr[27]_INST_0_i_25_n_0 ),
        .I5(\badr[27]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\badr[27]_INST_0_i_27_n_0 ),
        .I5(\badr[27]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[27]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\badr[28]_INST_0_i_26_n_0 ),
        .I5(\badr[28]_INST_0_i_27_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\badr[28]_INST_0_i_28_n_0 ),
        .I5(\badr[28]_INST_0_i_29_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[28]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\badr[29]_INST_0_i_25_n_0 ),
        .I5(\badr[29]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\badr[29]_INST_0_i_27_n_0 ),
        .I5(\badr[29]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[29]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_12 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\badr[30]_INST_0_i_25_n_0 ),
        .I5(\badr[30]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_13 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\badr[30]_INST_0_i_27_n_0 ),
        .I5(\badr[30]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[30]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_14 
       (.I0(\bank13/a0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/a0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\badr[31]_INST_0_i_51_n_0 ),
        .I5(\badr[31]_INST_0_i_52_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_15 
       (.I0(\bank13/a0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/a0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\badr[31]_INST_0_i_55_n_0 ),
        .I5(\badr[31]_INST_0_i_56_n_0 ),
        .O(\rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_49 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_80_n_0 ),
        .I4(\badr[31]_INST_0_i_81_n_0 ),
        .O(\bank13/a0buso2h/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_50 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[31]_INST_0_i_80_n_0 ),
        .O(\bank13/a0buso2h/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_53 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_57_n_0 ),
        .I3(\badr[31]_INST_0_i_81_n_0 ),
        .I4(\badr[31]_INST_0_i_80_n_0 ),
        .O(\bank13/a0buso2h/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a0buso2h/i_/badr[31]_INST_0_i_54 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[31]_INST_0_i_58_n_0 ),
        .I2(\badr[31]_INST_0_i_81_n_0 ),
        .I3(\badr[31]_INST_0_i_57_n_0 ),
        .I4(\badr[31]_INST_0_i_80_n_0 ),
        .O(\bank13/a0buso2h/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_36 
       (.I0(\rgf/bank13/gr24 [0]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [0]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_37 
       (.I0(\rgf/bank13/gr22 [0]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [0]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_38 
       (.I0(\rgf/bank13/gr20 [0]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [0]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_39 
       (.I0(\rgf/bank13/gr26 [0]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [0]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_39 
       (.I0(\rgf/bank13/gr24 [10]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [10]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_40 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [10]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_41 
       (.I0(\rgf/bank13/gr20 [10]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [10]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_42 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [10]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_39 
       (.I0(\rgf/bank13/gr24 [11]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [11]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_40 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [11]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_41 
       (.I0(\rgf/bank13/gr20 [11]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [11]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_42 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [11]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_40 
       (.I0(\rgf/bank13/gr24 [12]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [12]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_41 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [12]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_42 
       (.I0(\rgf/bank13/gr20 [12]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [12]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_43 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [12]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_42 
       (.I0(\rgf/bank13/gr24 [13]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [13]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_43 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [13]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_44 
       (.I0(\rgf/bank13/gr20 [13]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [13]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_45 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [13]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_35 
       (.I0(\rgf/bank13/gr24 [14]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [14]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_36 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [14]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_37 
       (.I0(\rgf/bank13/gr20 [14]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [14]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_38 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [14]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_105 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[0]_INST_0_i_25_n_0 ),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso2l/gr4_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_106 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso2l/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_107 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[15]_INST_0_i_131_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso2l/gr2_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_108 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso2l/gr1_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_109 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[0]_INST_0_i_25_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso2l/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_110 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(ctl_sela0_rn),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(\badr[15]_INST_0_i_132_n_0 ),
        .I4(\badr[0]_INST_0_i_25_n_0 ),
        .O(\bank13/a0buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_111 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(ctl_sela0_rn),
        .I3(\badr[15]_INST_0_i_131_n_0 ),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso2l/gr6_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_112 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[0]_INST_0_i_25_n_0 ),
        .I2(\badr[15]_INST_0_i_131_n_0 ),
        .I3(ctl_sela0_rn),
        .I4(\badr[15]_INST_0_i_132_n_0 ),
        .O(\bank13/a0buso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_40 
       (.I0(\rgf/bank13/gr24 [15]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [15]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_41 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [15]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_42 
       (.I0(\rgf/bank13/gr20 [15]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [15]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_43 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [15]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_35 
       (.I0(\rgf/bank13/gr24 [1]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [1]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_36 
       (.I0(\rgf/bank13/gr22 [1]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [1]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_37 
       (.I0(\rgf/bank13/gr20 [1]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [1]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_38 
       (.I0(\rgf/bank13/gr26 [1]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [1]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_35 
       (.I0(\rgf/bank13/gr24 [2]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [2]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_36 
       (.I0(\rgf/bank13/gr22 [2]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [2]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_37 
       (.I0(\rgf/bank13/gr20 [2]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [2]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_38 
       (.I0(\rgf/bank13/gr26 [2]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [2]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_35 
       (.I0(\rgf/bank13/gr24 [3]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [3]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_36 
       (.I0(\rgf/bank13/gr22 [3]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [3]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_37 
       (.I0(\rgf/bank13/gr20 [3]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [3]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_38 
       (.I0(\rgf/bank13/gr26 [3]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [3]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_36 
       (.I0(\rgf/bank13/gr24 [4]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [4]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_37 
       (.I0(\rgf/bank13/gr22 [4]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [4]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_38 
       (.I0(\rgf/bank13/gr20 [4]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [4]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_39 
       (.I0(\rgf/bank13/gr26 [4]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [4]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_39 
       (.I0(\rgf/bank13/gr24 [5]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [5]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_40 
       (.I0(\rgf/bank13/gr22 [5]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [5]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_41 
       (.I0(\rgf/bank13/gr20 [5]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [5]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_42 
       (.I0(\rgf/bank13/gr26 [5]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [5]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_39 
       (.I0(\rgf/bank13/gr24 [6]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [6]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_40 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [6]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_41 
       (.I0(\rgf/bank13/gr20 [6]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [6]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_42 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [6]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_39 
       (.I0(\rgf/bank13/gr24 [7]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [7]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_40 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [7]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_41 
       (.I0(\rgf/bank13/gr20 [7]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [7]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_42 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [7]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_40 
       (.I0(\rgf/bank13/gr24 [8]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [8]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_41 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [8]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_42 
       (.I0(\rgf/bank13/gr20 [8]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [8]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_43 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [8]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_39 
       (.I0(\rgf/bank13/gr24 [9]),
        .I1(\bank13/a0buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr23 [9]),
        .I3(\bank13/a0buso2l/gr3_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_40 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\bank13/a0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [9]),
        .I3(\bank13/a0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_41 
       (.I0(\rgf/bank13/gr20 [9]),
        .I1(\bank13/a0buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [9]),
        .I3(\bank13/a0buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_42 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\bank13/a0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [9]),
        .I3(\bank13/a0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_19 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [0]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [0]),
        .I4(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_20 
       (.I0(\rgf/bank13/gr00 [0]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [0]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_21 
       (.I0(\rgf/bank13/gr06 [0]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [0]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[0]_INST_0_i_42 
       (.I0(\rgf/bank13/gr02 [0]),
        .I1(\rgf/bank13/gr01 [0]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [10]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [10]),
        .I4(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [10]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [10]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[10]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\rgf/bank13/gr01 [10]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [11]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [11]),
        .I4(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [11]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [11]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[11]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\rgf/bank13/gr01 [11]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [12]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [12]),
        .I4(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [12]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [12]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[12]_INST_0_i_44 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\rgf/bank13/gr01 [12]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_26 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [13]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [13]),
        .I4(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_27 
       (.I0(\rgf/bank13/gr00 [13]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [13]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_28 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[13]_INST_0_i_47 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\rgf/bank13/gr01 [13]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_19 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [14]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [14]),
        .I4(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_20 
       (.I0(\rgf/bank13/gr00 [14]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [14]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_21 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[14]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\rgf/bank13/gr01 [14]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_22 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_69_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_23 
       (.I0(\rgf/bank13/gr00 [15]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [15]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_24 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_67 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_68 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[31]_INST_0_i_19_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_69 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\rgf/bank13/gr01 [15]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_69_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_70 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_71 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_67_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .O(\bank13/a1buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_72 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso/gr6_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a1buso/i_/badr[15]_INST_0_i_73 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso/gr5_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_19 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [1]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [1]),
        .I4(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_20 
       (.I0(\rgf/bank13/gr00 [1]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [1]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_21 
       (.I0(\rgf/bank13/gr06 [1]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [1]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[1]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [1]),
        .I1(\rgf/bank13/gr01 [1]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_19 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [2]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [2]),
        .I4(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_20 
       (.I0(\rgf/bank13/gr00 [2]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [2]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_21 
       (.I0(\rgf/bank13/gr06 [2]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [2]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[2]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [2]),
        .I1(\rgf/bank13/gr01 [2]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_19 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [3]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [3]),
        .I4(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_20 
       (.I0(\rgf/bank13/gr00 [3]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [3]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_21 
       (.I0(\rgf/bank13/gr06 [3]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [3]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [3]),
        .I1(\rgf/bank13/gr01 [3]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_19 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [4]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [4]),
        .I4(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_20 
       (.I0(\rgf/bank13/gr00 [4]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [4]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_21 
       (.I0(\rgf/bank13/gr06 [4]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [4]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[4]_INST_0_i_42 
       (.I0(\rgf/bank13/gr02 [4]),
        .I1(\rgf/bank13/gr01 [4]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [5]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [5]),
        .I4(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [5]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [5]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[5]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [5]),
        .I1(\rgf/bank13/gr01 [5]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [6]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [6]),
        .I4(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [6]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [6]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[6]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\rgf/bank13/gr01 [6]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [7]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [7]),
        .I4(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [7]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [7]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[7]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\rgf/bank13/gr01 [7]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [8]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [8]),
        .I4(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [8]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [8]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[8]_INST_0_i_44 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\rgf/bank13/gr01 [8]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_23 
       (.I0(\bank13/a1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [9]),
        .I2(\bank13/a1buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [9]),
        .I4(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_24 
       (.I0(\rgf/bank13/gr00 [9]),
        .I1(\bank13/a1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr07 [9]),
        .I3(\bank13/a1buso/gr7_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\bank13/a1buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\bank13/a1buso/gr5_bus1 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso/i_/badr[9]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\rgf/bank13/gr01 [9]),
        .I2(\grn[15]_i_4__7_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_36 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [14]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [14]),
        .I4(\rgf_c1bus_wb[10]_i_39_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_40_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[10]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[19]_i_43 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [15]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [15]),
        .I4(\rgf_c1bus_wb[19]_i_45_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_46_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[19]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_57 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [2]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [2]),
        .I4(\rgf_c1bus_wb[28]_i_75_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_76_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_59 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [1]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [1]),
        .I4(\rgf_c1bus_wb[28]_i_79_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_80_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_64 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [4]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [4]),
        .I4(\rgf_c1bus_wb[28]_i_85_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_86_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_66 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [3]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [3]),
        .I4(\rgf_c1bus_wb[28]_i_89_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_90_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[28]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso/i_/rgf_c1bus_wb[4]_i_29 
       (.I0(\bank13/a1buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [0]),
        .I2(\bank13/a1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [0]),
        .I4(\rgf_c1bus_wb[4]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_31_n_0 ),
        .O(\rgf/bank13/a1buso/i_/rgf_c1bus_wb[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [0]),
        .I1(\rgf/bank13/gr21 [0]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\badr[16]_INST_0_i_18_n_0 ),
        .I5(\badr[16]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[16]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [1]),
        .I1(\rgf/bank13/gr21 [1]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\badr[17]_INST_0_i_18_n_0 ),
        .I5(\badr[17]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[17]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [2]),
        .I1(\rgf/bank13/gr21 [2]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\badr[18]_INST_0_i_18_n_0 ),
        .I5(\badr[18]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[18]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [3]),
        .I1(\rgf/bank13/gr21 [3]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\badr[19]_INST_0_i_18_n_0 ),
        .I5(\badr[19]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[19]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [4]),
        .I1(\rgf/bank13/gr21 [4]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\badr[20]_INST_0_i_18_n_0 ),
        .I5(\badr[20]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[20]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [5]),
        .I1(\rgf/bank13/gr21 [5]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\badr[21]_INST_0_i_18_n_0 ),
        .I5(\badr[21]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[21]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\rgf/bank13/gr21 [6]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\badr[22]_INST_0_i_18_n_0 ),
        .I5(\badr[22]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[22]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\rgf/bank13/gr21 [7]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\badr[23]_INST_0_i_18_n_0 ),
        .I5(\badr[23]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[23]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\rgf/bank13/gr21 [8]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\badr[24]_INST_0_i_18_n_0 ),
        .I5(\badr[24]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[24]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\rgf/bank13/gr21 [9]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\badr[25]_INST_0_i_18_n_0 ),
        .I5(\badr[25]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[25]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\rgf/bank13/gr21 [10]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\badr[26]_INST_0_i_18_n_0 ),
        .I5(\badr[26]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[26]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\rgf/bank13/gr21 [11]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\badr[27]_INST_0_i_18_n_0 ),
        .I5(\badr[27]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[27]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\rgf/bank13/gr21 [12]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\badr[28]_INST_0_i_18_n_0 ),
        .I5(\badr[28]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[28]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\rgf/bank13/gr21 [13]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\badr[29]_INST_0_i_18_n_0 ),
        .I5(\badr[29]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[29]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_20 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\rgf/bank13/gr21 [14]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_6 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\badr[30]_INST_0_i_18_n_0 ),
        .I5(\badr[30]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_7 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[30]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_28 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_67_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .O(\bank13/a1buso2h/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_29 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2h/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_32 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2h/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_33 
       (.I0(\rgf/bank13/bank_sel00_out ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[31]_INST_0_i_19_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2h/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_34 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\rgf/bank13/gr21 [15]),
        .I2(\rgf/bank13/bank_sel00_out ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_8 
       (.I0(\bank13/a1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/a1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\badr[31]_INST_0_i_30_n_0 ),
        .I5(\badr[31]_INST_0_i_31_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_9 
       (.I0(\bank13/a1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/a1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_34_n_0 ),
        .O(\rgf/bank13/a1buso2h/i_/badr[31]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_22 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_23 
       (.I0(\rgf/bank13/gr20 [0]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [0]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [0]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [0]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43 
       (.I0(\rgf/bank13/gr22 [0]),
        .I1(\rgf/bank13/gr21 [0]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [10]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [10]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [10]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_44 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\rgf/bank13/gr21 [10]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [11]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [11]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [11]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_44 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\rgf/bank13/gr21 [11]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [12]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [12]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [12]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_45 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\rgf/bank13/gr21 [12]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_29 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_30 
       (.I0(\rgf/bank13/gr20 [13]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [13]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_31 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [13]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_48 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\rgf/bank13/gr21 [13]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_22 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_23 
       (.I0(\rgf/bank13/gr20 [14]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [14]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [14]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\rgf/bank13/gr21 [14]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_25 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_76_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_26 
       (.I0(\rgf/bank13/gr20 [15]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [15]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_27 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [15]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_74 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2l/gr3_bus1 ));
  LUT5 #(
    .INIT(32'h00000020)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_75 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[31]_INST_0_i_19_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_76 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\rgf/bank13/gr21 [15]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_77 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2l/gr0_bus1 ));
  LUT5 #(
    .INIT(32'h00800000)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_78 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_67_n_0 ),
        .I4(\badr[31]_INST_0_i_19_n_0 ),
        .O(\bank13/a1buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_79 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[15]_INST_0_i_15_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2l/gr6_bus1 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_80 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\badr[31]_INST_0_i_19_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[31]_INST_0_i_67_n_0 ),
        .O(\bank13/a1buso2l/gr5_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_22 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_23 
       (.I0(\rgf/bank13/gr20 [1]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [1]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [1]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [1]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [1]),
        .I1(\rgf/bank13/gr21 [1]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_22 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_23 
       (.I0(\rgf/bank13/gr20 [2]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [2]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [2]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [2]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [2]),
        .I1(\rgf/bank13/gr21 [2]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_22 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_23 
       (.I0(\rgf/bank13/gr20 [3]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [3]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [3]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [3]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [3]),
        .I1(\rgf/bank13/gr21 [3]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_22 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_23 
       (.I0(\rgf/bank13/gr20 [4]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [4]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_24 
       (.I0(\rgf/bank13/gr26 [4]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [4]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_43 
       (.I0(\rgf/bank13/gr22 [4]),
        .I1(\rgf/bank13/gr21 [4]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [5]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [5]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [5]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [5]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_44 
       (.I0(\rgf/bank13/gr22 [5]),
        .I1(\rgf/bank13/gr21 [5]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [6]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [6]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [6]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_44 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\rgf/bank13/gr21 [6]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [7]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [7]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [7]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_44 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\rgf/bank13/gr21 [7]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [8]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [8]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [8]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_45 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\rgf/bank13/gr21 [8]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_26 
       (.I0(\bank13/a1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/a1buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_27 
       (.I0(\rgf/bank13/gr20 [9]),
        .I1(\bank13/a1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr27 [9]),
        .I3(\bank13/a1buso2l/gr7_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\bank13/a1buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [9]),
        .I3(\bank13/a1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000C0A000)) 
    \rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_44 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\rgf/bank13/gr21 [9]),
        .I2(\badr[15]_INST_0_i_128_n_0 ),
        .I3(\badr[15]_INST_0_i_14_n_0 ),
        .I4(\badr[15]_INST_0_i_15_n_0 ),
        .I5(\badr[31]_INST_0_i_68_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_54 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\rgf_c1bus_wb[28]_i_71_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_72_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_60 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\rgf_c1bus_wb[28]_i_81_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_82_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_67 
       (.I0(\bank13/a1buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/a1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\rgf_c1bus_wb[28]_i_91_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_92_n_0 ),
        .O(\rgf/bank13/a1buso2l/i_/rgf_c1bus_wb[28]_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_25_n_0 ),
        .I1(\bank13/b0buso/gr1_bus1 ),
        .I2(\rgf/bank13/gr01 [0]),
        .I3(\bank13/b0buso/gr2_bus1 ),
        .I4(\rgf/bank13/gr02 [0]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [0]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [0]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_25 
       (.I0(\rgf/bank13/gr04 [0]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr03 [0]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26 
       (.I0(\rgf/bank13/gr06 [0]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [0]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[0]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_14 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [1]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [1]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_15 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_23_n_0 ),
        .I1(\bank13/b0buso/gr1_bus1 ),
        .I2(\rgf/bank13/gr01 [1]),
        .I3(\bank13/b0buso/gr2_bus1 ),
        .I4(\rgf/bank13/gr02 [1]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_22 
       (.I0(\rgf/bank13/gr06 [1]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [1]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [1]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr03 [1]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[1]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_14 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [2]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [2]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_15 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_23_n_0 ),
        .I1(\bank13/b0buso/gr1_bus1 ),
        .I2(\rgf/bank13/gr01 [2]),
        .I3(\bank13/b0buso/gr2_bus1 ),
        .I4(\rgf/bank13/gr02 [2]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_22 
       (.I0(\rgf/bank13/gr06 [2]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [2]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [2]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr03 [2]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[2]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_15 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [3]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [3]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_23_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_16 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_24_n_0 ),
        .I1(\bank13/b0buso/gr1_bus1 ),
        .I2(\rgf/bank13/gr01 [3]),
        .I3(\bank13/b0buso/gr2_bus1 ),
        .I4(\rgf/bank13/gr02 [3]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_23 
       (.I0(\rgf/bank13/gr06 [3]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [3]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_24 
       (.I0(\rgf/bank13/gr04 [3]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr03 [3]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[3]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_14 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [4]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [4]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_15 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_23_n_0 ),
        .I1(\bank13/b0buso/gr1_bus1 ),
        .I2(\rgf/bank13/gr01 [4]),
        .I3(\bank13/b0buso/gr2_bus1 ),
        .I4(\rgf/bank13/gr02 [4]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_22 
       (.I0(\rgf/bank13/gr06 [4]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_23 
       (.I0(\rgf/bank13/gr04 [4]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr03 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[4]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21 
       (.I0(\bank13/b0buso/gr7_bus1 ),
        .I1(\rgf/bank13/gr07 [5]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr00 [5]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_39_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_40_n_0 ),
        .I1(\bank13/b0buso/gr1_bus1 ),
        .I2(\rgf/bank13/gr01 [5]),
        .I3(\bank13/b0buso/gr2_bus1 ),
        .I4(\rgf/bank13/gr02 [5]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_39 
       (.I0(\rgf/bank13/gr06 [5]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr05 [5]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_40 
       (.I0(\rgf/bank13/gr04 [5]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr03 [5]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_41 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [1]),
        .O(\bank13/b0buso/gr1_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bbus_o[5]_INST_0_i_42 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .O(\bank13/b0buso/gr2_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [6]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_16 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [6]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [6]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_9 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/gr00 [6]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [6]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[6]_INST_0_i_16_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [7]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_16 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [7]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [7]),
        .I4(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_9 
       (.I0(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/gr00 [7]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [7]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bbus_o[7]_INST_0_i_16_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_23 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/gr00 [10]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [10]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_37 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [10]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_38 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [10]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [10]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_47 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[10]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_23 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/gr00 [11]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [11]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_37 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [11]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_38 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [11]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [11]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[11]_INST_0_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_27 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_56_n_0 ),
        .I1(\rgf/bank13/gr00 [12]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [12]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_57_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_56 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [12]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_57 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [12]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [12]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_74_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_74 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[12]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_18 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_32_n_0 ),
        .I1(\rgf/bank13/gr00 [13]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [13]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_33_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_32 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [13]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_33 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [13]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [13]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_42 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[13]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_19 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/gr00 [14]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [14]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_34_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_33 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [14]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_34 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [14]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [14]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_43 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[14]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_27 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_54_n_0 ),
        .I1(\rgf/bank13/gr00 [15]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [15]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_57_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_54 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [15]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_55 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .O(\bank13/b0buso/gr0_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_56 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [7]),
        .O(\bank13/b0buso/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_57 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [15]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_84_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_57_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_80 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .O(\bank13/b0buso/gr6_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_81 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [5]),
        .O(\bank13/b0buso/gr5_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_82 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [3]),
        .O(\bank13/b0buso/gr3_bus1 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_83 
       (.I0(\rgf/sreg/sr [1]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [0]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .O(\bank13/b0buso/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_84 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[15]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_19 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank13/gr00 [8]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [8]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_36_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_35 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [8]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_36 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [8]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [8]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_45 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[8]_INST_0_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_21 
       (.I0(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank13/gr00 [9]),
        .I2(\bank13/b0buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [9]),
        .I4(\bank13/b0buso/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_36_n_0 ),
        .O(\rgf/bank13/p_1_in3_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_35 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\bank13/b0buso/gr6_bus1 ),
        .I2(\rgf/bank13/gr05 [9]),
        .I3(\bank13/b0buso/gr5_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_36 
       (.I0(\bank13/b0buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [9]),
        .I2(\bank13/b0buso/gr4_bus1 ),
        .I3(\rgf/bank13/gr04 [9]),
        .I4(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_45_n_0 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_45 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\bank13/b0buso/gr2_bus1 ),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\bank13/b0buso/gr1_bus1 ),
        .O(\rgf/bank13/b0buso/i_/bdatw[9]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\bdatw[16]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\bdatw[16]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[16]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\bdatw[17]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\bdatw[17]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[17]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\bdatw[18]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\bdatw[18]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[18]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\bdatw[19]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\bdatw[19]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[19]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\bdatw[20]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\bdatw[20]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[20]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\bdatw[21]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\bdatw[21]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[21]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\bdatw[22]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\bdatw[22]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[22]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\bdatw[23]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\bdatw[23]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[23]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\bdatw[24]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\bdatw[24]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[24]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\bdatw[25]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\bdatw[25]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[25]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\bdatw[26]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\bdatw[26]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[26]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\bdatw[27]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\bdatw[27]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[27]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\bdatw[28]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\bdatw[28]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[28]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\bdatw[29]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\bdatw[29]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[29]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_11 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\bdatw[30]_INST_0_i_19_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_12 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\bdatw[30]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[30]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_21 
       (.I0(\bank13/b0buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/b0buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\bdatw[31]_INST_0_i_59_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_22 
       (.I0(\bank13/b0buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/b0buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\bdatw[31]_INST_0_i_62_n_0 ),
        .O(\rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_57 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [3]),
        .O(\bank13/b0buso2h/gr3_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_58 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [4]),
        .O(\bank13/b0buso2h/gr4_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_60 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [7]),
        .O(\bank13/b0buso2h/gr7_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b0buso2h/i_/bdatw[31]_INST_0_i_61 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b0bus_sel_0 [0]),
        .O(\bank13/b0buso2h/gr0_bus1 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_20 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_27_n_0 ),
        .I1(\bank13/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [0]),
        .I3(\bank13/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [0]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_21 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_27 
       (.I0(\rgf/bank13/gr24 [0]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr23 [0]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_28 
       (.I0(\rgf/bank13/gr26 [0]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [0]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[0]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_12 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_13 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_21_n_0 ),
        .I1(\bank13/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [1]),
        .I3(\bank13/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [1]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_20 
       (.I0(\rgf/bank13/gr26 [1]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [1]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_21 
       (.I0(\rgf/bank13/gr24 [1]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr23 [1]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[1]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_12 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_13 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_21_n_0 ),
        .I1(\bank13/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [2]),
        .I3(\bank13/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [2]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_20 
       (.I0(\rgf/bank13/gr26 [2]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [2]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_21 
       (.I0(\rgf/bank13/gr24 [2]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr23 [2]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[2]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_13 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_14 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_22_n_0 ),
        .I1(\bank13/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [3]),
        .I3(\bank13/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [3]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_21 
       (.I0(\rgf/bank13/gr26 [3]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [3]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_22 
       (.I0(\rgf/bank13/gr24 [3]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr23 [3]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[3]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_12 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_20_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_13 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_21_n_0 ),
        .I1(\bank13/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [4]),
        .I3(\bank13/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [4]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_20 
       (.I0(\rgf/bank13/gr26 [4]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_21 
       (.I0(\rgf/bank13/gr24 [4]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr23 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[4]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_19 
       (.I0(\bank13/b0buso2l/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_35_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_20 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_36_n_0 ),
        .I1(\bank13/b0buso2l/gr1_bus1 ),
        .I2(\rgf/bank13/gr21 [5]),
        .I3(\bank13/b0buso2l/gr2_bus1 ),
        .I4(\rgf/bank13/gr22 [5]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_35 
       (.I0(\rgf/bank13/gr26 [5]),
        .I1(\rgf/b0bus_sel_0 [6]),
        .I2(\rgf/bank13/gr25 [5]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [5]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_36 
       (.I0(\rgf/bank13/gr24 [5]),
        .I1(\rgf/b0bus_sel_0 [4]),
        .I2(\rgf/bank13/gr23 [5]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b0bus_sel_0 [3]),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [1]),
        .O(\bank13/b0buso2l/gr1_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[5]_INST_0_i_38 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [2]),
        .O(\bank13/b0buso2l/gr2_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_10 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/gr20 [6]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [6]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [6]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_18 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_22 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [6]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[6]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_10 
       (.I0(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/gr20 [7]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [7]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [7]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_18 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_22 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [7]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bbus_o[7]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_24 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank13/gr20 [10]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [10]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_40_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_39 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [10]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_40 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_48 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [10]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[10]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_24 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_39_n_0 ),
        .I1(\rgf/bank13/gr20 [11]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [11]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_40_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_39 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [11]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_40 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_48_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_48 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [11]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[11]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_28 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_58_n_0 ),
        .I1(\rgf/bank13/gr20 [12]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [12]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_59_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_58 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [12]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_58_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_59 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_75_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_75 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [12]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[12]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_19 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank13/gr20 [13]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [13]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_35_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_34 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [13]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_35 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_43_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_43 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [13]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[13]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_20 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank13/gr20 [14]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [14]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_36_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_35 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [14]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_36 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_44_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_44 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [14]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[14]_INST_0_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_28 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_58_n_0 ),
        .I1(\rgf/bank13/gr20 [15]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [15]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_61_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [15]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_58 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [15]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_58_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_59 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [0]),
        .O(\bank13/b0buso2l/gr0_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_60 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [7]),
        .O(\bank13/b0buso2l/gr7_bus1 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_61 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_89_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_61_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_85 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [6]),
        .O(\bank13/b0buso2l/gr6_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_86 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [5]),
        .O(\bank13/b0buso2l/gr5_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_87 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [3]),
        .O(\bank13/b0buso2l/gr3_bus1 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_88 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/sreg/sr [0]),
        .I2(\rgf/sreg/sr [1]),
        .I3(\rgf/b0bus_sel_0 [4]),
        .O(\bank13/b0buso2l/gr4_bus1 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_89 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [15]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[15]_INST_0_i_89_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_20 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/gr20 [8]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [8]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_37 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [8]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_38 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_46 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [8]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[8]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_22 
       (.I0(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/gr20 [9]),
        .I2(\bank13/b0buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [9]),
        .I4(\bank13/b0buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/p_0_in2_in [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_37 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\bank13/b0buso2l/gr6_bus1 ),
        .I2(\rgf/bank13/gr25 [9]),
        .I3(\bank13/b0buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_38 
       (.I0(\bank13/b0buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/b0buso2l/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_46_n_0 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_46 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\bank13/b0buso2l/gr2_bus1 ),
        .I2(\rgf/bank13/gr21 [9]),
        .I3(\bank13/b0buso2l/gr1_bus1 ),
        .O(\rgf/bank13/b0buso2l/i_/bdatw[9]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_15 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank13/gr00 [10]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [10]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [10]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [10]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_26 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [10]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [10]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [10]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [10]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[10]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_14 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_25_n_0 ),
        .I1(\rgf/bank13/gr00 [11]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [11]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_26_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_25 
       (.I0(\rgf/bank13/gr06 [11]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [11]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_26 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [11]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [11]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [11]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [11]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[11]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_20 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_48_n_0 ),
        .I1(\rgf/bank13/gr00 [12]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [12]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_49_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_39 
       (.I0(\bdatw[12]_INST_0_i_60_n_0 ),
        .I1(\bank13/b1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr04 [4]),
        .I3(\bdatw[12]_INST_0_i_61_n_0 ),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [4]),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_40 
       (.I0(\bdatw[12]_INST_0_i_62_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [4]),
        .I3(\bdatw[12]_INST_0_i_63_n_0 ),
        .I4(\bank13/b1buso/gr6_bus1 ),
        .I5(\rgf/bank13/gr06 [4]),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_48 
       (.I0(\rgf/bank13/gr06 [12]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [12]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_49 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [12]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [12]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_70_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_70 
       (.I0(\rgf/bank13/gr02 [12]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [12]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[12]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_13 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_24_n_0 ),
        .I1(\rgf/bank13/gr00 [13]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [13]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_25_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_24 
       (.I0(\rgf/bank13/gr06 [13]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [13]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_25 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [13]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [13]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_38 
       (.I0(\rgf/bank13/gr02 [13]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [13]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[13]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_12 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_21_n_0 ),
        .I1(\rgf/bank13/gr00 [14]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [14]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_21 
       (.I0(\rgf/bank13/gr06 [14]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [14]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_22 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [14]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [14]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37 
       (.I0(\rgf/bank13/gr02 [14]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [14]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[14]_INST_0_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_16 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_31_n_0 ),
        .I1(\rgf/bank13/gr00 [15]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [15]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_34_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_31 
       (.I0(\rgf/bank13/gr06 [15]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [15]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_32 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_63_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_33 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_0[1]),
        .I4(ctl_selb1_0[2]),
        .I5(ctl_selb1_rn[2]),
        .O(\bank13/b1buso/gr7_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_34 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [15]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [15]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_66_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_62 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_65 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso/gr3_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_66 
       (.I0(\rgf/bank13/gr02 [15]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [15]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[15]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_14 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_27_n_0 ),
        .I1(\rgf/bank13/gr00 [8]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [8]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_27 
       (.I0(\rgf/bank13/gr06 [8]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [8]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_28 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [8]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [8]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [8]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [8]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[8]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_15 
       (.I0(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27_n_0 ),
        .I1(\rgf/bank13/gr00 [9]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [9]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27 
       (.I0(\rgf/bank13/gr06 [9]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [9]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_28 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [9]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [9]),
        .I5(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_41_n_0 ),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_41 
       (.I0(\rgf/bank13/gr02 [9]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [9]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/bdatw[9]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_18 
       (.I0(\niss_dsp_b1[0]_INST_0_i_23_n_0 ),
        .I1(\bank13/b1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr04 [0]),
        .I3(\niss_dsp_b1[0]_INST_0_i_24_n_0 ),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [0]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_19 
       (.I0(\niss_dsp_b1[0]_INST_0_i_25_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [0]),
        .I3(\niss_dsp_b1[0]_INST_0_i_26_n_0 ),
        .I4(\bank13/b1buso/gr6_bus1 ),
        .I5(\rgf/bank13/gr06 [0]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_18 
       (.I0(\niss_dsp_b1[1]_INST_0_i_23_n_0 ),
        .I1(\bank13/b1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr04 [1]),
        .I3(\niss_dsp_b1[1]_INST_0_i_24_n_0 ),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [1]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_19 
       (.I0(\niss_dsp_b1[1]_INST_0_i_25_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [1]),
        .I3(\niss_dsp_b1[1]_INST_0_i_26_n_0 ),
        .I4(\bank13/b1buso/gr6_bus1 ),
        .I5(\rgf/bank13/gr06 [1]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[1]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_20 
       (.I0(\niss_dsp_b1[2]_INST_0_i_28_n_0 ),
        .I1(\bank13/b1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr04 [2]),
        .I3(\niss_dsp_b1[2]_INST_0_i_29_n_0 ),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [2]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_21 
       (.I0(\niss_dsp_b1[2]_INST_0_i_30_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [2]),
        .I3(\niss_dsp_b1[2]_INST_0_i_31_n_0 ),
        .I4(\bank13/b1buso/gr6_bus1 ),
        .I5(\rgf/bank13/gr06 [2]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[2]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_10 
       (.I0(\niss_dsp_b1[3]_INST_0_i_22_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [3]),
        .I3(\niss_dsp_b1[3]_INST_0_i_23_n_0 ),
        .I4(\bank13/b1buso/gr6_bus1 ),
        .I5(\rgf/bank13/gr06 [3]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_9 
       (.I0(\niss_dsp_b1[3]_INST_0_i_20_n_0 ),
        .I1(\bank13/b1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr04 [3]),
        .I3(\niss_dsp_b1[3]_INST_0_i_21_n_0 ),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [3]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[3]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_11 
       (.I0(\niss_dsp_b1[5]_INST_0_i_26_n_0 ),
        .I1(\bank13/b1buso/gr4_bus1 ),
        .I2(\rgf/bank13/gr04 [5]),
        .I3(\niss_dsp_b1[5]_INST_0_i_28_n_0 ),
        .I4(\bank13/b1buso/gr2_bus1 ),
        .I5(\rgf/bank13/gr02 [5]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_12 
       (.I0(\niss_dsp_b1[5]_INST_0_i_30_n_0 ),
        .I1(\bank13/b1buso/gr0_bus1 ),
        .I2(\rgf/bank13/gr00 [5]),
        .I3(\niss_dsp_b1[5]_INST_0_i_31_n_0 ),
        .I4(\bank13/b1buso/gr6_bus1 ),
        .I5(\rgf/bank13/gr06 [5]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_27 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_59_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_29 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_61_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[5]_INST_0_i_32 
       (.I0(\grn[15]_i_4__7_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_62_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso/gr6_bus1 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_15 
       (.I0(\rgf/bank13/gr06 [6]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [6]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_16 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [6]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [6]),
        .I5(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [6]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [6]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_9 
       (.I0(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/gr00 [6]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [6]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_16_n_0 ),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[6]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_15 
       (.I0(\rgf/bank13/gr06 [7]),
        .I1(\grn[15]_i_4__7_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr05 [7]),
        .I4(\bank13/b1buso/gr5_bus1 ),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_16 
       (.I0(\bank13/b1buso/gr3_bus1 ),
        .I1(\rgf/bank13/gr03 [7]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/bank13/gr04 [7]),
        .I5(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_21 
       (.I0(\rgf/bank13/gr02 [7]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr01 [7]),
        .I3(\grn[15]_i_4__7_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_9 
       (.I0(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_15_n_0 ),
        .I1(\rgf/bank13/gr00 [7]),
        .I2(\bank13/b1buso/gr0_bus1 ),
        .I3(\rgf/bank13/gr07 [7]),
        .I4(\bank13/b1buso/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_16_n_0 ),
        .O(\rgf/bank13/b1buso/i_/niss_dsp_b1[7]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [0]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [0]),
        .I4(\bdatw[16]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [0]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [0]),
        .I4(\bdatw[16]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[16]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [1]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [1]),
        .I4(\bdatw[17]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [1]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [1]),
        .I4(\bdatw[17]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[17]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [2]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [2]),
        .I4(\bdatw[18]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [2]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [2]),
        .I4(\bdatw[18]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[18]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [3]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [3]),
        .I4(\bdatw[19]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [3]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [3]),
        .I4(\bdatw[19]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[19]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [4]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [4]),
        .I4(\bdatw[20]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [4]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [4]),
        .I4(\bdatw[20]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[20]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [5]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [5]),
        .I4(\bdatw[21]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [5]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [5]),
        .I4(\bdatw[21]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[21]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [6]),
        .I4(\bdatw[22]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [6]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [6]),
        .I4(\bdatw[22]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[22]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [7]),
        .I4(\bdatw[23]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [7]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [7]),
        .I4(\bdatw[23]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[23]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [8]),
        .I4(\bdatw[24]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [8]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [8]),
        .I4(\bdatw[24]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[24]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [9]),
        .I4(\bdatw[25]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [9]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [9]),
        .I4(\bdatw[25]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[25]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [10]),
        .I4(\bdatw[26]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [10]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [10]),
        .I4(\bdatw[26]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[26]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [11]),
        .I4(\bdatw[27]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [11]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [11]),
        .I4(\bdatw[27]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[27]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [12]),
        .I4(\bdatw[28]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [12]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [12]),
        .I4(\bdatw[28]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[28]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [13]),
        .I4(\bdatw[29]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [13]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [13]),
        .I4(\bdatw[29]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[29]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_17 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [14]),
        .I4(\bdatw[30]_INST_0_i_21_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_18 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [14]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [14]),
        .I4(\bdatw[30]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[30]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_38 
       (.I0(\bank13/b1buso2h/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\bank13/b1buso2h/gr4_bus1 ),
        .I3(\rgf/bank13/gr24 [15]),
        .I4(\bdatw[31]_INST_0_i_96_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_39 
       (.I0(\bank13/b1buso2h/gr7_bus1 ),
        .I1(\rgf/bank13/gr27 [15]),
        .I2(\bank13/b1buso2h/gr0_bus1 ),
        .I3(\rgf/bank13/gr20 [15]),
        .I4(\bdatw[31]_INST_0_i_99_n_0 ),
        .O(\rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_94 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [3]),
        .O(\bank13/b1buso2h/gr3_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_95 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .O(\bank13/b1buso2h/gr4_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_97 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [7]),
        .O(\bank13/b1buso2h/gr7_bus1 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf/bank13/b1buso2h/i_/bdatw[31]_INST_0_i_98 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/b1bus_sel_0 [0]),
        .O(\bank13/b1buso2h/gr0_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_16 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_27_n_0 ),
        .I1(\rgf/bank13/gr20 [10]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [10]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_27 
       (.I0(\rgf/bank13/gr26 [10]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [10]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_28 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [10]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [10]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [10]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [10]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[10]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_15 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_27_n_0 ),
        .I1(\rgf/bank13/gr20 [11]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [11]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_28_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_27 
       (.I0(\rgf/bank13/gr26 [11]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [11]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_28 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [11]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [11]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [11]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [11]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[11]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_21 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_50_n_0 ),
        .I1(\rgf/bank13/gr20 [12]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [12]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_51_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_41 
       (.I0(\bdatw[12]_INST_0_i_64_n_0 ),
        .I1(\bank13/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr24 [4]),
        .I3(\bdatw[12]_INST_0_i_65_n_0 ),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [4]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_42 
       (.I0(\bdatw[12]_INST_0_i_66_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [4]),
        .I3(\bdatw[12]_INST_0_i_67_n_0 ),
        .I4(\bank13/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank13/gr26 [4]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_50 
       (.I0(\rgf/bank13/gr26 [12]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [12]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_51 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [12]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [12]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_71_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_71 
       (.I0(\rgf/bank13/gr22 [12]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [12]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[12]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_14 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank13/gr20 [13]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [13]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_27_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_26 
       (.I0(\rgf/bank13/gr26 [13]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [13]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_27 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [13]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [13]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_39_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_39 
       (.I0(\rgf/bank13/gr22 [13]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [13]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[13]_INST_0_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_13 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/gr20 [14]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [14]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_24_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_23 
       (.I0(\rgf/bank13/gr26 [14]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [14]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_24 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [14]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [14]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38 
       (.I0(\rgf/bank13/gr22 [14]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [14]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[14]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_17 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_35_n_0 ),
        .I1(\rgf/bank13/gr20 [15]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [15]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_38_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_35 
       (.I0(\rgf/bank13/gr26 [15]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [15]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\bdatw[15]_INST_0_i_63_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso2l/gr0_bus1 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_37 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(\bdatw[31]_INST_0_i_12_n_0 ),
        .I3(ctl_selb1_0[1]),
        .I4(ctl_selb1_0[2]),
        .I5(ctl_selb1_rn[2]),
        .O(\bank13/b1buso2l/gr7_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_38 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [15]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [15]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_69_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_67 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso2l/gr5_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_68 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\bdatw[15]_INST_0_i_64_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso2l/gr3_bus1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_69 
       (.I0(\rgf/bank13/gr22 [15]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [15]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[15]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_15 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank13/gr20 [8]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [8]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_30_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_29 
       (.I0(\rgf/bank13/gr26 [8]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [8]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_30 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [8]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [8]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [8]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [8]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[8]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_16 
       (.I0(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29_n_0 ),
        .I1(\rgf/bank13/gr20 [9]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [9]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_30_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29 
       (.I0(\rgf/bank13/gr26 [9]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [9]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_30 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [9]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [9]),
        .I5(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_42_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_42 
       (.I0(\rgf/bank13/gr22 [9]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [9]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/bdatw[9]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_20 
       (.I0(\niss_dsp_b1[0]_INST_0_i_27_n_0 ),
        .I1(\bank13/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr24 [0]),
        .I3(\niss_dsp_b1[0]_INST_0_i_28_n_0 ),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [0]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_21 
       (.I0(\niss_dsp_b1[0]_INST_0_i_29_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [0]),
        .I3(\niss_dsp_b1[0]_INST_0_i_30_n_0 ),
        .I4(\bank13/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank13/gr26 [0]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[0]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_20 
       (.I0(\niss_dsp_b1[1]_INST_0_i_27_n_0 ),
        .I1(\bank13/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr24 [1]),
        .I3(\niss_dsp_b1[1]_INST_0_i_28_n_0 ),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [1]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_21 
       (.I0(\niss_dsp_b1[1]_INST_0_i_29_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [1]),
        .I3(\niss_dsp_b1[1]_INST_0_i_30_n_0 ),
        .I4(\bank13/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[1]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_22 
       (.I0(\niss_dsp_b1[2]_INST_0_i_32_n_0 ),
        .I1(\bank13/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr24 [2]),
        .I3(\niss_dsp_b1[2]_INST_0_i_33_n_0 ),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [2]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_23 
       (.I0(\niss_dsp_b1[2]_INST_0_i_34_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [2]),
        .I3(\niss_dsp_b1[2]_INST_0_i_35_n_0 ),
        .I4(\bank13/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank13/gr26 [2]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[2]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_11 
       (.I0(\niss_dsp_b1[3]_INST_0_i_24_n_0 ),
        .I1(\bank13/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr24 [3]),
        .I3(\niss_dsp_b1[3]_INST_0_i_25_n_0 ),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [3]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_12 
       (.I0(\niss_dsp_b1[3]_INST_0_i_26_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [3]),
        .I3(\niss_dsp_b1[3]_INST_0_i_27_n_0 ),
        .I4(\bank13/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[3]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_13 
       (.I0(\niss_dsp_b1[5]_INST_0_i_33_n_0 ),
        .I1(\bank13/b1buso2l/gr4_bus1 ),
        .I2(\rgf/bank13/gr24 [5]),
        .I3(\niss_dsp_b1[5]_INST_0_i_35_n_0 ),
        .I4(\bank13/b1buso2l/gr2_bus1 ),
        .I5(\rgf/bank13/gr22 [5]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEAFFEAFFEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_14 
       (.I0(\niss_dsp_b1[5]_INST_0_i_37_n_0 ),
        .I1(\bank13/b1buso2l/gr0_bus1 ),
        .I2(\rgf/bank13/gr20 [5]),
        .I3(\niss_dsp_b1[5]_INST_0_i_38_n_0 ),
        .I4(\bank13/b1buso2l/gr6_bus1 ),
        .I5(\rgf/bank13/gr26 [5]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_34 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_59_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso2l/gr4_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_36 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_61_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso2l/gr2_bus1 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[5]_INST_0_i_39 
       (.I0(\badr[15]_INST_0_i_128_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_62_n_0 ),
        .I2(ctl_selb1_rn[0]),
        .I3(\bdatw[31]_INST_0_i_12_n_0 ),
        .I4(ctl_selb1_0[1]),
        .I5(ctl_selb1_0[2]),
        .O(\bank13/b1buso2l/gr6_bus1 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_10 
       (.I0(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/gr20 [6]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [6]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [6]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [6]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_18 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [6]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [6]),
        .I5(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_22 
       (.I0(\rgf/bank13/gr22 [6]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [6]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[6]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_10 
       (.I0(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_17_n_0 ),
        .I1(\rgf/bank13/gr20 [7]),
        .I2(\bank13/b1buso2l/gr0_bus1 ),
        .I3(\rgf/bank13/gr27 [7]),
        .I4(\bank13/b1buso2l/gr7_bus1 ),
        .I5(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_18_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFF808080)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_17 
       (.I0(\rgf/bank13/gr26 [7]),
        .I1(\badr[15]_INST_0_i_128_n_0 ),
        .I2(\rgf/b1bus_sel_0 [6]),
        .I3(\rgf/bank13/gr25 [7]),
        .I4(\bank13/b1buso2l/gr5_bus1 ),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8888888)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_18 
       (.I0(\bank13/b1buso2l/gr3_bus1 ),
        .I1(\rgf/bank13/gr23 [7]),
        .I2(\rgf/b1bus_sel_0 [4]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/bank13/gr24 [7]),
        .I5(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_22_n_0 ),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_22 
       (.I0(\rgf/bank13/gr22 [7]),
        .I1(\rgf/b1bus_sel_0 [2]),
        .I2(\rgf/bank13/gr21 [7]),
        .I3(\badr[15]_INST_0_i_128_n_0 ),
        .I4(\rgf/b1bus_sel_0 [1]),
        .O(\rgf/bank13/b1buso2l/i_/niss_dsp_b1[7]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[0]_INST_0_i_11 
       (.I0(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[0]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_37_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_38_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[0]_INST_0_i_39_n_0 ),
        .O(\rgf/a0bus_b13 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[0]_INST_0_i_5 
       (.I0(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[0]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_23_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[0]_INST_0_i_24_n_0 ),
        .O(\rgf/a1bus_b13 [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[10]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[10]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[10]_INST_0_i_42_n_0 ),
        .O(\rgf/a0bus_b13 [10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[10]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[10]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[10]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[11]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[11]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[11]_INST_0_i_42_n_0 ),
        .O(\rgf/a0bus_b13 [11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[11]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[11]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[11]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[12]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[12]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_42_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[12]_INST_0_i_43_n_0 ),
        .O(\rgf/a0bus_b13 [12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[12]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[12]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[12]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[13]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_40_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[13]_INST_0_i_41_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_42_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_43_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_44_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[13]_INST_0_i_45_n_0 ),
        .O(\rgf/a0bus_b13 [13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[13]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_26_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_27_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[13]_INST_0_i_28_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_29_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_30_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[13]_INST_0_i_31_n_0 ),
        .O(\rgf/a1bus_b13 [13]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[14]_INST_0_i_11 
       (.I0(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[14]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_37_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[14]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_b13 [14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[14]_INST_0_i_5 
       (.I0(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[14]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_23_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[14]_INST_0_i_24_n_0 ),
        .O(\rgf/a1bus_b13 [14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[15]_INST_0_i_12 
       (.I0(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[15]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_42_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[15]_INST_0_i_43_n_0 ),
        .O(\rgf/a0bus_b13 [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[15]_INST_0_i_6 
       (.I0(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_22_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_23_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[15]_INST_0_i_24_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_25_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_26_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[15]_INST_0_i_27_n_0 ),
        .O(\rgf/a1bus_b13 [15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[1]_INST_0_i_11 
       (.I0(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[1]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_37_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[1]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_b13 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[1]_INST_0_i_5 
       (.I0(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[1]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_23_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[1]_INST_0_i_24_n_0 ),
        .O(\rgf/a1bus_b13 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[2]_INST_0_i_11 
       (.I0(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[2]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_37_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[2]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_b13 [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[2]_INST_0_i_5 
       (.I0(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[2]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_23_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[2]_INST_0_i_24_n_0 ),
        .O(\rgf/a1bus_b13 [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[3]_INST_0_i_11 
       (.I0(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_33_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[3]_INST_0_i_34_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_35_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_36_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_37_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[3]_INST_0_i_38_n_0 ),
        .O(\rgf/a0bus_b13 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[3]_INST_0_i_5 
       (.I0(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[3]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_23_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[3]_INST_0_i_24_n_0 ),
        .O(\rgf/a1bus_b13 [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[4]_INST_0_i_11 
       (.I0(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_34_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[4]_INST_0_i_35_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_36_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_37_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_38_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[4]_INST_0_i_39_n_0 ),
        .O(\rgf/a0bus_b13 [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[4]_INST_0_i_5 
       (.I0(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_19_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_20_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[4]_INST_0_i_21_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_22_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_23_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[4]_INST_0_i_24_n_0 ),
        .O(\rgf/a1bus_b13 [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[5]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[5]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[5]_INST_0_i_42_n_0 ),
        .O(\rgf/a0bus_b13 [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[5]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[5]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[5]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[6]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[6]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[6]_INST_0_i_42_n_0 ),
        .O(\rgf/a0bus_b13 [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[6]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[6]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[6]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[7]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[7]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[7]_INST_0_i_42_n_0 ),
        .O(\rgf/a0bus_b13 [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[7]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[7]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[7]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [7]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[8]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_38_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[8]_INST_0_i_39_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_40_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_41_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_42_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[8]_INST_0_i_43_n_0 ),
        .O(\rgf/a0bus_b13 [8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[8]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[8]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[8]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [8]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[9]_INST_0_i_13 
       (.I0(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_37_n_0 ),
        .I1(\rgf/bank13/a0buso/i_/badr[9]_INST_0_i_38_n_0 ),
        .I2(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_39_n_0 ),
        .I3(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_40_n_0 ),
        .I4(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_41_n_0 ),
        .I5(\rgf/bank13/a0buso2l/i_/badr[9]_INST_0_i_42_n_0 ),
        .O(\rgf/a0bus_b13 [9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf/bank13/badr[9]_INST_0_i_7 
       (.I0(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_23_n_0 ),
        .I1(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_24_n_0 ),
        .I2(\rgf/bank13/a1buso/i_/badr[9]_INST_0_i_25_n_0 ),
        .I3(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_26_n_0 ),
        .I4(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_27_n_0 ),
        .I5(\rgf/bank13/a1buso2l/i_/badr[9]_INST_0_i_28_n_0 ),
        .O(\rgf/a1bus_b13 [9]));
  FDRE \rgf/bank13/grn00/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[0]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[10]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[11]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[12]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[13]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[14]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[15]_i_2__11_n_0 ),
        .Q(\rgf/bank13/gr00 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[1]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[2]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[3]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[4]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[5]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[6]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[7]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[8]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn00/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__27_n_0 ),
        .D(\grn[9]_i_1__11_n_0 ),
        .Q(\rgf/bank13/gr00 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[0]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[10]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[11]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[12]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[13]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[14]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[15]_i_2__10_n_0 ),
        .Q(\rgf/bank13/gr01 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[1]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[2]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[3]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[4]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[5]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[6]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[7]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[8]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn01/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__19_n_0 ),
        .D(\grn[9]_i_1__10_n_0 ),
        .Q(\rgf/bank13/gr01 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[0]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[10]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[11]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[12]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[13]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[14]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[15]_i_2__12_n_0 ),
        .Q(\rgf/bank13/gr02 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[1]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[2]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[3]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[4]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[5]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[6]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[7]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[8]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn02/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__18_n_0 ),
        .D(\grn[9]_i_1__12_n_0 ),
        .Q(\rgf/bank13/gr02 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[0]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[10]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[11]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[12]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[13]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[14]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[15]_i_2__9_n_0 ),
        .Q(\rgf/bank13/gr03 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[1]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[2]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[3]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[4]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[5]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[6]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[7]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[8]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn03/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__23_n_0 ),
        .D(\grn[9]_i_1__9_n_0 ),
        .Q(\rgf/bank13/gr03 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[0]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[10]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[11]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[12]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[13]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[14]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[15]_i_2__13_n_0 ),
        .Q(\rgf/bank13/gr04 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[1]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[2]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[3]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[4]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[5]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[6]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[7]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[8]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn04/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__21_n_0 ),
        .D(\grn[9]_i_1__13_n_0 ),
        .Q(\rgf/bank13/gr04 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[0]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[10]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[11]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[12]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[13]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[14]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[15]_i_2__8_n_0 ),
        .Q(\rgf/bank13/gr05 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[1]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[2]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[3]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[4]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[5]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[6]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[7]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[8]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn05/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__22_n_0 ),
        .D(\grn[9]_i_1__8_n_0 ),
        .Q(\rgf/bank13/gr05 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[0]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[10]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[11]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[12]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[13]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[14]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[15]_i_2__14_n_0 ),
        .Q(\rgf/bank13/gr06 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[1]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[2]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[3]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[4]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[5]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[6]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[7]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[8]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn06/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__20_n_0 ),
        .D(\grn[9]_i_1__14_n_0 ),
        .Q(\rgf/bank13/gr06 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[0]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[10]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[11]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[12]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[13]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[14]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[15]_i_2__7_n_0 ),
        .Q(\rgf/bank13/gr07 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[1]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[2]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[3]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[4]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[5]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[6]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[7]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[8]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn07/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__17_n_0 ),
        .D(\grn[9]_i_1__7_n_0 ),
        .Q(\rgf/bank13/gr07 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[0]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[10]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[11]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[12]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[13]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[14]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[15]_i_2__23_n_0 ),
        .Q(\rgf/bank13/gr20 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[1]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[2]_i_1__22_n_0 ),
        .Q(\rgf/bank13/gr20 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[3]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[4]_i_1__22_n_0 ),
        .Q(\rgf/bank13/gr20 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[5]_i_1__22_n_0 ),
        .Q(\rgf/bank13/gr20 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[6]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[7]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[8]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn20/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__29_n_0 ),
        .D(\grn[9]_i_1__23_n_0 ),
        .Q(\rgf/bank13/gr20 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[0]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[10]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[11]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[12]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[13]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[14]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[15]_i_2__24_n_0 ),
        .Q(\rgf/bank13/gr21 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[1]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[2]_i_1__21_n_0 ),
        .Q(\rgf/bank13/gr21 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[3]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[4]_i_1__21_n_0 ),
        .Q(\rgf/bank13/gr21 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[5]_i_1__21_n_0 ),
        .Q(\rgf/bank13/gr21 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[6]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[7]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[8]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn21/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__10_n_0 ),
        .D(\grn[9]_i_1__24_n_0 ),
        .Q(\rgf/bank13/gr21 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[0]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[10]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[11]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[12]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[13]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[14]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[15]_i_2__25_n_0 ),
        .Q(\rgf/bank13/gr22 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[1]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[2]_i_1__20_n_0 ),
        .Q(\rgf/bank13/gr22 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[3]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[4]_i_1__20_n_0 ),
        .Q(\rgf/bank13/gr22 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[5]_i_1__20_n_0 ),
        .Q(\rgf/bank13/gr22 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[6]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[7]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[8]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn22/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__9_n_0 ),
        .D(\grn[9]_i_1__25_n_0 ),
        .Q(\rgf/bank13/gr22 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[0]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[10]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[11]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[12]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[13]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[14]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[15]_i_2__26_n_0 ),
        .Q(\rgf/bank13/gr23 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[1]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[2]_i_1__19_n_0 ),
        .Q(\rgf/bank13/gr23 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[3]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[4]_i_1__19_n_0 ),
        .Q(\rgf/bank13/gr23 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[5]_i_1__19_n_0 ),
        .Q(\rgf/bank13/gr23 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[6]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[7]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[8]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn23/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__25_n_0 ),
        .D(\grn[9]_i_1__26_n_0 ),
        .Q(\rgf/bank13/gr23 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[0]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[10]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[11]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[12]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[13]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[14]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[15]_i_2__27_n_0 ),
        .Q(\rgf/bank13/gr24 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[1]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[2]_i_1__18_n_0 ),
        .Q(\rgf/bank13/gr24 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[3]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[4]_i_1__18_n_0 ),
        .Q(\rgf/bank13/gr24 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[5]_i_1__18_n_0 ),
        .Q(\rgf/bank13/gr24 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[6]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[7]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[8]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn24/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__8_n_0 ),
        .D(\grn[9]_i_1__27_n_0 ),
        .Q(\rgf/bank13/gr24 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[0]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[10]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[11]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[12]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[13]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[14]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[15]_i_2__28_n_0 ),
        .Q(\rgf/bank13/gr25 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[1]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[2]_i_1__17_n_0 ),
        .Q(\rgf/bank13/gr25 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[3]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[4]_i_1__17_n_0 ),
        .Q(\rgf/bank13/gr25 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[5]_i_1__17_n_0 ),
        .Q(\rgf/bank13/gr25 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[6]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[7]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[8]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn25/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__7_n_0 ),
        .D(\grn[9]_i_1__28_n_0 ),
        .Q(\rgf/bank13/gr25 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[0]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[10]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[11]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[12]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[13]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[14]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[15]_i_2__29_n_0 ),
        .Q(\rgf/bank13/gr26 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[1]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[2]_i_1__16_n_0 ),
        .Q(\rgf/bank13/gr26 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[3]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[4]_i_1__16_n_0 ),
        .Q(\rgf/bank13/gr26 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[5]_i_1__16_n_0 ),
        .Q(\rgf/bank13/gr26 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[6]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[7]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[8]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn26/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__6_n_0 ),
        .D(\grn[9]_i_1__29_n_0 ),
        .Q(\rgf/bank13/gr26 [9]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[0] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[0]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [0]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[10] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[10]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [10]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[11] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[11]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [11]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[12] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[12]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [12]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[13] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[13]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [13]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[14] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[14]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [14]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[15] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[15]_i_2__30_n_0 ),
        .Q(\rgf/bank13/gr27 [15]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[1] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[1]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [1]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[2] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[2]_i_1__15_n_0 ),
        .Q(\rgf/bank13/gr27 [2]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[3] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[3]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [3]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[4] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[4]_i_1__15_n_0 ),
        .Q(\rgf/bank13/gr27 [4]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[5] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[5]_i_1__15_n_0 ),
        .Q(\rgf/bank13/gr27 [5]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[6] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[6]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [6]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[7] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[7]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [7]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[8] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[8]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [8]),
        .R(\alu1/div/p_0_in__0 ));
  FDRE \rgf/bank13/grn27/grn_reg[9] 
       (.C(clk),
        .CE(\grn[15]_i_1__5_n_0 ),
        .D(\grn[9]_i_1__30_n_0 ),
        .Q(\rgf/bank13/gr27 [9]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [0]),
        .Q(\rgf/ivec/iv [0]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [10]),
        .Q(\rgf/ivec/iv [10]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [11]),
        .Q(\rgf/ivec/iv [11]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [12]),
        .Q(\rgf/ivec/iv [12]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [13]),
        .Q(\rgf/ivec/iv [13]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [14]),
        .Q(\rgf/ivec/iv [14]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [15]),
        .Q(\rgf/ivec/iv [15]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [1]),
        .Q(\rgf/ivec/iv [1]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [2]),
        .Q(\rgf/ivec/iv [2]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [3]),
        .Q(\rgf/ivec/iv [3]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [4]),
        .Q(\rgf/ivec/iv [4]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [5]),
        .Q(\rgf/ivec/iv [5]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [6]),
        .Q(\rgf/ivec/iv [6]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [7]),
        .Q(\rgf/ivec/iv [7]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [8]),
        .Q(\rgf/ivec/iv [8]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/ivec/iv_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/ivec/p_1_in [9]),
        .Q(\rgf/ivec/iv [9]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [0]),
        .Q(\rgf/pcnt/pc [0]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [10]),
        .Q(\rgf/pcnt/pc [10]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [11]),
        .Q(\rgf/pcnt/pc [11]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [12]),
        .Q(\rgf/pcnt/pc [12]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [13]),
        .Q(\rgf/pcnt/pc [13]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [14]),
        .Q(\rgf/pcnt/pc [14]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [15]),
        .Q(\rgf/pcnt/pc [15]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [1]),
        .Q(\rgf/pcnt/pc [1]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [2]),
        .Q(\rgf/pcnt/pc [2]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [3]),
        .Q(\rgf/pcnt/pc [3]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [4]),
        .Q(\rgf/pcnt/pc [4]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [5]),
        .Q(\rgf/pcnt/pc [5]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [6]),
        .Q(\rgf/pcnt/pc [6]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [7]),
        .Q(\rgf/pcnt/pc [7]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [8]),
        .Q(\rgf/pcnt/pc [8]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/pcnt/pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/pcnt/p_1_in [9]),
        .Q(\rgf/pcnt/pc [9]),
        .R(\alu1/div/p_0_in__0 ));
  LUT3 #(
    .INIT(8'h54)) 
    \rgf/rctl/grn[15]_i_4 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [1]),
        .O(\rgf/bank_sel [2]));
  LUT3 #(
    .INIT(8'h45)) 
    \rgf/rctl/grn[15]_i_5 
       (.I0(\rgf/sreg/sr [0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/sreg/sr [1]),
        .O(\rgf/bank_sel [0]));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[0]),
        .Q(\rgf/rctl/rgf_c0bus_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[10] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[10]),
        .Q(\rgf/rctl/rgf_c0bus_wb [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[11] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[11]),
        .Q(\rgf/rctl/rgf_c0bus_wb [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[12] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[12]),
        .Q(\rgf/rctl/rgf_c0bus_wb [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[13] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[13]),
        .Q(\rgf/rctl/rgf_c0bus_wb [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[14] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[14]),
        .Q(\rgf/rctl/rgf_c0bus_wb [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[15] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[15]),
        .Q(\rgf/rctl/rgf_c0bus_wb [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[16] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[16]),
        .Q(\rgf/rctl/rgf_c0bus_wb [16]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[17] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[17]),
        .Q(\rgf/rctl/rgf_c0bus_wb [17]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[18] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[18]),
        .Q(\rgf/rctl/rgf_c0bus_wb [18]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[19] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[19]),
        .Q(\rgf/rctl/rgf_c0bus_wb [19]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[1]),
        .Q(\rgf/rctl/rgf_c0bus_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[20] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[20]),
        .Q(\rgf/rctl/rgf_c0bus_wb [20]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[21] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[21]),
        .Q(\rgf/rctl/rgf_c0bus_wb [21]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[22] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[22]),
        .Q(\rgf/rctl/rgf_c0bus_wb [22]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[23] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[23]),
        .Q(\rgf/rctl/rgf_c0bus_wb [23]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[24] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[24]),
        .Q(\rgf/rctl/rgf_c0bus_wb [24]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[25] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[25]),
        .Q(\rgf/rctl/rgf_c0bus_wb [25]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[26] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[26]),
        .Q(\rgf/rctl/rgf_c0bus_wb [26]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[27] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[27]),
        .Q(\rgf/rctl/rgf_c0bus_wb [27]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[28] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[28]),
        .Q(\rgf/rctl/rgf_c0bus_wb [28]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[29] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[29]),
        .Q(\rgf/rctl/rgf_c0bus_wb [29]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[2]),
        .Q(\rgf/rctl/rgf_c0bus_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[30] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[30]),
        .Q(\rgf/rctl/rgf_c0bus_wb [30]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[31] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[31]),
        .Q(\rgf/rctl/rgf_c0bus_wb [31]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[3] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[3]),
        .Q(\rgf/rctl/rgf_c0bus_wb [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[4] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[4]),
        .Q(\rgf/rctl/rgf_c0bus_wb [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[5] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[5]),
        .Q(\rgf/rctl/rgf_c0bus_wb [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[6] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[6]),
        .Q(\rgf/rctl/rgf_c0bus_wb [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[7] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[7]),
        .Q(\rgf/rctl/rgf_c0bus_wb [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[8] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[8]),
        .Q(\rgf/rctl/rgf_c0bus_wb [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c0bus_wb_reg[9] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(c0bus[9]),
        .Q(\rgf/rctl/rgf_c0bus_wb [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[0]),
        .Q(\rgf/rctl/rgf_c1bus_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[10] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[10]),
        .Q(\rgf/rctl/rgf_c1bus_wb [10]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[11] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[11]),
        .Q(\rgf/rctl/rgf_c1bus_wb [11]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[12] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[12]),
        .Q(\rgf/rctl/rgf_c1bus_wb [12]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[13] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[13]),
        .Q(\rgf/rctl/rgf_c1bus_wb [13]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[14] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[14]),
        .Q(\rgf/rctl/rgf_c1bus_wb [14]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[15] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[15]),
        .Q(\rgf/rctl/rgf_c1bus_wb [15]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[16] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[16]),
        .Q(\rgf/rctl/rgf_c1bus_wb [16]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[17] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[17]),
        .Q(\rgf/rctl/rgf_c1bus_wb [17]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[18] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[18]),
        .Q(\rgf/rctl/rgf_c1bus_wb [18]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[19] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[19]),
        .Q(\rgf/rctl/rgf_c1bus_wb [19]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[1]),
        .Q(\rgf/rctl/rgf_c1bus_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[20] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[20]),
        .Q(\rgf/rctl/rgf_c1bus_wb [20]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[21] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[21]),
        .Q(\rgf/rctl/rgf_c1bus_wb [21]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[22] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[22]),
        .Q(\rgf/rctl/rgf_c1bus_wb [22]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[23] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[23]),
        .Q(\rgf/rctl/rgf_c1bus_wb [23]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[24] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[24]),
        .Q(\rgf/rctl/rgf_c1bus_wb [24]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[25] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[25]),
        .Q(\rgf/rctl/rgf_c1bus_wb [25]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[26] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[26]),
        .Q(\rgf/rctl/rgf_c1bus_wb [26]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[27] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[27]),
        .Q(\rgf/rctl/rgf_c1bus_wb [27]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[28] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[28]),
        .Q(\rgf/rctl/rgf_c1bus_wb [28]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[29] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[29]),
        .Q(\rgf/rctl/rgf_c1bus_wb [29]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[2]),
        .Q(\rgf/rctl/rgf_c1bus_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[30] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[30]),
        .Q(\rgf/rctl/rgf_c1bus_wb [30]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[31] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[31]),
        .Q(\rgf/rctl/rgf_c1bus_wb [31]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[3] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[3]),
        .Q(\rgf/rctl/rgf_c1bus_wb [3]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[4] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[4]),
        .Q(\rgf/rctl/rgf_c1bus_wb [4]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[5] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[5]),
        .Q(\rgf/rctl/rgf_c1bus_wb [5]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[6] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[6]),
        .Q(\rgf/rctl/rgf_c1bus_wb [6]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[7] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[7]),
        .Q(\rgf/rctl/rgf_c1bus_wb [7]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[8] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[8]),
        .Q(\rgf/rctl/rgf_c1bus_wb [8]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_c1bus_wb_reg[9] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(c1bus[9]),
        .Q(\rgf/rctl/rgf_c1bus_wb [9]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_rn_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(ctl_selc0_rn),
        .Q(\rgf/rctl/rgf_selc0_rn_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_rn_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(\rgf_selc0_rn_wb[1]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc0_rn_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_rn_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(\rgf_selc0_rn_wb[2]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc0_rn_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_stat_reg 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(\rgf/rctl/p_2_in ),
        .Q(\rgf/rctl/rgf_selc0_stat ),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(ctl_selc0[0]),
        .Q(\rgf/rctl/rgf_selc0_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc0_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc0_stat_i_2_n_0),
        .D(ctl_selc0[1]),
        .Q(\rgf/rctl/rgf_selc0_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_rn_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(ctl_selc1_rn),
        .Q(\rgf/rctl/rgf_selc1_rn_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_rn_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(\rgf_selc1_rn_wb[1]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc1_rn_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_rn_wb_reg[2] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(\rgf_selc1_rn_wb[2]_i_1_n_0 ),
        .Q(\rgf/rctl/rgf_selc1_rn_wb [2]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_stat_reg 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(rgf_selc1_stat_i_2_n_0),
        .Q(\rgf/rctl/rgf_selc1_stat ),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_wb_reg[0] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(ctl_selc1[0]),
        .Q(\rgf/rctl/rgf_selc1_wb [0]),
        .R(rgf_selc0_stat_i_1_n_0));
  FDRE \rgf/rctl/rgf_selc1_wb_reg[1] 
       (.C(clk),
        .CE(rgf_selc1_stat_i_1_n_0),
        .D(ctl_selc1[1]),
        .Q(\rgf/rctl/rgf_selc1_wb [1]),
        .R(rgf_selc0_stat_i_1_n_0));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[0]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [0]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[10]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [10]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[11]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [11]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[12]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [12]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[13]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [13]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[14]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [14]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[15]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [15]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[16]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [16]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[17]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [17]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[18]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [18]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[19]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [19]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[1]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [1]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[20]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [20]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[21]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [21]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[22]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [22]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[23]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [23]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[24]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [24]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[25]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [25]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[26]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [26]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[27]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [27]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[28]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [28]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[29]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [29]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[2]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [2]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[30]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [30]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[31]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [31]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[3]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [3]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[4]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [4]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[5]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [5]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[6]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [6]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[7]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [7]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[8]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [8]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sptr/sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp[9]_i_1_n_0 ),
        .Q(\rgf/sptr/sp [9]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [0]),
        .Q(\rgf/sreg/sr [0]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [10]),
        .Q(\rgf/sreg/sr [10]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [11]),
        .Q(\rgf/sreg/sr [11]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [12]),
        .Q(\rgf/sreg/sr [12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [13]),
        .Q(\rgf/sreg/sr [13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [14]),
        .Q(\rgf/sreg/sr [14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [15]),
        .Q(\rgf/sreg/sr [15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [1]),
        .Q(\rgf/sreg/sr [1]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [2]),
        .Q(\rgf/sreg/sr [2]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [3]),
        .Q(\rgf/sreg/sr [3]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [4]),
        .Q(\rgf/sreg/sr [4]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [5]),
        .Q(\rgf/sreg/sr [5]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [6]),
        .Q(\rgf/sreg/sr [6]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [7]),
        .Q(\rgf/sreg/sr [7]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [8]),
        .Q(\rgf/sreg/sr [8]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/sreg/sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/sreg/p_0_in__0 [9]),
        .Q(\rgf/sreg/sr [9]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [0]),
        .Q(\rgf/treg/tr [0]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [10]),
        .Q(\rgf/treg/tr [10]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [11]),
        .Q(\rgf/treg/tr [11]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [12]),
        .Q(\rgf/treg/tr [12]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [13]),
        .Q(\rgf/treg/tr [13]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [14]),
        .Q(\rgf/treg/tr [14]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [15]),
        .Q(\rgf/treg/tr [15]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [16]),
        .Q(\rgf/treg/tr [16]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [17]),
        .Q(\rgf/treg/tr [17]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [18]),
        .Q(\rgf/treg/tr [18]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [19]),
        .Q(\rgf/treg/tr [19]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [1]),
        .Q(\rgf/treg/tr [1]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [20]),
        .Q(\rgf/treg/tr [20]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [21]),
        .Q(\rgf/treg/tr [21]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [22]),
        .Q(\rgf/treg/tr [22]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [23]),
        .Q(\rgf/treg/tr [23]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [24]),
        .Q(\rgf/treg/tr [24]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [25]),
        .Q(\rgf/treg/tr [25]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [26]),
        .Q(\rgf/treg/tr [26]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [27]),
        .Q(\rgf/treg/tr [27]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [28]),
        .Q(\rgf/treg/tr [28]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [29]),
        .Q(\rgf/treg/tr [29]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [2]),
        .Q(\rgf/treg/tr [2]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [30]),
        .Q(\rgf/treg/tr [30]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [31]),
        .Q(\rgf/treg/tr [31]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [3]),
        .Q(\rgf/treg/tr [3]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [4]),
        .Q(\rgf/treg/tr [4]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [5]),
        .Q(\rgf/treg/tr [5]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [6]),
        .Q(\rgf/treg/tr [6]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [7]),
        .Q(\rgf/treg/tr [7]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [8]),
        .Q(\rgf/treg/tr [8]),
        .R(\alu1/div/p_0_in__0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \rgf/treg/tr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\rgf/treg/p_1_in [9]),
        .Q(\rgf/treg/tr [9]),
        .R(\alu1/div/p_0_in__0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[0]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[0]),
        .I2(\rgf_c0bus_wb[0]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_5_n_0 ),
        .O(c0bus[0]));
  LUT6 #(
    .INIT(64'hBBBBBBBBFBBBBBBB)) 
    \rgf_c0bus_wb[0]_i_10 
       (.I0(\rgf_c0bus_wb[0]_i_20_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[0]_i_21_n_0 ),
        .I3(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_18_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[0]_i_11 
       (.I0(a0bus_0[24]),
        .I1(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I2(a0bus_0[0]),
        .O(\rgf_c0bus_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c0bus_wb[0]_i_12 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(a0bus_0[8]),
        .I3(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I4(a0bus_0[0]),
        .O(\rgf_c0bus_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC0AEC0EE00EA00AA)) 
    \rgf_c0bus_wb[0]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I2(a0bus_0[0]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hD1)) 
    \rgf_c0bus_wb[0]_i_14 
       (.I0(\rgf_c0bus_wb[17]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[0]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h080D)) 
    \rgf_c0bus_wb[0]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[17]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000A033)) 
    \rgf_c0bus_wb[0]_i_17 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\rgf_c0bus_wb[17]_i_10_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[0]_i_18 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c0bus_wb[0]_i_19 
       (.I0(\rgf_c0bus_wb[25]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_22_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_28_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[0]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [0]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[0]),
        .I4(\rgf_c0bus_wb[0]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000B8FFB8)) 
    \rgf_c0bus_wb[0]_i_20 
       (.I0(\rgf_c0bus_wb[16]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_23_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hF7)) 
    \rgf_c0bus_wb[0]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[0]_i_22 
       (.I0(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[0]_i_23 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c0bus_wb[0]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[0]_i_9_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[0]_i_4 
       (.I0(bdatr[0]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[0]_i_5 
       (.I0(bdatr[8]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[0]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[0]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3]_i_11_n_7 ),
        .I2(\alu0/div/rem [0]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [0]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[0]_i_7 
       (.I0(\rgf_c0bus_wb[0]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c0bus_wb[0]_i_8 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[0]_i_15_n_0 ),
        .I5(\rgf_c0bus_wb[0]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAFBAA)) 
    \rgf_c0bus_wb[0]_i_9 
       (.I0(\rgf_c0bus_wb[0]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_19_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[10]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[10]),
        .I2(bdatr[10]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_3_n_0 ),
        .O(c0bus[10]));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[10]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[26]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[10]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h5030)) 
    \rgf_c0bus_wb[10]_i_11 
       (.I0(\rgf_c0bus_wb[27]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_18_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[10]_i_12 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \rgf_c0bus_wb[10]_i_13 
       (.I0(\rgf_c0bus_wb[18]_i_15_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c0bus_wb[10]_i_14 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[26]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[10]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \rgf_c0bus_wb[10]_i_16 
       (.I0(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c0bus_wb[10]_i_17 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[10]),
        .I2(b0bus_0[10]),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(a0bus_0[18]),
        .O(\rgf_c0bus_wb[10]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \rgf_c0bus_wb[10]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(a0bus_0[10]),
        .I2(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I4(b0bus_0[10]),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[10]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[10]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[10]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_67_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_70_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[10]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[9]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[10]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[10]_i_23 
       (.I0(\rgf_c0bus_wb[2]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h084C)) 
    \rgf_c0bus_wb[10]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[10]_i_25 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[9]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[10]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[10]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[10]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAEA)) 
    \rgf_c0bus_wb[10]_i_27 
       (.I0(\rgf_c0bus_wb[26]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I2(a0bus_0[10]),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(b0bus_0[10]),
        .O(\rgf_c0bus_wb[10]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hCFCFCFC055555555)) 
    \rgf_c0bus_wb[10]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I1(\alu0/asr0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul_a_i [17]),
        .I4(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[10]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [10]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[10]),
        .I4(\rgf_c0bus_wb[10]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[10]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[10]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBB00AF00AF00)) 
    \rgf_c0bus_wb[10]_i_5 
       (.I0(\rgf_c0bus_wb[10]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_14_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[10]_i_6 
       (.I0(\rgf_c0bus_wb[10]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_16_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[10]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_i_20_n_5 ),
        .I2(\alu0/div/rem [10]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [10]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h8FFF8F00)) 
    \rgf_c0bus_wb[10]_i_8 
       (.I0(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_18_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I4(\rgf_c0bus_wb_reg[10]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[10]_i_9 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[10]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[11]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[11]),
        .I2(bdatr[11]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_3_n_0 ),
        .O(c0bus[11]));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[11]_i_10 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[11]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[11]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c0bus_wb[11]_i_12 
       (.I0(\rgf_c0bus_wb[27]_i_33_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[11]_i_13 
       (.I0(\rgf_c0bus_wb[27]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[11]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[11]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[10]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[11]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[11]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[11]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[11]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c0bus_wb[11]_i_19 
       (.I0(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[11]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h5FC050C000000000)) 
    \rgf_c0bus_wb[11]_i_21 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[19]),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_33_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[11]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(b0bus_0[11]),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I4(a0bus_0[11]),
        .O(\rgf_c0bus_wb[11]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c0bus_wb[11]_i_23 
       (.I0(a0bus_0[3]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(a0bus_0[11]),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(b0bus_0[11]),
        .O(\rgf_c0bus_wb[11]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[11]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[11]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[11]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[11]_i_25 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c0bus_wb[11]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[11]_i_27 
       (.I0(\rgf_c0bus_wb[15]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[11]_i_28 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[10]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[11]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [11]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[11]),
        .I4(\rgf_c0bus_wb[11]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h5556555655555556)) 
    \rgf_c0bus_wb[11]_i_33 
       (.I0(a0bus_0[11]),
        .I1(p_2_in1_in[11]),
        .I2(\rgf/b0bus_out/bdatw[11]_INST_0_i_11_n_0 ),
        .I3(\rgf/b0bus_out/bdatw[11]_INST_0_i_10_n_0 ),
        .I4(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_36_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[11]_i_34 
       (.I0(\alu0/mul_a_i [17]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [18]),
        .I3(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[11]_i_35 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [11]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[11]));
  LUT6 #(
    .INIT(64'h5AAAAAAABBBBBBBB)) 
    \rgf_c0bus_wb[11]_i_36 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\fch/ir0 [10]),
        .I2(\bdatw[11]_INST_0_i_19_n_0 ),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [1]),
        .I5(ctl_selb0_0),
        .O(\rgf_c0bus_wb[11]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[11]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c0bus_wb[11]_i_5 
       (.I0(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_13_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[11]_i_6 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[11]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[11]_i_7 
       (.I0(\rgf_c0bus_wb[11]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[11]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_19_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[11]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_i_20_n_4 ),
        .I2(\alu0/div/rem [11]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [11]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[11]_i_9 
       (.I0(\rgf_c0bus_wb[11]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_22_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_23_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[12]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[12]),
        .I2(bdatr[12]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_3_n_0 ),
        .O(c0bus[12]));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[12]_i_10 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[12]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[12]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00EF00EF00FF0000)) 
    \rgf_c0bus_wb[12]_i_12 
       (.I0(\rgf_c0bus_wb[28]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[12]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[12]_i_14 
       (.I0(\rgf_c0bus_wb[28]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[12]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[11]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[12]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[12]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[12]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[12]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c0bus_wb[12]_i_19 
       (.I0(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[12]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[12]_i_20 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c0bus_wb[12]_i_21 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[12]),
        .I2(b0bus_0[12]),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(a0bus_0[20]),
        .O(\rgf_c0bus_wb[12]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \rgf_c0bus_wb[12]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(a0bus_0[12]),
        .I2(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I4(b0bus_0[12]),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[12]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_39_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c0bus_wb[12]_i_25 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[12]_i_26 
       (.I0(\rgf_c0bus_wb[12]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[12]_i_27 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[11]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[12]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[12]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[12]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c0bus_wb[12]_i_29 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(a0bus_0[12]),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(b0bus_0[12]),
        .O(\rgf_c0bus_wb[12]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[12]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [12]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[12]),
        .I4(\rgf_c0bus_wb[12]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[12]_i_30 
       (.I0(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'h888B8B8B)) 
    \rgf_c0bus_wb[12]_i_31 
       (.I0(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_45_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[12]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[12]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c0bus_wb[12]_i_5 
       (.I0(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[12]_i_6 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[12]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[12]_i_7 
       (.I0(\rgf_c0bus_wb[12]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_19_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[12]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_n_7 ),
        .I2(\alu0/div/rem [12]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [12]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h8FFF8F00)) 
    \rgf_c0bus_wb[12]_i_9 
       (.I0(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_22_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I4(\rgf_c0bus_wb_reg[12]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[13]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[13]),
        .I2(bdatr[13]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_3_n_0 ),
        .O(c0bus[13]));
  LUT6 #(
    .INIT(64'h4F444F4F4F444444)) 
    \rgf_c0bus_wb[13]_i_10 
       (.I0(\rgf_c0bus_wb[29]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I2(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[13]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[29]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00EF00EF00FF0000)) 
    \rgf_c0bus_wb[13]_i_12 
       (.I0(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[13]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h5030)) 
    \rgf_c0bus_wb[13]_i_14 
       (.I0(\rgf_c0bus_wb[30]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_19_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[13]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[12]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[13]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[13]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[13]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[13]_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[13]_i_19 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[13]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c0bus_wb[13]_i_20 
       (.I0(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h44C0CC0044C00000)) 
    \rgf_c0bus_wb[13]_i_21 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_29_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I5(a0bus_0[21]),
        .O(\rgf_c0bus_wb[13]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[13]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(b0bus_0[13]),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I4(a0bus_0[13]),
        .O(\rgf_c0bus_wb[13]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c0bus_wb[13]_i_23 
       (.I0(a0bus_0[5]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(b0bus_0[13]),
        .I4(a0bus_0[13]),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[13]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[13]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[13]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[13]_i_25 
       (.I0(\rgf_c0bus_wb[5]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c0bus_wb[13]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[13]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_64_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[13]_i_28 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[12]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h55555556)) 
    \rgf_c0bus_wb[13]_i_29 
       (.I0(a0bus_0[13]),
        .I1(p_2_in1_in[13]),
        .I2(\rgf/b0bus_out/bdatw[13]_INST_0_i_9_n_0 ),
        .I3(\rgf/b0bus_out/bdatw[13]_INST_0_i_8_n_0 ),
        .I4(\bdatw[13]_INST_0_i_7_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[13]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [13]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[13]),
        .I4(\rgf_c0bus_wb[13]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c0bus_wb[13]_i_30 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'h27FF2700)) 
    \rgf_c0bus_wb[13]_i_31 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[15]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[13]_i_32 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [13]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[13]));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[13]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c0bus_wb[13]_i_5 
       (.I0(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[13]_i_6 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[13]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[13]_i_7 
       (.I0(\rgf_c0bus_wb[13]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_20_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[13]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_n_6 ),
        .I2(\alu0/div/quo [13]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [13]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[13]_i_9 
       (.I0(\rgf_c0bus_wb[13]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_22_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[13]_i_23_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[13]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[14]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[14]),
        .I2(bdatr[14]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_3_n_0 ),
        .O(c0bus[14]));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c0bus_wb[14]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I3(a0bus_0[31]),
        .O(\rgf_c0bus_wb[14]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[14]_i_11 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FAFC0AFC)) 
    \rgf_c0bus_wb[14]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_43_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_15_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[14]_i_13 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c0bus_wb[14]_i_14 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h1DFF)) 
    \rgf_c0bus_wb[14]_i_15 
       (.I0(\rgf_c0bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h3808F8C800000000)) 
    \rgf_c0bus_wb[14]_i_16 
       (.I0(a0bus_0[22]),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_25_n_0 ),
        .I4(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[14]_i_17 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(b0bus_0[14]),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I4(a0bus_0[14]),
        .O(\rgf_c0bus_wb[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c0bus_wb[14]_i_18 
       (.I0(a0bus_0[6]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(b0bus_0[14]),
        .I4(a0bus_0[14]),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[14]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[14]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[14]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c0bus_wb[14]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[14]_i_20 
       (.I0(\rgf_c0bus_wb[30]_i_16_n_0 ),
        .I1(\remden[31]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[14]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[14]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[13]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[14]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c0bus_wb[14]_i_23 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[14]_i_24 
       (.I0(\rgf_c0bus_wb[30]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h55555556)) 
    \rgf_c0bus_wb[14]_i_25 
       (.I0(a0bus_0[14]),
        .I1(p_2_in1_in[14]),
        .I2(\rgf/b0bus_out/bdatw[14]_INST_0_i_10_n_0 ),
        .I3(\rgf/b0bus_out/bdatw[14]_INST_0_i_9_n_0 ),
        .I4(\bdatw[14]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFA0A0C0CFC0CF)) 
    \rgf_c0bus_wb[14]_i_26 
       (.I0(\rgf_c0bus_wb[20]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_38_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h15FF1500)) 
    \rgf_c0bus_wb[14]_i_27 
       (.I0(\rgf_c0bus_wb[30]_i_45_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[14]_i_28 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [14]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[14]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [14]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[14]),
        .I4(\rgf_c0bus_wb[14]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h8A88AAAA)) 
    \rgf_c0bus_wb[14]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFAF00BB00BB00)) 
    \rgf_c0bus_wb[14]_i_5 
       (.I0(\rgf_c0bus_wb[14]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_14_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hE2E200E2)) 
    \rgf_c0bus_wb[14]_i_6 
       (.I0(\rgf_c0bus_wb[14]_i_12_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_13_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c0bus_wb[14]_i_7 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[13]),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[14]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_n_5 ),
        .I2(\alu0/div/quo [14]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [14]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[14]_i_9 
       (.I0(\rgf_c0bus_wb[14]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_17_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_18_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[15]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[15]),
        .I2(bdatr[15]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_3_n_0 ),
        .O(c0bus[15]));
  LUT6 #(
    .INIT(64'hCFC0DFDFCFC0D0D0)) 
    \rgf_c0bus_wb[15]_i_10 
       (.I0(\rgf_c0bus_wb[15]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_21_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[15]_i_22_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[15]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFB51FB51FB11BB11)) 
    \rgf_c0bus_wb[15]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h08000888)) 
    \rgf_c0bus_wb[15]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFF70)) 
    \rgf_c0bus_wb[15]_i_14 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[14]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCDDCFCFFFDDCFCF)) 
    \rgf_c0bus_wb[15]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_44_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF8A80)) 
    \rgf_c0bus_wb[15]_i_16 
       (.I0(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_41_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_44_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_c0bus_wb[15]_i_18 
       (.I0(\rgf_c0bus_wb[31]_i_42_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c0bus_wb[15]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_5_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c0bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hDDCFDFFF)) 
    \rgf_c0bus_wb[15]_i_20 
       (.I0(b0bus_0[15]),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[15]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEFEEE00000000)) 
    \rgf_c0bus_wb[15]_i_21 
       (.I0(\rgf_c0bus_wb[15]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_35_n_0 ),
        .I3(b0bus_0[15]),
        .I4(a0bus_0[15]),
        .I5(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hBAAABABABAAABAAA)) 
    \rgf_c0bus_wb[15]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_57_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[15]),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(b0bus_0[15]),
        .O(\rgf_c0bus_wb[15]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[15]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[15]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[15]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c0bus_wb[15]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_25 
       (.I0(\rgf_c0bus_wb[28]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[15]_i_26 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[15]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_36_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[15]_i_28 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[14]),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[15]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [15]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[15]),
        .I4(\rgf_c0bus_wb[15]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8888888888888880)) 
    \rgf_c0bus_wb[15]_i_33 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(p_2_in1_in[7]),
        .I3(\rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[7]_INST_0_i_3_n_0 ),
        .I5(\bbus_o[7]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c0bus_wb[15]_i_34 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(a0bus_0[23]),
        .O(\rgf_c0bus_wb[15]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[15]_i_35 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hF022F077)) 
    \rgf_c0bus_wb[15]_i_36 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[15]),
        .I2(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h8A888A88AAAA8A88)) 
    \rgf_c0bus_wb[15]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_12_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hD000FFFFD000D000)) 
    \rgf_c0bus_wb[15]_i_5 
       (.I0(\rgf_c0bus_wb[15]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_13_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hA0AAEEEEA0AAE0EE)) 
    \rgf_c0bus_wb[15]_i_6 
       (.I0(\rgf_c0bus_wb[15]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_23_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[15]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c0bus_wb[15]_i_7 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c0bus_wb[15]_i_8 
       (.I0(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I1(\alu0/mul/mul_rslt ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[15]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[15]_i_19_n_4 ),
        .I2(\alu0/div/quo [15]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [15]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[16]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[16]),
        .I2(bdatr[16]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_3_n_0 ),
        .O(c0bus[16]));
  LUT6 #(
    .INIT(64'h5151514040405140)) 
    \rgf_c0bus_wb[16]_i_10 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(a0bus_0[31]),
        .I3(\rgf_c0bus_wb[23]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[16]_i_11 
       (.I0(\rgf_c0bus_wb[16]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hDDC8DDDDDDC88888)) 
    \rgf_c0bus_wb[16]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[16]_i_13 
       (.I0(\rgf_c0bus_wb[16]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c0bus_wb[16]_i_14 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[15]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c0bus_wb[16]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[16]_i_16 
       (.I0(\rgf_c0bus_wb[16]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_27_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h55015F01F501FF01)) 
    \rgf_c0bus_wb[16]_i_17 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_32_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c0bus_wb[16]_i_18 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[16]_i_19 
       (.I0(\rgf_c0bus_wb[16]_i_35_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_36_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[16]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[16]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[16]),
        .I2(a0bus_0[16]),
        .O(\rgf_c0bus_wb[16]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[16]_i_21 
       (.I0(a0bus_0[24]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[16]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[16]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[16]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[19]_i_11_n_7 ),
        .O(\rgf_c0bus_wb[16]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[16]_i_24 
       (.I0(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[17]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c0bus_wb[16]_i_25 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[16]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_62_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[16]_i_27 
       (.I0(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_56_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_52_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[16]_i_28 
       (.I0(\rgf_c0bus_wb[16]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \rgf_c0bus_wb[16]_i_29 
       (.I0(\rgf_c0bus_wb[7]_i_37_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[16]_i_3 
       (.I0(\rgf_c0bus_wb[16]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_9_n_0 ),
        .I2(niss_dsp_c0[16]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[16]_i_30 
       (.I0(\rgf_c0bus_wb[24]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[16]_i_31 
       (.I0(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[16]_i_32 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[16]_i_33 
       (.I0(\rgf_c0bus_wb[25]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[16]_i_34 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[15]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[16]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[16]_i_35 
       (.I0(a0bus_0[8]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[16]),
        .I4(a0bus_0[16]),
        .O(\rgf_c0bus_wb[16]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[16]_i_36 
       (.I0(a0bus_0[16]),
        .I1(b0bus_0[16]),
        .O(\rgf_c0bus_wb[16]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFD08)) 
    \rgf_c0bus_wb[16]_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[16]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[15]),
        .O(\rgf_c0bus_wb[16]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c0bus_wb[16]_i_38 
       (.I0(\rgf_c0bus_wb[22]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\alu0/mul_a_i [20]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\alu0/mul_a_i [21]),
        .I5(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hB8BBB8BBB8BBB888)) 
    \rgf_c0bus_wb[16]_i_39 
       (.I0(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\alu0/asr0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\alu0/mul_a_i [17]),
        .I5(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h8A88AAAA8A888A88)) 
    \rgf_c0bus_wb[16]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hF011F0DD)) 
    \rgf_c0bus_wb[16]_i_40 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[16]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000FF1010)) 
    \rgf_c0bus_wb[16]_i_5 
       (.I0(\rgf_c0bus_wb[16]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_16_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h545454FF55FF55FF)) 
    \rgf_c0bus_wb[16]_i_6 
       (.I0(\rgf_c0bus_wb[16]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_11_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_18_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[16]_i_7 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[16]_i_8 
       (.I0(\rgf_c0bus_wb[16]_i_19_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[16]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_23_n_0 ),
        .I2(\alu0/div/quo [16]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [16]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[16]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[17]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[17]),
        .I2(bdatr[17]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_3_n_0 ),
        .O(c0bus[17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[17]_i_10 
       (.I0(\rgf_c0bus_wb[25]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E2E2FFCC3300)) 
    \rgf_c0bus_wb[17]_i_11 
       (.I0(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[17]_i_12 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[16]),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[17]_i_13 
       (.I0(\rgf_c0bus_wb[25]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[17]_i_14 
       (.I0(\rgf_c0bus_wb[17]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E2E2FFCC3300)) 
    \rgf_c0bus_wb[17]_i_15 
       (.I0(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_c0bus_wb[17]_i_16 
       (.I0(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[17]_i_17 
       (.I0(\rgf_c0bus_wb[17]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[17]_i_18 
       (.I0(\rgf_c0bus_wb[17]_i_26_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_27_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[17]_i_19 
       (.I0(a0bus_0[25]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[17]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[17]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[17]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[17]),
        .I2(a0bus_0[17]),
        .O(\rgf_c0bus_wb[17]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[17]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[17]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[17]_i_22 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\alu0/art/add/tout [18]),
        .O(\rgf_c0bus_wb[17]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[17]_i_23 
       (.I0(\rgf_c0bus_wb[17]_i_28_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[17]_i_24 
       (.I0(\rgf_c0bus_wb[17]_i_30_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[17]_i_25 
       (.I0(\rgf_c0bus_wb[23]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[17]_i_31_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[17]_i_26 
       (.I0(a0bus_0[9]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[17]),
        .I4(a0bus_0[17]),
        .O(\rgf_c0bus_wb[17]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[17]_i_27 
       (.I0(a0bus_0[17]),
        .I1(b0bus_0[17]),
        .O(\rgf_c0bus_wb[17]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[17]_i_28 
       (.I0(a0bus_0[19]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[20]),
        .O(\rgf_c0bus_wb[17]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[17]_i_29 
       (.I0(a0bus_0[17]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[18]),
        .O(\rgf_c0bus_wb[17]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[17]_i_3 
       (.I0(\rgf_c0bus_wb[17]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_9_n_0 ),
        .I2(niss_dsp_c0[17]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[17]_i_30 
       (.I0(a0bus_0[20]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[19]),
        .O(\rgf_c0bus_wb[17]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[17]_i_31 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[19]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul_a_i [20]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[17]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[17]_i_32 
       (.I0(\alu0/mul_a_i [17]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [18]),
        .I3(\rgf/sreg/sr [8]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[17]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[17]_i_4 
       (.I0(\rgf_c0bus_wb[17]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEEEAAAEA)) 
    \rgf_c0bus_wb[17]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c0bus_wb[17]_i_6 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[17]_i_7 
       (.I0(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[17]_i_8 
       (.I0(\rgf_c0bus_wb[17]_i_18_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[17]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[17]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_22_n_0 ),
        .I2(\alu0/div/rem [17]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [17]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[17]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[18]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[18]),
        .I2(bdatr[18]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_3_n_0 ),
        .O(c0bus[18]));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[18]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_11 
       (.I0(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[18]_i_12 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\alu0/mul_a_i [17]),
        .O(\rgf_c0bus_wb[18]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[18]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[18]_i_14 
       (.I0(\rgf_c0bus_wb[18]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[18]_i_15 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_16 
       (.I0(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFB8FFFF)) 
    \rgf_c0bus_wb[18]_i_17 
       (.I0(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[18]_i_18 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[18]_i_19 
       (.I0(\rgf_c0bus_wb[18]_i_36_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_37_n_0 ),
        .I5(\rgf_c0bus_wb[26]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[18]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[18]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[18]),
        .I2(a0bus_0[18]),
        .O(\rgf_c0bus_wb[18]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[18]_i_21 
       (.I0(a0bus_0[26]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[18]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[18]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[18]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[19]_i_11_n_5 ),
        .O(\rgf_c0bus_wb[18]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[18]_i_24 
       (.I0(\rgf_c0bus_wb[30]_i_48_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_25 
       (.I0(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_51_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_43_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[18]_i_27 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_39_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[18]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[18]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[18]_i_3 
       (.I0(\rgf_c0bus_wb[18]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_9_n_0 ),
        .I2(niss_dsp_c0[18]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h8B8B88BB)) 
    \rgf_c0bus_wb[18]_i_30 
       (.I0(\rgf_c0bus_wb[30]_i_62_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(a0bus_0[18]),
        .I3(a0bus_0[17]),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[18]_i_31 
       (.I0(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_56_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_52_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[18]_i_32 
       (.I0(\rgf_c0bus_wb[20]_i_33_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[18]_i_33 
       (.I0(\rgf_c0bus_wb[20]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c0bus_wb[18]_i_34 
       (.I0(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\alu0/mul_a_i [26]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\alu0/mul_a_i [27]),
        .I5(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFEFF5400)) 
    \rgf_c0bus_wb[18]_i_35 
       (.I0(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I1(\alu0/mul_a_i [30]),
        .I2(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[18]_i_36 
       (.I0(a0bus_0[10]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[18]),
        .I4(a0bus_0[18]),
        .O(\rgf_c0bus_wb[18]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[18]_i_37 
       (.I0(a0bus_0[18]),
        .I1(b0bus_0[18]),
        .O(\rgf_c0bus_wb[18]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[18]_i_38 
       (.I0(a0bus_0[18]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[19]),
        .O(\rgf_c0bus_wb[18]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[18]_i_39 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[19]),
        .I2(\alu0/mul_a_i [18]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[18]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[18]_i_4 
       (.I0(\rgf_c0bus_wb[18]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[18]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[18]_i_6 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[18]_i_7 
       (.I0(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[18]_i_8 
       (.I0(\rgf_c0bus_wb[18]_i_19_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[18]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_23_n_0 ),
        .I2(\alu0/div/rem [18]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [18]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[18]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[19]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[19]),
        .I2(bdatr[19]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(p_2_in[19]),
        .O(c0bus[19]));
  LUT5 #(
    .INIT(32'hEEEEE000)) 
    \rgf_c0bus_wb[19]_i_10 
       (.I0(\rgf_c0bus_wb[19]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[19]_i_12 
       (.I0(\rgf_c0bus_wb[19]_i_31_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_32_n_0 ),
        .I5(\rgf_c0bus_wb[27]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[19]_i_13 
       (.I0(a0bus_0[27]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[19]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[19]),
        .I2(a0bus_0[19]),
        .O(\rgf_c0bus_wb[19]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[19]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[19]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[19]_i_16 
       (.I0(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[19]_i_17 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\alu0/mul_a_i [18]),
        .O(\rgf_c0bus_wb[19]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFF00E2E2)) 
    \rgf_c0bus_wb[19]_i_18 
       (.I0(\rgf_c0bus_wb[28]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[19]_i_19 
       (.I0(\rgf_c0bus_wb[27]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[19]_i_2 
       (.I0(\rgf_c0bus_wb[19]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .I2(niss_dsp_c0[19]),
        .I3(\rgf_c0bus_wb[19]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_5_n_0 ),
        .O(p_2_in[19]));
  LUT5 #(
    .INIT(32'h7FFF7F00)) 
    \rgf_c0bus_wb[19]_i_20 
       (.I0(a0bus_0[31]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[19]_i_21 
       (.I0(\rgf_c0bus_wb[19]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_c0bus_wb[19]_i_22 
       (.I0(\rgf_c0bus_wb[27]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[19]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[19]),
        .O(\rgf_c0bus_wb[19]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[19]_i_24 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[18]),
        .O(\rgf_c0bus_wb[19]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[19]_i_25 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[17]),
        .O(\rgf_c0bus_wb[19]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hD8)) 
    \rgf_c0bus_wb[19]_i_26 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[16]),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[19]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[19]_i_27 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[19]),
        .I2(b0bus_0[19]),
        .I3(\sr[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c0bus_wb[19]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[19]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[19]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[19]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[19]_i_31 
       (.I0(a0bus_0[11]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[19]),
        .I4(a0bus_0[19]),
        .O(\rgf_c0bus_wb[19]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[19]_i_32 
       (.I0(a0bus_0[19]),
        .I1(b0bus_0[19]),
        .O(\rgf_c0bus_wb[19]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[19]_i_33 
       (.I0(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_41_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[19]_i_34 
       (.I0(\remden[31]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[19]_i_4 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb_reg[19]_i_11_n_4 ),
        .I2(\alu0/div/quo [19]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [19]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[19]_i_5 
       (.I0(\rgf_c0bus_wb[19]_i_12_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[19]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[19]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[19]_i_6 
       (.I0(\rgf_c0bus_wb[2]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[19]_i_7 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[19]_i_8 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[19]_i_9 
       (.I0(\rgf_c0bus_wb[19]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[1]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[1]),
        .I2(\rgf_c0bus_wb[1]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_5_n_0 ),
        .O(c0bus[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFF45444545)) 
    \rgf_c0bus_wb[1]_i_10 
       (.I0(\rgf_c0bus_wb[1]_i_19_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[17]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[1]_i_11 
       (.I0(a0bus_0[25]),
        .I1(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c0bus_wb[1]_i_12 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(a0bus_0[1]),
        .I3(a0bus_0[9]),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[1]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(a0bus_0[1]),
        .I3(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[1]_i_14 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[1]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[17]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[1]_i_16 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c0bus_wb[1]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_26_n_0 ),
        .I4(a0bus_0[0]),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFD50000)) 
    \rgf_c0bus_wb[1]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_31_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF04C404C404C4)) 
    \rgf_c0bus_wb[1]_i_19 
       (.I0(\rgf_c0bus_wb[17]_i_14_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_23_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[1]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [1]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[1]),
        .I4(\rgf_c0bus_wb[1]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \rgf_c0bus_wb[1]_i_20 
       (.I0(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \rgf_c0bus_wb[1]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000021333330213)) 
    \rgf_c0bus_wb[1]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c0bus_wb[1]_i_23 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[1]_i_24 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[1]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[1]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[1]_i_4 
       (.I0(bdatr[1]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[1]_i_5 
       (.I0(bdatr[9]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[1]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[1]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3]_i_11_n_6 ),
        .I2(\alu0/div/quo [1]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [1]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[1]_i_7 
       (.I0(\rgf_c0bus_wb[1]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[1]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[1]_i_8 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[1]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[1]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h000000F2)) 
    \rgf_c0bus_wb[1]_i_9 
       (.I0(\rgf_c0bus_wb[1]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[1]_i_17_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[1]_i_18_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[20]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[20]),
        .I2(bdatr[20]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_3_n_0 ),
        .O(c0bus[20]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[20]_i_10 
       (.I0(\rgf_c0bus_wb[28]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_22_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[20]_i_11 
       (.I0(\rgf_c0bus_wb[20]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[20]_i_12 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[19]),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFCC3300B8B8B8B8)) 
    \rgf_c0bus_wb[20]_i_13 
       (.I0(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[20]_i_14 
       (.I0(\rgf_c0bus_wb[28]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[20]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[20]_i_16 
       (.I0(\rgf_c0bus_wb[20]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B8FFFFFFFF)) 
    \rgf_c0bus_wb[20]_i_17 
       (.I0(\rgf_c0bus_wb[20]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[20]_i_18 
       (.I0(\rgf_c0bus_wb[20]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\remden[31]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[20]_i_19 
       (.I0(\rgf_c0bus_wb[20]_i_31_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_32_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[20]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[20]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[20]_i_20 
       (.I0(a0bus_0[28]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[20]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[20]),
        .I2(a0bus_0[20]),
        .O(\rgf_c0bus_wb[20]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[20]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[20]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[20]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[23]_i_24_n_7 ),
        .O(\rgf_c0bus_wb[20]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[20]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_50_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_51_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[20]_i_25 
       (.I0(\rgf_c0bus_wb[22]_i_29_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[20]_i_26 
       (.I0(\rgf_c0bus_wb[22]_i_31_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c0bus_wb[20]_i_27 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[20]_i_28 
       (.I0(a0bus_0[4]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[20]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[20]_i_29 
       (.I0(a0bus_0[2]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[20]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[20]_i_3 
       (.I0(\rgf_c0bus_wb[20]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_9_n_0 ),
        .I2(niss_dsp_c0[20]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[20]_i_30 
       (.I0(\rgf_c0bus_wb[22]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[20]_i_31 
       (.I0(a0bus_0[12]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[20]),
        .I4(a0bus_0[20]),
        .O(\rgf_c0bus_wb[20]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[20]_i_32 
       (.I0(a0bus_0[20]),
        .I1(b0bus_0[20]),
        .O(\rgf_c0bus_wb[20]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[20]_i_33 
       (.I0(a0bus_0[20]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[21]),
        .O(\rgf_c0bus_wb[20]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[20]_i_34 
       (.I0(\alu0/mul_a_i [20]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [21]),
        .I3(\rgf/sreg/sr [8]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[20]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[20]_i_4 
       (.I0(\rgf_c0bus_wb[20]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[20]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[20]_i_6 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[20]_i_7 
       (.I0(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[20]_i_8 
       (.I0(\rgf_c0bus_wb[20]_i_19_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[20]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[20]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_23_n_0 ),
        .I2(\alu0/div/quo [20]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [20]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[21]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[21]),
        .I2(bdatr[21]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[21]_i_3_n_0 ),
        .O(c0bus[21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_10 
       (.I0(\rgf_c0bus_wb[21]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_11 
       (.I0(\rgf_c0bus_wb[21]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[21]_i_12 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\alu0/mul_a_i [20]),
        .O(\rgf_c0bus_wb[21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF33CC00E2E2E2E2)) 
    \rgf_c0bus_wb[21]_i_13 
       (.I0(\rgf_c0bus_wb[30]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_27_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_14 
       (.I0(\rgf_c0bus_wb[21]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[21]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_16 
       (.I0(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hEFECE3E0FFFFFFFF)) 
    \rgf_c0bus_wb[21]_i_17 
       (.I0(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_33_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000CDC8CDC8)) 
    \rgf_c0bus_wb[21]_i_18 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\remden[31]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_35_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[21]_i_19 
       (.I0(\rgf_c0bus_wb[21]_i_36_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_37_n_0 ),
        .I5(\rgf_c0bus_wb[29]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[21]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[21]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[21]),
        .I2(a0bus_0[21]),
        .O(\rgf_c0bus_wb[21]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[21]_i_21 
       (.I0(a0bus_0[29]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[21]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[21]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[21]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_67_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_68_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[21]_i_24 
       (.I0(\rgf_c0bus_wb[25]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[21]_i_25 
       (.I0(\rgf_c0bus_wb[31]_i_64_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c0bus_wb[21]_i_26 
       (.I0(a0bus_0[31]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[21]_i_27 
       (.I0(\rgf_c0bus_wb[21]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[21]_i_28 
       (.I0(\rgf_c0bus_wb[25]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_53_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[21]_i_29 
       (.I0(\rgf_c0bus_wb[31]_i_76_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_72_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_73_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[21]_i_3 
       (.I0(\rgf_c0bus_wb[21]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_9_n_0 ),
        .I2(niss_dsp_c0[21]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF777700037774)) 
    \rgf_c0bus_wb[21]_i_30 
       (.I0(a0bus_0[31]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[21]_i_31 
       (.I0(\rgf_c0bus_wb[23]_i_40_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[21]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[21]_i_32 
       (.I0(a0bus_0[5]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[21]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[21]_i_33 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[21]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[21]_i_34 
       (.I0(\alu0/mul_a_i [29]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [30]),
        .I3(\rgf/sreg/sr [8]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[21]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[21]_i_35 
       (.I0(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_41_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[21]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[21]_i_36 
       (.I0(a0bus_0[13]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[21]),
        .I4(a0bus_0[21]),
        .O(\rgf_c0bus_wb[21]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[21]_i_37 
       (.I0(a0bus_0[21]),
        .I1(b0bus_0[21]),
        .O(\rgf_c0bus_wb[21]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[21]_i_38 
       (.I0(a0bus_0[21]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[22]),
        .O(\rgf_c0bus_wb[21]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[21]_i_39 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[22]),
        .I2(\alu0/mul_a_i [21]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[21]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[21]_i_4 
       (.I0(\rgf_c0bus_wb[21]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[21]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[21]_i_6 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[21]_i_7 
       (.I0(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[21]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[21]_i_8 
       (.I0(\rgf_c0bus_wb[21]_i_19_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[21]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[21]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb_reg[23]_i_24_n_6 ),
        .I2(\alu0/div/rem [21]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [21]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[21]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[22]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[22]),
        .I2(bdatr[22]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_3_n_0 ),
        .O(c0bus[22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_10 
       (.I0(\rgf_c0bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[22]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_26_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[22]_i_12 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\alu0/mul_a_i [21]),
        .O(\rgf_c0bus_wb[22]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \rgf_c0bus_wb[22]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_14 
       (.I0(\rgf_c0bus_wb[30]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[22]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_16 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \rgf_c0bus_wb[22]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_37_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_36_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[22]_i_18 
       (.I0(\rgf_c0bus_wb[22]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \rgf_c0bus_wb[22]_i_19 
       (.I0(\rgf_c0bus_wb[22]_i_27_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[22]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[22]_i_20 
       (.I0(a0bus_0[30]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[22]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[22]),
        .I2(a0bus_0[22]),
        .O(\rgf_c0bus_wb[22]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[22]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[22]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[22]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[23]_i_24_n_5 ),
        .O(\rgf_c0bus_wb[22]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[22]_i_24 
       (.I0(\rgf_c0bus_wb[28]_i_44_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[22]_i_25 
       (.I0(\rgf_c0bus_wb[22]_i_30_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[22]_i_26 
       (.I0(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_33_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[22]_i_27 
       (.I0(a0bus_0[14]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[22]),
        .I4(a0bus_0[22]),
        .O(\rgf_c0bus_wb[22]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[22]_i_28 
       (.I0(a0bus_0[22]),
        .I1(b0bus_0[22]),
        .O(\rgf_c0bus_wb[22]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[22]_i_29 
       (.I0(a0bus_0[26]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[27]),
        .O(\rgf_c0bus_wb[22]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[22]_i_3 
       (.I0(\rgf_c0bus_wb[22]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_9_n_0 ),
        .I2(niss_dsp_c0[22]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[22]_i_30 
       (.I0(a0bus_0[25]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[24]),
        .O(\rgf_c0bus_wb[22]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[22]_i_31 
       (.I0(a0bus_0[22]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[23]),
        .O(\rgf_c0bus_wb[22]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB8B8)) 
    \rgf_c0bus_wb[22]_i_32 
       (.I0(\alu0/mul_a_i [26]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [27]),
        .I3(\rgf/sreg/sr [8]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[22]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hDDF588A0)) 
    \rgf_c0bus_wb[22]_i_33 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[24]),
        .I2(a0bus_0[25]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[22]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hDDF588A0)) 
    \rgf_c0bus_wb[22]_i_34 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[22]),
        .I2(a0bus_0[23]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[22]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[22]_i_4 
       (.I0(\rgf_c0bus_wb[22]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[22]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c0bus_wb[22]_i_6 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c0bus_wb[22]_i_7 
       (.I0(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[22]_i_8 
       (.I0(\rgf_c0bus_wb[22]_i_19_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[22]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_23_n_0 ),
        .I2(\alu0/div/rem [22]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [22]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[22]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[23]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[23]),
        .I2(bdatr[23]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_3_n_0 ),
        .O(c0bus[23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_10 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[23]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[23]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_46_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000BBBBBBBB)) 
    \rgf_c0bus_wb[23]_i_13 
       (.I0(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[23]_i_14 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_15 
       (.I0(\rgf_c0bus_wb[23]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rgf_c0bus_wb[23]_i_17 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_39_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[23]_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[22]),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[23]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[23]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[23]_i_20 
       (.I0(\rgf_c0bus_wb[23]_i_30_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_31_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_60_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[23]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[23]),
        .I2(a0bus_0[23]),
        .O(\rgf_c0bus_wb[23]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[23]_i_22 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[23]_i_23 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[23]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c0bus_wb[23]_i_25 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[23]_i_26 
       (.I0(\rgf_c0bus_wb[25]_i_42_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[23]_i_27 
       (.I0(\rgf_c0bus_wb[25]_i_41_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_40_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[23]_i_28 
       (.I0(\rgf_c0bus_wb[21]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \rgf_c0bus_wb[23]_i_29 
       (.I0(\rgf_c0bus_wb[27]_i_45_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[23]_i_3 
       (.I0(\rgf_c0bus_wb[23]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_9_n_0 ),
        .I2(niss_dsp_c0[23]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[23]_i_30 
       (.I0(a0bus_0[15]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[23]),
        .I4(a0bus_0[23]),
        .O(\rgf_c0bus_wb[23]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[23]_i_31 
       (.I0(a0bus_0[23]),
        .I1(b0bus_0[23]),
        .O(\rgf_c0bus_wb[23]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_32 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[23]),
        .O(\rgf_c0bus_wb[23]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_33 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[22]),
        .O(\rgf_c0bus_wb[23]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_34 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[21]),
        .O(\rgf_c0bus_wb[23]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[23]_i_35 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[20]),
        .O(\rgf_c0bus_wb[23]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[23]_i_36 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[23]),
        .I2(b0bus_0[23]),
        .I3(\sr[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[23]_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[22]),
        .I2(b0bus_0[22]),
        .I3(\sr[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h0111011101115555)) 
    \rgf_c0bus_wb[23]_i_4 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_11_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[23]_i_40 
       (.I0(a0bus_0[23]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[24]),
        .O(\rgf_c0bus_wb[23]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hDDF588A0)) 
    \rgf_c0bus_wb[23]_i_41 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[23]),
        .I2(a0bus_0[24]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[23]_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hCF88CF8F)) 
    \rgf_c0bus_wb[23]_i_5 
       (.I0(\rgf_c0bus_wb[23]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFB8)) 
    \rgf_c0bus_wb[23]_i_6 
       (.I0(\rgf_c0bus_wb[23]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[23]_i_7 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[23]_i_8 
       (.I0(\rgf_c0bus_wb[23]_i_20_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[23]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb_reg[23]_i_24_n_4 ),
        .I2(\alu0/div/rem [23]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [23]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[23]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[24]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[24]),
        .I2(bdatr[24]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(p_2_in[24]),
        .O(c0bus[24]));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[24]_i_10 
       (.I0(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[24]_i_11 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_7 ),
        .O(\rgf_c0bus_wb[24]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBFFBBBBBBCC88888)) 
    \rgf_c0bus_wb[24]_i_12 
       (.I0(\rgf_c0bus_wb[24]_i_24_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(a0bus_0[24]),
        .I3(b0bus_0[24]),
        .I4(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[24]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[24]),
        .I2(a0bus_0[24]),
        .O(\rgf_c0bus_wb[24]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[24]_i_14 
       (.I0(a0bus_0[16]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[24]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I3(a0bus_0[24]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h5C)) 
    \rgf_c0bus_wb[24]_i_16 
       (.I0(\rgf_c0bus_wb[7]_i_37_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_17 
       (.I0(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[24]_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[23]),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_19 
       (.I0(\rgf_c0bus_wb[16]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[24]_i_2 
       (.I0(\rgf_c0bus_wb[24]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .I2(niss_dsp_c0[24]),
        .I3(\rgf_c0bus_wb[24]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[24]_i_5_n_0 ),
        .O(p_2_in[24]));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[24]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[24]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[24]_i_21 
       (.I0(\rgf_c0bus_wb[28]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I4(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_22 
       (.I0(\rgf_c0bus_wb[28]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \rgf_c0bus_wb[24]_i_23 
       (.I0(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I1(a0bus_0[0]),
        .I2(\rgf_c0bus_wb[16]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[24]_i_24 
       (.I0(a0bus_0[0]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[24]_i_25 
       (.I0(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[24]_i_26 
       (.I0(\rgf_c0bus_wb[28]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[24]_i_27 
       (.I0(\rgf_c0bus_wb[20]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_52_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_28 
       (.I0(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_62_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[24]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c0bus_wb[24]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[24]_i_9_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[24]_i_30 
       (.I0(\alu0/mul_a_i [26]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [27]),
        .I3(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[22]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[24]_i_4 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_11_n_0 ),
        .I2(\alu0/div/quo [24]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [24]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \rgf_c0bus_wb[24]_i_5 
       (.I0(\rgf_c0bus_wb[24]_i_12_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_14_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[24]_i_6 
       (.I0(\rgf_c0bus_wb[24]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[24]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[24]_i_7 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[24]_i_8 
       (.I0(\rgf_c0bus_wb[24]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \rgf_c0bus_wb[24]_i_9 
       (.I0(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[24]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[25]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[25]),
        .I2(bdatr[25]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_3_n_0 ),
        .O(c0bus[25]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_10 
       (.I0(\rgf_c0bus_wb[25]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \rgf_c0bus_wb[25]_i_11 
       (.I0(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[25]_i_12 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[24]),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_13 
       (.I0(\rgf_c0bus_wb[25]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rgf_c0bus_wb[25]_i_14 
       (.I0(\rgf_c0bus_wb[25]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_32_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_15 
       (.I0(\rgf_c0bus_wb[25]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFF00FEFE)) 
    \rgf_c0bus_wb[25]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[25]_i_17 
       (.I0(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_36_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[25]_i_18 
       (.I0(\rgf_c0bus_wb[25]_i_37_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_38_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[25]_i_19 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[25]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[25]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[25]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[25]),
        .I2(a0bus_0[25]),
        .O(\rgf_c0bus_wb[25]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[25]_i_21 
       (.I0(a0bus_0[17]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[25]_i_22 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_6 ),
        .O(\rgf_c0bus_wb[25]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_67_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_68_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_24 
       (.I0(\rgf_c0bus_wb[20]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_25 
       (.I0(\rgf_c0bus_wb[25]_i_40_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_26 
       (.I0(\rgf_c0bus_wb[27]_i_44_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_64_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_28 
       (.I0(\rgf_c0bus_wb[21]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_76_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_72_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[25]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_43_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[25]_i_3 
       (.I0(\rgf_c0bus_wb[25]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_9_n_0 ),
        .I2(niss_dsp_c0[25]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_30 
       (.I0(\rgf_c0bus_wb[31]_i_54_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_55_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_31 
       (.I0(\rgf_c0bus_wb[31]_i_56_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_48_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[25]_i_32 
       (.I0(\rgf_c0bus_wb[31]_i_73_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c0bus_wb[25]_i_33 
       (.I0(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(a0bus_0[17]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[16]),
        .O(\rgf_c0bus_wb[25]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[25]_i_34 
       (.I0(\remden[31]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[25]_i_35 
       (.I0(a0bus_0[1]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[0]),
        .O(\rgf_c0bus_wb[25]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hB8FF)) 
    \rgf_c0bus_wb[25]_i_36 
       (.I0(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[25]_i_37 
       (.I0(a0bus_0[1]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[25]),
        .I4(a0bus_0[25]),
        .O(\rgf_c0bus_wb[25]_i_37_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[25]_i_38 
       (.I0(a0bus_0[25]),
        .I1(b0bus_0[25]),
        .O(\rgf_c0bus_wb[25]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[25]_i_39 
       (.I0(\rgf_c0bus_wb[18]_i_38_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_70_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[25]_i_4 
       (.I0(\rgf_c0bus_wb[25]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[25]_i_40 
       (.I0(a0bus_0[27]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[28]),
        .O(\rgf_c0bus_wb[25]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[25]_i_41 
       (.I0(a0bus_0[25]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[26]),
        .O(\rgf_c0bus_wb[25]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[25]_i_42 
       (.I0(a0bus_0[29]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[25]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[25]_i_43 
       (.I0(a0bus_0[31]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[25]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[25]_i_44 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[25]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul_a_i [26]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[25]_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[25]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[25]_i_6 
       (.I0(\rgf_c0bus_wb[25]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c0bus_wb[25]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hACAFACAFACAFA0A3)) 
    \rgf_c0bus_wb[25]_i_8 
       (.I0(\rgf_c0bus_wb[25]_i_18_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[25]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_22_n_0 ),
        .I2(\alu0/div/quo [25]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [25]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[25]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[26]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[26]),
        .I2(bdatr[26]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(p_2_in[26]),
        .O(c0bus[26]));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[26]_i_10 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_5 ),
        .O(\rgf_c0bus_wb[26]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBFFBBBBBBCC88888)) 
    \rgf_c0bus_wb[26]_i_11 
       (.I0(\rgf_c0bus_wb[26]_i_23_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(a0bus_0[26]),
        .I3(b0bus_0[26]),
        .I4(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I5(\rgf_c0bus_wb[26]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[26]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[26]),
        .I2(a0bus_0[26]),
        .O(\rgf_c0bus_wb[26]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[26]_i_13 
       (.I0(a0bus_0[18]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[26]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I3(a0bus_0[26]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFCC3300E2E2E2E2)) 
    \rgf_c0bus_wb[26]_i_15 
       (.I0(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[26]_i_16 
       (.I0(\rgf_c0bus_wb[18]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[26]_i_17 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[25]),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[26]_i_18 
       (.I0(\rgf_c0bus_wb[18]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \rgf_c0bus_wb[26]_i_19 
       (.I0(\rgf_c0bus_wb[17]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[26]_i_2 
       (.I0(\rgf_c0bus_wb[26]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .I2(niss_dsp_c0[26]),
        .I3(\rgf_c0bus_wb[26]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_5_n_0 ),
        .O(p_2_in[26]));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[26]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_35_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FEAEFEAE)) 
    \rgf_c0bus_wb[26]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_31_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000B8FF0000)) 
    \rgf_c0bus_wb[26]_i_22 
       (.I0(\rgf_c0bus_wb[30]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[26]_i_23 
       (.I0(a0bus_0[2]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[26]_i_24 
       (.I0(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[26]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[26]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[26]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[26]_i_4 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_10_n_0 ),
        .I2(\alu0/div/quo [26]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [26]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \rgf_c0bus_wb[26]_i_5 
       (.I0(\rgf_c0bus_wb[26]_i_11_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[26]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[26]_i_13_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[26]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[26]_i_6 
       (.I0(\rgf_c0bus_wb[26]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[26]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[26]_i_7 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[26]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[26]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[26]_i_8 
       (.I0(\rgf_c0bus_wb[26]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c0bus_wb[26]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[26]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[26]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[26]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[27]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[27]),
        .I2(bdatr[27]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[27]_i_3_n_0 ),
        .O(c0bus[27]));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[27]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_11 
       (.I0(\rgf_c0bus_wb[27]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[27]_i_12 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\alu0/mul_a_i [26]),
        .O(\rgf_c0bus_wb[27]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_13 
       (.I0(\rgf_c0bus_wb[27]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[27]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hEF40)) 
    \rgf_c0bus_wb[27]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \rgf_c0bus_wb[27]_i_16 
       (.I0(\rgf_c0bus_wb[27]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAAA7555)) 
    \rgf_c0bus_wb[27]_i_17 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[27]_i_18 
       (.I0(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[27]_i_19 
       (.I0(\rgf_c0bus_wb[27]_i_34_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_35_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[27]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[27]_i_20 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[27]),
        .I2(a0bus_0[27]),
        .O(\rgf_c0bus_wb[27]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[27]_i_21 
       (.I0(a0bus_0[19]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[27]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[27]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_67_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c0bus_wb[27]_i_25 
       (.I0(a0bus_0[17]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[16]),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[27]_i_26 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[27]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_68_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_64_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[27]_i_28 
       (.I0(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_76_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_72_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_73_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \rgf_c0bus_wb[27]_i_29 
       (.I0(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_33_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_45_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[27]_i_3 
       (.I0(\rgf_c0bus_wb[27]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_9_n_0 ),
        .I2(niss_dsp_c0[27]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[27]_i_30 
       (.I0(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[27]_i_31 
       (.I0(\alu0/mul_a_i [29]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [30]),
        .I3(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[27]_i_46_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[27]_i_32 
       (.I0(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h2EEEEEEEFFFFFFFF)) 
    \rgf_c0bus_wb[27]_i_33 
       (.I0(\rgf_c0bus_wb[23]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[31]),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[27]_i_34 
       (.I0(a0bus_0[3]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[27]),
        .I4(a0bus_0[27]),
        .O(\rgf_c0bus_wb[27]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[27]_i_35 
       (.I0(a0bus_0[27]),
        .I1(b0bus_0[27]),
        .O(\rgf_c0bus_wb[27]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_36 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[27]),
        .O(\rgf_c0bus_wb[27]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[26]),
        .O(\rgf_c0bus_wb[27]_i_37_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_38 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[25]),
        .O(\rgf_c0bus_wb[27]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[27]_i_39 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[24]),
        .O(\rgf_c0bus_wb[27]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[27]_i_4 
       (.I0(\rgf_c0bus_wb[27]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[27]_i_42 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[25]),
        .I2(b0bus_0[25]),
        .I3(\sr[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_42_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[27]_i_43 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[24]),
        .I2(b0bus_0[24]),
        .I3(\sr[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[27]_i_44 
       (.I0(a0bus_0[31]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[27]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[27]_i_45 
       (.I0(\rgf_c0bus_wb[30]_i_59_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[25]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[27]_i_46 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[28]),
        .I2(\alu0/mul_a_i [27]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[27]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[27]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[27]_i_6 
       (.I0(\rgf_c0bus_wb[27]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c0bus_wb[27]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[27]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[27]_i_8 
       (.I0(\rgf_c0bus_wb[27]_i_19_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_21_n_0 ),
        .I5(\rgf_c0bus_wb[27]_i_22_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[27]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_4 ),
        .I2(\alu0/div/rem [27]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [27]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[28]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[28]),
        .I2(bdatr[28]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_3_n_0 ),
        .O(c0bus[28]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[28]_i_10 
       (.I0(\rgf_c0bus_wb[28]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_11 
       (.I0(\rgf_c0bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[28]_i_12 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\alu0/mul_a_i [27]),
        .O(\rgf_c0bus_wb[28]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[28]_i_13 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \rgf_c0bus_wb[28]_i_14 
       (.I0(\rgf_c0bus_wb[28]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_31_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hEF40)) 
    \rgf_c0bus_wb[28]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCFCAC5C0CFCACFCA)) 
    \rgf_c0bus_wb[28]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I5(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \rgf_c0bus_wb[28]_i_17 
       (.I0(\rgf_c0bus_wb[28]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[28]_i_18 
       (.I0(\rgf_c0bus_wb[28]_i_36_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_37_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[28]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[28]),
        .I2(a0bus_0[28]),
        .O(\rgf_c0bus_wb[28]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[28]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[28]_i_20 
       (.I0(a0bus_0[20]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[28]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[28]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \rgf_c0bus_wb[28]_i_22 
       (.I0(a0bus_0[17]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[18]),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_43_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_23 
       (.I0(\rgf_c0bus_wb[30]_i_44_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_24 
       (.I0(\rgf_c0bus_wb[23]_i_27_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[28]_i_25 
       (.I0(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_39_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[28]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_51_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_48_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[28]_i_27 
       (.I0(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_56_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_52_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[28]_i_28 
       (.I0(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h5F5030305F503F30)) 
    \rgf_c0bus_wb[28]_i_29 
       (.I0(a0bus_0[31]),
        .I1(a0bus_0[30]),
        .I2(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[28]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[28]_i_3 
       (.I0(\rgf_c0bus_wb[28]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_9_n_0 ),
        .I2(niss_dsp_c0[28]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_30 
       (.I0(\rgf_c0bus_wb[30]_i_61_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_58_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_31 
       (.I0(\rgf_c0bus_wb[28]_i_40_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_60_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \rgf_c0bus_wb[28]_i_32 
       (.I0(\rgf_c0bus_wb[28]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_62_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0FFFFEFE00000)) 
    \rgf_c0bus_wb[28]_i_33 
       (.I0(\alu0/mul_a_i [30]),
        .I1(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\remden[31]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[28]_i_34 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[0]),
        .O(\rgf_c0bus_wb[28]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_35 
       (.I0(\rgf_c0bus_wb[28]_i_43_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[28]_i_36 
       (.I0(a0bus_0[4]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[28]),
        .I4(a0bus_0[28]),
        .O(\rgf_c0bus_wb[28]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[28]_i_37 
       (.I0(a0bus_0[28]),
        .I1(b0bus_0[28]),
        .O(\rgf_c0bus_wb[28]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_38 
       (.I0(\rgf_c0bus_wb[21]_i_38_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[28]_i_39 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[28]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[28]_i_4 
       (.I0(\rgf_c0bus_wb[28]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[28]_i_40 
       (.I0(a0bus_0[22]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[21]),
        .O(\rgf_c0bus_wb[28]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[28]_i_41 
       (.I0(\rgf_c0bus_wb[30]_i_63_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[17]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[28]_i_42 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[28]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul_a_i [29]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[28]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[28]_i_43 
       (.I0(a0bus_0[31]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[28]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[28]_i_44 
       (.I0(a0bus_0[29]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[28]),
        .O(\rgf_c0bus_wb[28]_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[28]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[28]_i_6 
       (.I0(\rgf_c0bus_wb[28]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c0bus_wb[28]_i_7 
       (.I0(\rgf_c0bus_wb[28]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B888BBBBBB8B)) 
    \rgf_c0bus_wb[28]_i_8 
       (.I0(\rgf_c0bus_wb[28]_i_18_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[28]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb_reg[29]_i_11_n_7 ),
        .I2(\alu0/div/rem [28]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo__0 [28]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[28]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF88F8)) 
    \rgf_c0bus_wb[29]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[29]),
        .I2(bdatr[29]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(p_2_in[29]),
        .O(c0bus[29]));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[29]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[29]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c0bus_wb[29]_i_12 
       (.I0(\rgf_c0bus_wb[29]_i_32_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_33_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[29]_i_13 
       (.I0(a0bus_0[21]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c0bus_wb[29]_i_14 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[29]),
        .I2(a0bus_0[29]),
        .O(\rgf_c0bus_wb[29]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \rgf_c0bus_wb[29]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[29]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[29]_i_16 
       (.I0(\rgf_c0bus_wb[21]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[29]_i_17 
       (.I0(\rgf_c0bus_wb[21]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c0bus_wb[29]_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[28]),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[29]_i_19 
       (.I0(\rgf_c0bus_wb[21]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \rgf_c0bus_wb[29]_i_2 
       (.I0(\rgf_c0bus_wb[29]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .I2(niss_dsp_c0[29]),
        .I3(\rgf_c0bus_wb[29]_i_4_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_5_n_0 ),
        .O(p_2_in[29]));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[29]_i_20 
       (.I0(\rgf_c0bus_wb[25]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_24_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hEF40)) 
    \rgf_c0bus_wb[29]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[29]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \rgf_c0bus_wb[29]_i_23 
       (.I0(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_24 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .O(\rgf_c0bus_wb[29]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_25 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[30]),
        .O(\rgf_c0bus_wb[29]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_26 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[29]),
        .O(\rgf_c0bus_wb[29]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[29]_i_27 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[28]),
        .O(\rgf_c0bus_wb[29]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \rgf_c0bus_wb[29]_i_28 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(\alu0/art/p_0_in__0 ),
        .O(\rgf_c0bus_wb[29]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[29]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[29]_i_6_n_0 ),
        .I2(\rgf_c0bus_wb[29]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[29]_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c0bus_wb[29]_i_31 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[28]),
        .I2(b0bus_0[28]),
        .I3(\sr[6]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[29]_i_32 
       (.I0(a0bus_0[5]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[29]),
        .I4(a0bus_0[29]),
        .O(\rgf_c0bus_wb[29]_i_32_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[29]_i_33 
       (.I0(a0bus_0[29]),
        .I1(b0bus_0[29]),
        .O(\rgf_c0bus_wb[29]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c0bus_wb[29]_i_34 
       (.I0(\remden[31]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\alu0/mul_a_i [29]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\alu0/mul_a_i [30]),
        .I5(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[29]_i_4 
       (.I0(\rgf_c0bus_wb[29]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb_reg[29]_i_11_n_6 ),
        .I2(\alu0/div/quo__0 [29]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [29]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB888B8B8BB8BBBBB)) 
    \rgf_c0bus_wb[29]_i_5 
       (.I0(\rgf_c0bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[29]_i_13_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_14_n_0 ),
        .I5(\rgf_c0bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[29]_i_6 
       (.I0(\rgf_c0bus_wb[29]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[29]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[29]_i_7 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[29]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[29]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[29]_i_8 
       (.I0(\rgf_c0bus_wb[29]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c0bus_wb[29]_i_9 
       (.I0(\rgf_c0bus_wb[29]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[29]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[29]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[29]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEFE)) 
    \rgf_c0bus_wb[2]_i_1 
       (.I0(\rgf_c0bus_wb[2]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_7_n_0 ),
        .O(c0bus[2]));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \rgf_c0bus_wb[2]_i_10 
       (.I0(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h002E002E0000002E)) 
    \rgf_c0bus_wb[2]_i_11 
       (.I0(\rgf_c0bus_wb[2]_i_19_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c0bus_wb[2]_i_12 
       (.I0(\rgf_c0bus_wb[2]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_24_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_20_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c0bus_wb[2]_i_13 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h505F30305F5F3F3F)) 
    \rgf_c0bus_wb[2]_i_14 
       (.I0(a0bus_0[26]),
        .I1(a0bus_0[2]),
        .I2(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I3(a0bus_0[10]),
        .I4(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[2]_i_15 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(a0bus_0[2]),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \rgf_c0bus_wb[2]_i_16 
       (.I0(\rgf/sreg/sr [8]),
        .I1(p_2_in1_in[5]),
        .I2(\rgf/b0bus_out/bbus_o[5]_INST_0_i_6_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[5]_INST_0_i_5_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[5]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[2]_i_17 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[1]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[2]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[2]_i_18 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBB888B8)) 
    \rgf_c0bus_wb[2]_i_19 
       (.I0(\rgf_c0bus_wb[2]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_19_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[2]_i_2 
       (.I0(cbus_i[2]),
        .I1(ccmd[4]),
        .O(\rgf_c0bus_wb[2]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c0bus_wb[2]_i_20 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h00088808)) 
    \rgf_c0bus_wb[2]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c0bus_wb[2]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFFD080D080)) 
    \rgf_c0bus_wb[2]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_31_n_0 ),
        .I4(a0bus_0[1]),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E2FFFFFFFF)) 
    \rgf_c0bus_wb[2]_i_24 
       (.I0(\rgf_c0bus_wb[27]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_32_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_33_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \rgf_c0bus_wb[2]_i_25 
       (.I0(\rgf_c0bus_wb[18]_i_33_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[2]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c0bus_wb[2]_i_27 
       (.I0(\rgf_c0bus_wb[2]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(a0bus_0[31]),
        .I5(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h5C5F)) 
    \rgf_c0bus_wb[2]_i_28 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(a0bus_0[2]),
        .O(\rgf_c0bus_wb[2]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAA45BB45FFFFFFFF)) 
    \rgf_c0bus_wb[2]_i_29 
       (.I0(\rgf_c0bus_wb[2]_i_36_n_0 ),
        .I1(ctl_selb0_0),
        .I2(\fch/ir0 [4]),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(\fch/ir0 [5]),
        .I5(\bbus_o[5]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[2]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [2]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[2]),
        .I4(\rgf_c0bus_wb[2]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c0bus_wb[2]_i_30 
       (.I0(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[2]_i_31 
       (.I0(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_67_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'h8AFF8A00)) 
    \rgf_c0bus_wb[2]_i_32 
       (.I0(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[2]_i_33 
       (.I0(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[2]_i_34 
       (.I0(\rgf_c0bus_wb[28]_i_42_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\remden[31]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5050503F303F3)) 
    \rgf_c0bus_wb[2]_i_35 
       (.I0(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_67_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_38_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAA2AA)) 
    \rgf_c0bus_wb[2]_i_36 
       (.I0(ctl_selb0_0),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [1]),
        .O(\rgf_c0bus_wb[2]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hF5DDF088)) 
    \rgf_c0bus_wb[2]_i_37 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(\alu0/mul_a_i [30]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[2]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hDFD58F80)) 
    \rgf_c0bus_wb[2]_i_38 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[16]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\alu0/mul_a_i [17]),
        .I4(a0bus_0[15]),
        .O(\rgf_c0bus_wb[2]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[2]_i_4 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h55FD000055FD55FD)) 
    \rgf_c0bus_wb[2]_i_5 
       (.I0(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_12_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_13_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[2]_i_6 
       (.I0(bdatr[10]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[2]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[2]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[2]_i_7 
       (.I0(bdatr[2]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[2]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3]_i_11_n_5 ),
        .I2(\alu0/div/rem [2]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [2]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[2]_i_9 
       (.I0(\rgf_c0bus_wb[2]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[30]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[30]),
        .I2(bdatr[30]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_3_n_0 ),
        .O(c0bus[30]));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_10 
       (.I0(\rgf_c0bus_wb[30]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c0bus_wb[30]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_27_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[30]_i_12 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I2(\alu0/mul_a_i [29]),
        .O(\rgf_c0bus_wb[30]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c0bus_wb[30]_i_13 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[30]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_14 
       (.I0(\rgf_c0bus_wb[30]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \rgf_c0bus_wb[30]_i_15 
       (.I0(\rgf_c0bus_wb[30]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_33_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFF11100000)) 
    \rgf_c0bus_wb[30]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\alu0/mul_a_i [30]),
        .I3(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I5(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hEEFFE0FFA0FFA0FF)) 
    \rgf_c0bus_wb[30]_i_17 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[30]_i_35_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I4(\remden[31]_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c0bus_wb[30]_i_18 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_36_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \rgf_c0bus_wb[30]_i_19 
       (.I0(\rgf_c0bus_wb[30]_i_38_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_17_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c0bus_wb[30]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \rgf_c0bus_wb[30]_i_20 
       (.I0(\rgf_c0bus_wb[30]_i_39_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_40_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_20_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[30]_i_21 
       (.I0(a0bus_0[22]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c0bus_wb[30]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[30]),
        .I2(a0bus_0[30]),
        .O(\rgf_c0bus_wb[30]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[30]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I3(a0bus_0[30]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[30]_i_24 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[29]_i_11_n_5 ),
        .O(\rgf_c0bus_wb[30]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \rgf_c0bus_wb[30]_i_25 
       (.I0(\rgf_c0bus_wb[30]_i_43_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_44_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h1010505F1F1F505F)) 
    \rgf_c0bus_wb[30]_i_26 
       (.I0(\rgf_c0bus_wb[30]_i_45_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[30]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_27 
       (.I0(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[30]_i_28 
       (.I0(\rgf_c0bus_wb[30]_i_48_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_51_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[30]_i_29 
       (.I0(\rgf_c0bus_wb[30]_i_52_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_53_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_54_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_55_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[30]_i_3 
       (.I0(\rgf_c0bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_9_n_0 ),
        .I2(niss_dsp_c0[30]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c0bus_wb[30]_i_30 
       (.I0(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_56_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_57_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[30]_i_31 
       (.I0(\rgf_c0bus_wb[30]_i_58_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_59_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[30]_i_32 
       (.I0(\rgf_c0bus_wb[30]_i_60_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_61_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[30]_i_33 
       (.I0(\rgf_c0bus_wb[30]_i_62_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_63_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h0151FEAE)) 
    \rgf_c0bus_wb[30]_i_34 
       (.I0(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[30]_i_35 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_36 
       (.I0(\rgf_c0bus_wb[20]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_56_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[30]_i_37 
       (.I0(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h55FF565655FFFFFF)) 
    \rgf_c0bus_wb[30]_i_38 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(a0bus_0[30]),
        .I4(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[30]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c0bus_wb[30]_i_39 
       (.I0(a0bus_0[6]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I3(b0bus_0[30]),
        .I4(a0bus_0[30]),
        .O(\rgf_c0bus_wb[30]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c0bus_wb[30]_i_4 
       (.I0(\rgf_c0bus_wb[30]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_11_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_12_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[30]_i_40 
       (.I0(a0bus_0[30]),
        .I1(b0bus_0[30]),
        .O(\rgf_c0bus_wb[30]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h2222222222222220)) 
    \rgf_c0bus_wb[30]_i_41 
       (.I0(\rgf_c0bus_wb[30]_i_64_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I2(\bdatw[15]_INST_0_i_11_n_0 ),
        .I3(\rgf/b0bus_out/bdatw[15]_INST_0_i_12_n_0 ),
        .I4(\rgf/b0bus_out/bdatw[15]_INST_0_i_13_n_0 ),
        .I5(p_2_in1_in[15]),
        .O(\rgf_c0bus_wb[30]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[30]_i_42 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_43 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[16]),
        .O(\rgf_c0bus_wb[30]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_44 
       (.I0(a0bus_0[13]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[14]),
        .O(\rgf_c0bus_wb[30]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[30]_i_45 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_46 
       (.I0(a0bus_0[3]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[30]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_47 
       (.I0(a0bus_0[1]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[2]),
        .O(\rgf_c0bus_wb[30]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_48 
       (.I0(a0bus_0[7]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[30]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_49 
       (.I0(a0bus_0[5]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[30]_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c0bus_wb[30]_i_5 
       (.I0(\rgf_c0bus_wb[30]_i_13_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_50 
       (.I0(a0bus_0[11]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[30]_i_50_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_51 
       (.I0(a0bus_0[9]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[30]_i_51_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_52 
       (.I0(a0bus_0[8]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[30]_i_52_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_53 
       (.I0(a0bus_0[10]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[30]_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_54 
       (.I0(a0bus_0[12]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[30]_i_54_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[30]_i_55 
       (.I0(a0bus_0[13]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[14]),
        .O(\rgf_c0bus_wb[30]_i_55_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_56 
       (.I0(a0bus_0[6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[30]_i_56_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[30]_i_57 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[30]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[30]_i_58 
       (.I0(a0bus_0[28]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[27]),
        .O(\rgf_c0bus_wb[30]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[30]_i_59 
       (.I0(a0bus_0[29]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[30]_i_59_n_0 ));
  LUT5 #(
    .INIT(32'h0000FF47)) 
    \rgf_c0bus_wb[30]_i_6 
       (.I0(\rgf_c0bus_wb[30]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\remden[31]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[30]_i_60 
       (.I0(a0bus_0[24]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[23]),
        .O(\rgf_c0bus_wb[30]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h3333333333333353)) 
    \rgf_c0bus_wb[30]_i_61 
       (.I0(a0bus_0[26]),
        .I1(a0bus_0[25]),
        .I2(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I3(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I5(p_2_in1_in[0]),
        .O(\rgf_c0bus_wb[30]_i_61_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c0bus_wb[30]_i_62 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[16]),
        .O(\rgf_c0bus_wb[30]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h3333333333333353)) 
    \rgf_c0bus_wb[30]_i_63 
       (.I0(a0bus_0[18]),
        .I1(a0bus_0[17]),
        .I2(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I3(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I4(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I5(p_2_in1_in[0]),
        .O(\rgf_c0bus_wb[30]_i_63_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[30]_i_64 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[30]_i_65 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [15]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[15]));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c0bus_wb[30]_i_7 
       (.I0(\rgf_c0bus_wb[30]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \rgf_c0bus_wb[30]_i_8 
       (.I0(\rgf_c0bus_wb[30]_i_20_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_21_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_22_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[30]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_24_n_0 ),
        .I2(\alu0/div/rem [30]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo__0 [30]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[30]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[31]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[31]),
        .I2(bdatr[31]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_4_n_0 ),
        .O(c0bus[31]));
  LUT6 #(
    .INIT(64'h11F111F1FFFF11F1)) 
    \rgf_c0bus_wb[31]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I2(\alu0/div/quo__0 [31]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [31]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c0bus_wb[31]_i_11 
       (.I0(\alu0/mul/mul_rslt ),
        .I1(\niss_dsp_a0[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[31]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c0bus_wb[31]_i_12 
       (.I0(a0bus_0[31]),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[31]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c0bus_wb[31]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I1(\alu0/mul_a_i [30]),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[31]_i_14 
       (.I0(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[31]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c0bus_wb[31]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_39_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_40_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_41_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h04F8)) 
    \rgf_c0bus_wb[31]_i_16 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[31]_i_42_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[31]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_43_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[22]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFF8F)) 
    \rgf_c0bus_wb[31]_i_18 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[31]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\remden[31]_i_3_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c0bus_wb[31]_i_2 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [1]),
        .O(\rgf_c0bus_wb[31]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFF4FCF4F)) 
    \rgf_c0bus_wb[31]_i_20 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBBBFFFB)) 
    \rgf_c0bus_wb[31]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_44_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_10_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_45_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[31]_i_22 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[31]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_46_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_48_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_50_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c0bus_wb[31]_i_25 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_51_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_52_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_27 
       (.I0(\rgf_c0bus_wb[31]_i_53_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_54_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEAAAB0002AAA8)) 
    \rgf_c0bus_wb[31]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_55_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_56_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c0bus_wb[31]_i_29 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_49_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'h000E0E0E)) 
    \rgf_c0bus_wb[31]_i_3 
       (.I0(\rgf_c0bus_wb[31]_i_5_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_6_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_7_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c0bus_wb[31]_i_30 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[31]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hAEEA)) 
    \rgf_c0bus_wb[31]_i_31 
       (.I0(\rgf_c0bus_wb[31]_i_57_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I2(b0bus_0[31]),
        .I3(a0bus_0[31]),
        .O(\rgf_c0bus_wb[31]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0F8F8F0F0F0F0)) 
    \rgf_c0bus_wb[31]_i_32 
       (.I0(a0bus_0[31]),
        .I1(b0bus_0[31]),
        .I2(\rgf_c0bus_wb[23]_i_22_n_0 ),
        .I3(b0bus_0[15]),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hFFA8)) 
    \rgf_c0bus_wb[31]_i_33 
       (.I0(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I1(b0bus_0[31]),
        .I2(a0bus_0[31]),
        .I3(\rgf_c0bus_wb[31]_i_60_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[31]_i_34 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c0bus_wb[31]_i_35 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .O(\rgf_c0bus_wb[31]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_36 
       (.I0(\sr[6]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_62_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hEFFFFFFF)) 
    \rgf_c0bus_wb[31]_i_37 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(div_crdy0),
        .O(\rgf_c0bus_wb[31]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \rgf_c0bus_wb[31]_i_38 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(div_crdy0),
        .I4(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[31]_i_39 
       (.I0(\rgf_c0bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_64_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \rgf_c0bus_wb[31]_i_4 
       (.I0(\rgf_c0bus_wb[31]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_10_n_0 ),
        .I2(niss_dsp_c0[31]),
        .I3(\rgf_c0bus_wb[31]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c0bus_wb[31]_i_40 
       (.I0(\rgf_c0bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(a0bus_0[31]),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[31]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_41 
       (.I0(\rgf_c0bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_67_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_68_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_69_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c0bus_wb[31]_i_42 
       (.I0(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c0bus_wb[31]_i_43 
       (.I0(\rgf_c0bus_wb[18]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_70_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_71_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c0bus_wb[31]_i_44 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[23]_i_25_n_0 ),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c0bus_wb[31]_i_45 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_46 
       (.I0(\rgf_c0bus_wb[31]_i_72_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_73_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_74_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_47 
       (.I0(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_33_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_76_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_48 
       (.I0(a0bus_0[25]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[24]),
        .O(\rgf_c0bus_wb[31]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \rgf_c0bus_wb[31]_i_49 
       (.I0(p_2_in1_in[4]),
        .I1(\rgf/b0bus_out/bbus_o[4]_INST_0_i_5_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[4]_INST_0_i_4_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[4]_INST_0_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_78_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[31]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h8888888A8A8A888A)) 
    \rgf_c0bus_wb[31]_i_5 
       (.I0(\rgf_c0bus_wb[31]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_13_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_50 
       (.I0(a0bus_0[27]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[26]),
        .O(\rgf_c0bus_wb[31]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_51 
       (.I0(a0bus_0[29]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[28]),
        .O(\rgf_c0bus_wb[31]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_52 
       (.I0(a0bus_0[31]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[30]),
        .O(\rgf_c0bus_wb[31]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_53 
       (.I0(a0bus_0[17]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[16]),
        .O(\rgf_c0bus_wb[31]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_54 
       (.I0(a0bus_0[19]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[18]),
        .O(\rgf_c0bus_wb[31]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_55 
       (.I0(a0bus_0[21]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[20]),
        .O(\rgf_c0bus_wb[31]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h00000004FFFFFFF7)) 
    \rgf_c0bus_wb[31]_i_56 
       (.I0(a0bus_0[23]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[22]),
        .O(\rgf_c0bus_wb[31]_i_56_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_57 
       (.I0(a0bus_0[7]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_57_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_58 
       (.I0(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_58_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_59 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFF4FFF4)) 
    \rgf_c0bus_wb[31]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[31]_i_60 
       (.I0(a0bus_0[23]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h5555555400000000)) 
    \rgf_c0bus_wb[31]_i_61 
       (.I0(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I1(\bbus_o[7]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/bbus_o[7]_INST_0_i_3_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[7]_INST_0_i_4_n_0 ),
        .I4(p_2_in1_in[7]),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_61_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_c0bus_wb[31]_i_62 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_62_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_63 
       (.I0(a0bus_0[4]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[31]_i_63_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_64 
       (.I0(a0bus_0[2]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[3]),
        .O(\rgf_c0bus_wb[31]_i_64_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_65 
       (.I0(a0bus_0[0]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[1]),
        .O(\rgf_c0bus_wb[31]_i_65_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c0bus_wb[31]_i_66 
       (.I0(a0bus_0[12]),
        .I1(a0bus_0[13]),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_66_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_67 
       (.I0(a0bus_0[10]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[11]),
        .O(\rgf_c0bus_wb[31]_i_67_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_68 
       (.I0(a0bus_0[8]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[9]),
        .O(\rgf_c0bus_wb[31]_i_68_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_69 
       (.I0(a0bus_0[6]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[31]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \rgf_c0bus_wb[31]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_28_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h555555515555555D)) 
    \rgf_c0bus_wb[31]_i_70 
       (.I0(a0bus_0[17]),
        .I1(\bbus_o[0]_INST_0_i_2_n_0 ),
        .I2(\rgf/b0bus_out/rgf_c0bus_wb[31]_i_77_n_0 ),
        .I3(\rgf/b0bus_out/bbus_o[0]_INST_0_i_6_n_0 ),
        .I4(p_2_in1_in[0]),
        .I5(a0bus_0[16]),
        .O(\rgf_c0bus_wb[31]_i_70_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_71 
       (.I0(a0bus_0[14]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[15]),
        .O(\rgf_c0bus_wb[31]_i_71_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_72 
       (.I0(a0bus_0[9]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[8]),
        .O(\rgf_c0bus_wb[31]_i_72_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_73 
       (.I0(a0bus_0[11]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[10]),
        .O(\rgf_c0bus_wb[31]_i_73_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_74 
       (.I0(a0bus_0[13]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[12]),
        .O(\rgf_c0bus_wb[31]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_75 
       (.I0(a0bus_0[15]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[14]),
        .O(\rgf_c0bus_wb[31]_i_75_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[31]_i_76 
       (.I0(a0bus_0[7]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[31]_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h0AF15FF1FFFFFFFF)) 
    \rgf_c0bus_wb[31]_i_78 
       (.I0(ctl_selb0_0),
        .I1(\fch/ir0 [3]),
        .I2(\rgf_c0bus_wb[31]_i_82_n_0 ),
        .I3(\bdatw[31]_INST_0_i_7_n_0 ),
        .I4(\fch/ir0 [4]),
        .I5(\bbus_o[5]_INST_0_i_2_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_78_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[31]_i_79 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [7]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[31]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \rgf_c0bus_wb[31]_i_82 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [2]),
        .O(\rgf_c0bus_wb[31]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[31]_i_9 
       (.I0(\rgf_c0bus_wb[31]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_32_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_33_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[31]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[3]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[3]),
        .I2(\rgf_c0bus_wb[3]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[3]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_5_n_0 ),
        .O(c0bus[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFF45444545)) 
    \rgf_c0bus_wb[3]_i_10 
       (.I0(\rgf_c0bus_wb[3]_i_19_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_20_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0043CC4C3373FF7F)) 
    \rgf_c0bus_wb[3]_i_12 
       (.I0(a0bus_0[27]),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I4(a0bus_0[3]),
        .I5(\rgf_c0bus_wb[3]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[3]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(a0bus_0[3]),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[3]_i_14 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_28_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_22_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[3]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[19]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[3]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[3]_i_16 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_29_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c0bus_wb[3]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_27_n_0 ),
        .I4(a0bus_0[2]),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFD50000)) 
    \rgf_c0bus_wb[3]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[11]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_27_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4070437340704070)) 
    \rgf_c0bus_wb[3]_i_19 
       (.I0(\rgf_c0bus_wb[20]_i_14_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[19]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_22_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[3]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [3]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[3]),
        .I4(\rgf_c0bus_wb[3]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[3]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[3]_i_20 
       (.I0(\rgf_c0bus_wb[28]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[19]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \rgf_c0bus_wb[3]_i_21 
       (.I0(\rgf_c0bus_wb[2]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_10_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[19]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000030FFFFFFDD)) 
    \rgf_c0bus_wb[3]_i_22 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[3]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h0FDD)) 
    \rgf_c0bus_wb[3]_i_27 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(a0bus_0[11]),
        .I2(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \rgf_c0bus_wb[3]_i_28 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[11]_i_34_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000015155550151)) 
    \rgf_c0bus_wb[3]_i_29 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[28]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[3]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c0bus_wb[3]_i_30 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[3]_i_31 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[2]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[3]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[3]_i_4 
       (.I0(bdatr[3]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[3]_i_5 
       (.I0(bdatr[11]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[3]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[3]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[3]_i_11_n_4 ),
        .I2(\alu0/div/rem [3]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [3]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c0bus_wb[3]_i_7 
       (.I0(\rgf_c0bus_wb[3]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[3]_i_8 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[3]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h000000F2)) 
    \rgf_c0bus_wb[3]_i_9 
       (.I0(\rgf_c0bus_wb[3]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_17_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[3]_i_18_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[4]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[4]),
        .I2(\rgf_c0bus_wb[4]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_5_n_0 ),
        .O(c0bus[4]));
  LUT5 #(
    .INIT(32'h5F4F554F)) 
    \rgf_c0bus_wb[4]_i_10 
       (.I0(\rgf_c0bus_wb[4]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_21_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[4]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[4]_i_11 
       (.I0(a0bus_0[28]),
        .I1(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I2(a0bus_0[4]),
        .O(\rgf_c0bus_wb[4]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c0bus_wb[4]_i_12 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(a0bus_0[12]),
        .I3(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I4(a0bus_0[4]),
        .O(\rgf_c0bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC000FFFFC0006C00)) 
    \rgf_c0bus_wb[4]_i_13 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(a0bus_0[4]),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[4]_i_14 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[20]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[4]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[20]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[4]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c0bus_wb[4]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[20]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[4]_i_17 
       (.I0(\rgf_c0bus_wb[20]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFE200E2)) 
    \rgf_c0bus_wb[4]_i_18 
       (.I0(\rgf_c0bus_wb[21]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_23_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c0bus_wb[4]_i_19 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[4]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [4]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[4]),
        .I4(\rgf_c0bus_wb[4]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c0bus_wb[4]_i_20 
       (.I0(\rgf_c0bus_wb[12]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[21]_i_29_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h20F070F0)) 
    \rgf_c0bus_wb[4]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[12]_i_26_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \rgf_c0bus_wb[4]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_30_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[4]_i_23 
       (.I0(\rgf_c0bus_wb[20]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[20]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[28]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[4]_i_24 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[3]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[4]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h008F)) 
    \rgf_c0bus_wb[4]_i_25 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[3]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[4]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[4]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[4]_i_4 
       (.I0(bdatr[12]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[4]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[4]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[4]_i_5 
       (.I0(bdatr[4]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[4]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_12_n_7 ),
        .I2(\alu0/div/rem [4]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [4]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[4]_i_7 
       (.I0(\rgf_c0bus_wb[4]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[4]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[4]_i_8 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c0bus_wb[4]_i_9 
       (.I0(\rgf_c0bus_wb[4]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[4]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[4]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[5]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[5]),
        .I2(\rgf_c0bus_wb[5]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_5_n_0 ),
        .O(c0bus[5]));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c0bus_wb[5]_i_10 
       (.I0(\rgf_c0bus_wb[5]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_20_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_21_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h5F4F554F)) 
    \rgf_c0bus_wb[5]_i_11 
       (.I0(\rgf_c0bus_wb[5]_i_22_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_23_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[5]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[5]_i_12 
       (.I0(a0bus_0[29]),
        .I1(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I2(a0bus_0[5]),
        .O(\rgf_c0bus_wb[5]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c0bus_wb[5]_i_13 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(a0bus_0[13]),
        .I3(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I4(a0bus_0[5]),
        .O(\rgf_c0bus_wb[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h8800FFFF88006A00)) 
    \rgf_c0bus_wb[5]_i_14 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(a0bus_0[5]),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[5]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[5]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h004080C0)) 
    \rgf_c0bus_wb[5]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[21]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h74)) 
    \rgf_c0bus_wb[5]_i_17 
       (.I0(\rgf_c0bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFDFFFCFF)) 
    \rgf_c0bus_wb[5]_i_18 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_27_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[5]_i_19 
       (.I0(\rgf_c0bus_wb[21]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[5]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [5]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[5]),
        .I4(\rgf_c0bus_wb[5]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[5]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h2222222230333000)) 
    \rgf_c0bus_wb[5]_i_20 
       (.I0(\rgf_c0bus_wb[5]_i_26_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c0bus_wb[5]_i_21 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c0bus_wb[5]_i_22 
       (.I0(\rgf_c0bus_wb[13]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_29_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_18_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h20F070F0)) 
    \rgf_c0bus_wb[5]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_28_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_28_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[13]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[5]_i_24 
       (.I0(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_35_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \rgf_c0bus_wb[5]_i_25 
       (.I0(\rgf_c0bus_wb[17]_i_31_n_0 ),
        .I1(\rgf_c0bus_wb[17]_i_32_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_37_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[5]_i_26 
       (.I0(\rgf_c0bus_wb[25]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[21]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[5]_i_27 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[4]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[5]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h008F)) 
    \rgf_c0bus_wb[5]_i_28 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[4]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[5]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c0bus_wb[5]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[5]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[5]_i_4 
       (.I0(bdatr[13]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[5]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[5]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[5]_i_5 
       (.I0(bdatr[5]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[5]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[5]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_12_n_6 ),
        .I2(\alu0/div/rem [5]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [5]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[5]_i_7 
       (.I0(\rgf_c0bus_wb[5]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[5]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \rgf_c0bus_wb[5]_i_8 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h2222222200022202)) 
    \rgf_c0bus_wb[5]_i_9 
       (.I0(\rgf_c0bus_wb[5]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_17_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I4(a0bus_0[31]),
        .I5(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[5]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hF8F8FFF8)) 
    \rgf_c0bus_wb[6]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[6]),
        .I2(\rgf_c0bus_wb[6]_i_2_n_0 ),
        .I3(bdatr[6]),
        .I4(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .O(c0bus[6]));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[6]_i_10 
       (.I0(\rgf_c0bus_wb[6]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_21_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[6]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[6]_i_11 
       (.I0(a0bus_0[30]),
        .I1(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I2(a0bus_0[6]),
        .O(\rgf_c0bus_wb[6]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c0bus_wb[6]_i_12 
       (.I0(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(a0bus_0[6]),
        .I3(a0bus_0[14]),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c0bus_wb[6]_i_13 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(a0bus_0[6]),
        .I3(\bbus_o[6]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[6]_i_14 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_22_n_0 ),
        .I4(\rgf_c0bus_wb[22]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[6]_i_15 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_22_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[22]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[6]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h5030)) 
    \rgf_c0bus_wb[6]_i_17 
       (.I0(\rgf_c0bus_wb[23]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_13_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h2222222230333000)) 
    \rgf_c0bus_wb[6]_i_18 
       (.I0(\rgf_c0bus_wb[6]_i_23_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_41_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_43_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c0bus_wb[6]_i_19 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hEFEEEFEFEFEEEEEE)) 
    \rgf_c0bus_wb[6]_i_2 
       (.I0(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I3(bdatr[6]),
        .I4(\mem/read_cyc [0]),
        .I5(bdatr[14]),
        .O(\rgf_c0bus_wb[6]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[6]_i_20 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_46_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h20F070F0)) 
    \rgf_c0bus_wb[6]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_41_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h74777444)) 
    \rgf_c0bus_wb[6]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_41_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_26_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c0bus_wb[6]_i_23 
       (.I0(\rgf_c0bus_wb[22]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[6]_i_24 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[5]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[6]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h008F)) 
    \rgf_c0bus_wb[6]_i_25 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[5]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[6]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c0bus_wb[6]_i_26 
       (.I0(\alu0/mul_a_i [20]),
        .I1(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I2(\alu0/mul_a_i [21]),
        .I3(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[18]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[6]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [6]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[6]),
        .I4(\rgf_c0bus_wb[6]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[6]_i_4 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c0bus_wb[6]_i_5 
       (.I0(\mem/read_cyc [3]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .O(\rgf_c0bus_wb[6]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[6]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_12_n_5 ),
        .I2(\alu0/div/rem [6]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [6]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[6]_i_7 
       (.I0(\rgf_c0bus_wb[6]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_13_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[6]_i_8 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c0bus_wb[6]_i_9 
       (.I0(\rgf_c0bus_wb[6]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[6]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_18_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \rgf_c0bus_wb[7]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[7]),
        .I2(\rgf_c0bus_wb[7]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_5_n_0 ),
        .O(c0bus[7]));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c0bus_wb[7]_i_10 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c0bus_wb[7]_i_26_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h5F4F554F)) 
    \rgf_c0bus_wb[7]_i_11 
       (.I0(\rgf_c0bus_wb[7]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_29_n_0 ),
        .I3(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[7]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c0bus_wb[7]_i_13 
       (.I0(a0bus_0[31]),
        .I1(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I2(a0bus_0[7]),
        .O(\rgf_c0bus_wb[7]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[7]_i_14 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \rgf_c0bus_wb[7]_i_15 
       (.I0(b0bus_0[7]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(a0bus_0[15]),
        .I3(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I4(a0bus_0[7]),
        .O(\rgf_c0bus_wb[7]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_16 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \rgf_c0bus_wb[7]_i_17 
       (.I0(\rgf_c0bus_wb[7]_i_35_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(b0bus_0[7]),
        .I3(a0bus_0[7]),
        .I4(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[7]_i_18 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_36_n_0 ),
        .I4(\rgf_c0bus_wb[23]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[7]_i_19 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_36_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[23]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[7]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[7]_i_2 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [7]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[7]),
        .I4(\rgf_c0bus_wb[7]_i_6_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c0bus_wb[7]_i_20 
       (.I0(\rgf_c0bus_wb[23]_i_13_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[7]_i_21 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[7]_i_22 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_23 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c0bus_wb[7]_i_24 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[6]),
        .O(\rgf_c0bus_wb[7]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \rgf_c0bus_wb[7]_i_25 
       (.I0(\bbus_o[2]_INST_0_i_1_n_0 ),
        .I1(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\bbus_o[3]_INST_0_i_1_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[7]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c0bus_wb[7]_i_27 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[23]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h0050F3500050F050)) 
    \rgf_c0bus_wb[7]_i_28 
       (.I0(\rgf_c0bus_wb[16]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_47_n_0 ),
        .I5(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'h80F0D0F0)) 
    \rgf_c0bus_wb[7]_i_29 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_37_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_38_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[7]_i_3 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_9_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_11_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[7]_i_34 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_34_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \rgf_c0bus_wb[7]_i_35 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[7]_i_36 
       (.I0(\rgf_c0bus_wb[7]_i_37_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \rgf_c0bus_wb[7]_i_37 
       (.I0(\rgf_c0bus_wb[30]_i_44_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_50_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_51_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_48_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c0bus_wb[7]_i_38 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_24_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[7]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_c0bus_wb[7]_i_4 
       (.I0(bdatr[7]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E2000000)) 
    \rgf_c0bus_wb[7]_i_5 
       (.I0(bdatr[15]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[7]),
        .I3(\mem/read_cyc [2]),
        .I4(\mem/read_cyc [1]),
        .I5(\mem/read_cyc [3]),
        .O(\rgf_c0bus_wb[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[7]_i_6 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_12_n_4 ),
        .I2(\alu0/div/rem [7]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [7]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c0bus_wb[7]_i_7 
       (.I0(\rgf_c0bus_wb[7]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_17_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[7]_i_8 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_18_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCFDDCFDDFFFFCFDD)) 
    \rgf_c0bus_wb[7]_i_9 
       (.I0(\rgf_c0bus_wb[7]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[7]_i_21_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_22_n_0 ),
        .I3(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I4(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[23]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[8]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[8]),
        .I2(bdatr[8]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_3_n_0 ),
        .O(c0bus[8]));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[8]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_21_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[8]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[8]_i_11 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[8]_i_12 
       (.I0(\rgf_c0bus_wb[24]_i_19_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \rgf_c0bus_wb[8]_i_13 
       (.I0(\rgf_c0bus_wb[24]_i_22_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_24_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c0bus_wb[8]_i_14 
       (.I0(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[24]_i_17_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_10_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_21_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c0bus_wb[8]_i_15 
       (.I0(\rgf_c0bus_wb[25]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_22_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00002F7F)) 
    \rgf_c0bus_wb[8]_i_16 
       (.I0(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_23_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_24_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hD1FFD133D133D1FF)) 
    \rgf_c0bus_wb[8]_i_17 
       (.I0(a0bus_0[16]),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(a0bus_0[8]),
        .I5(b0bus_0[8]),
        .O(\rgf_c0bus_wb[8]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \rgf_c0bus_wb[8]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I1(a0bus_0[8]),
        .I2(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I4(b0bus_0[8]),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \rgf_c0bus_wb[8]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h74777444)) 
    \rgf_c0bus_wb[8]_i_20 
       (.I0(\rgf_c0bus_wb[25]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[14]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_38_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\rgf_c0bus_wb[16]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[8]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[7]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[8]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hB888B8B8)) 
    \rgf_c0bus_wb[8]_i_22 
       (.I0(\rgf_c0bus_wb[31]_i_75_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_34_n_0 ),
        .I3(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c0bus_wb[8]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c0bus_wb[8]_i_23 
       (.I0(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .I4(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_39_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[8]_i_24 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[7]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[8]_i_25 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[8]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[8]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hEEAAEEEA)) 
    \rgf_c0bus_wb[8]_i_26 
       (.I0(\rgf_c0bus_wb[24]_i_24_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I2(b0bus_0[8]),
        .I3(a0bus_0[8]),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[8]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [8]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[8]),
        .I4(\rgf_c0bus_wb[8]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[8]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_10_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c0bus_wb[8]_i_5 
       (.I0(\rgf_c0bus_wb[8]_i_11_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_12_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_14_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[8]_i_6 
       (.I0(\rgf_c0bus_wb[8]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_11_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[8]_i_16_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[8]_i_7 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_i_20_n_7 ),
        .I2(\alu0/div/quo [8]),
        .I3(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .I4(\alu0/div/rem [8]),
        .I5(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h4FFF4F00)) 
    \rgf_c0bus_wb[8]_i_8 
       (.I0(\rgf_c0bus_wb[8]_i_17_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[8]_i_18_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I4(\rgf_c0bus_wb_reg[8]_i_19_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h4F444F4F4F444444)) 
    \rgf_c0bus_wb[8]_i_9 
       (.I0(\rgf_c0bus_wb[24]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .I2(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[8]_i_20_n_0 ),
        .O(\rgf_c0bus_wb[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \rgf_c0bus_wb[9]_i_1 
       (.I0(ccmd[4]),
        .I1(cbus_i[9]),
        .I2(bdatr[9]),
        .I3(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_3_n_0 ),
        .O(c0bus[9]));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c0bus_wb[9]_i_10 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[25]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c0bus_wb[9]_i_11 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_24_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_15_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\rgf_c0bus_wb[9]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c0bus_wb[9]_i_12 
       (.I0(\rgf_c0bus_wb[25]_i_36_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[26]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h3500)) 
    \rgf_c0bus_wb[9]_i_13 
       (.I0(\rgf_c0bus_wb[25]_i_13_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_19_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c0bus_wb[9]_i_14 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c0bus_wb[9]_i_15 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[8]),
        .I2(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[9]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c0bus_wb[9]_i_16 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[25]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c0bus_wb[9]_i_17 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_15_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c0bus_wb[9]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_28_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c0bus_wb[9]_i_19 
       (.I0(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_26_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_27_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_27_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c0bus_wb[9]_i_2 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_6_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h44C0CC0044C00000)) 
    \rgf_c0bus_wb[9]_i_20 
       (.I0(\bbus_o[1]_INST_0_i_1_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_20_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_28_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I5(a0bus_0[17]),
        .O(\rgf_c0bus_wb[9]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c0bus_wb[9]_i_21 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(b0bus_0[9]),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I4(a0bus_0[9]),
        .O(\rgf_c0bus_wb[9]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c0bus_wb[9]_i_22 
       (.I0(a0bus_0[1]),
        .I1(\rgf_c0bus_wb[30]_i_42_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_59_n_0 ),
        .I3(b0bus_0[9]),
        .I4(a0bus_0[9]),
        .I5(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c0bus_wb[9]_i_23 
       (.I0(\rgf_c0bus_wb[31]_i_61_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(b0bus_0[9]),
        .I3(\niss_dsp_a0[32]_INST_0_i_5_n_0 ),
        .I4(a0bus_0[9]),
        .I5(\rgf_c0bus_wb[7]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \rgf_c0bus_wb[9]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I4(\rgf_c0bus_wb[17]_i_25_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c0bus_wb[9]_i_25 
       (.I0(\rgf_c0bus_wb[18]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_30_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c0bus_wb[9]_i_26 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[18]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[13]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c0bus_wb[9]_i_27 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(a0bus_0[8]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h5556555655555556)) 
    \rgf_c0bus_wb[9]_i_28 
       (.I0(a0bus_0[9]),
        .I1(p_2_in1_in[9]),
        .I2(\rgf/b0bus_out/bdatw[9]_INST_0_i_9_n_0 ),
        .I3(\rgf/b0bus_out/bdatw[9]_INST_0_i_8_n_0 ),
        .I4(\bbus_o[5]_INST_0_i_2_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_31_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \rgf_c0bus_wb[9]_i_29 
       (.I0(\rgf_c0bus_wb[16]_i_37_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c0bus_wb[9]_i_3 
       (.I0(\rgf_c0bus_wb[15]_i_7_n_0 ),
        .I1(\alu0/mul/mulh [9]),
        .I2(\rgf_c0bus_wb[15]_i_8_n_0 ),
        .I3(niss_dsp_c0[9]),
        .I4(\rgf_c0bus_wb[9]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c0bus_wb[9]_i_30 
       (.I0(\bdatw[31]_INST_0_i_6_n_0 ),
        .I1(\fch/eir [9]),
        .I2(\bdatw[31]_INST_0_i_7_n_0 ),
        .O(p_2_in1_in[9]));
  LUT6 #(
    .INIT(64'hA6AAAAAAA6AAFFFF)) 
    \rgf_c0bus_wb[9]_i_31 
       (.I0(\bdatw[31]_INST_0_i_7_n_0 ),
        .I1(\bdatw[11]_INST_0_i_19_n_0 ),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .I4(ctl_selb0_0),
        .I5(\fch/ir0 [8]),
        .O(\rgf_c0bus_wb[9]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c0bus_wb[9]_i_4 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_10_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_11_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c0bus_wb[9]_i_5 
       (.I0(\rgf_c0bus_wb[9]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_13_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c0bus_wb[9]_i_6 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[9]_i_15_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_16_n_0 ),
        .I4(\rgf_c0bus_wb[9]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[13]_i_18_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c0bus_wb[9]_i_7 
       (.I0(\rgf_c0bus_wb[9]_i_18_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_14_n_0 ),
        .I2(\rgf_c0bus_wb[9]_i_12_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_19_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c0bus_wb[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c0bus_wb[9]_i_8 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c0bus_wb_reg[11]_i_20_n_6 ),
        .I2(\alu0/div/rem [9]),
        .I3(\rgf_c0bus_wb[31]_i_38_n_0 ),
        .I4(\alu0/div/quo [9]),
        .I5(\rgf_c0bus_wb[31]_i_37_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c0bus_wb[9]_i_9 
       (.I0(\rgf_c0bus_wb[9]_i_20_n_0 ),
        .I1(\rgf_c0bus_wb[9]_i_21_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_22_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[9]_i_23_n_0 ),
        .O(\rgf_c0bus_wb[9]_i_9_n_0 ));
  MUXF7 \rgf_c0bus_wb_reg[10]_i_19 
       (.I0(\rgf_c0bus_wb[10]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_27_n_0 ),
        .O(\rgf_c0bus_wb_reg[10]_i_19_n_0 ),
        .S(\niss_dsp_a0[32]_INST_0_i_4_n_0 ));
  CARRY4 \rgf_c0bus_wb_reg[11]_i_20 
       (.CI(\rgf_c0bus_wb_reg[7]_i_12_n_0 ),
        .CO({\rgf_c0bus_wb_reg[11]_i_20_n_0 ,\rgf_c0bus_wb_reg[11]_i_20_n_1 ,\rgf_c0bus_wb_reg[11]_i_20_n_2 ,\rgf_c0bus_wb_reg[11]_i_20_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a0bus_0[11:8]),
        .O({\rgf_c0bus_wb_reg[11]_i_20_n_4 ,\rgf_c0bus_wb_reg[11]_i_20_n_5 ,\rgf_c0bus_wb_reg[11]_i_20_n_6 ,\rgf_c0bus_wb_reg[11]_i_20_n_7 }),
        .S({\art/add/rgf_c0bus_wb[11]_i_29_n_0 ,\art/add/rgf_c0bus_wb[11]_i_30_n_0 ,\art/add/rgf_c0bus_wb[11]_i_31_n_0 ,\art/add/rgf_c0bus_wb[11]_i_32_n_0 }));
  MUXF7 \rgf_c0bus_wb_reg[12]_i_23 
       (.I0(\rgf_c0bus_wb[12]_i_28_n_0 ),
        .I1(\rgf_c0bus_wb[12]_i_29_n_0 ),
        .O(\rgf_c0bus_wb_reg[12]_i_23_n_0 ),
        .S(\niss_dsp_a0[32]_INST_0_i_4_n_0 ));
  CARRY4 \rgf_c0bus_wb_reg[15]_i_19 
       (.CI(\rgf_c0bus_wb_reg[11]_i_20_n_0 ),
        .CO({\rgf_c0bus_wb_reg[15]_i_19_n_0 ,\rgf_c0bus_wb_reg[15]_i_19_n_1 ,\rgf_c0bus_wb_reg[15]_i_19_n_2 ,\rgf_c0bus_wb_reg[15]_i_19_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a0bus_0[15:12]),
        .O({\rgf_c0bus_wb_reg[15]_i_19_n_4 ,\rgf_c0bus_wb_reg[15]_i_19_n_5 ,\rgf_c0bus_wb_reg[15]_i_19_n_6 ,\rgf_c0bus_wb_reg[15]_i_19_n_7 }),
        .S({\art/add/rgf_c0bus_wb[15]_i_29_n_0 ,\art/add/rgf_c0bus_wb[15]_i_30_n_0 ,\art/add/rgf_c0bus_wb[15]_i_31_n_0 ,\art/add/rgf_c0bus_wb[15]_i_32_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[19]_i_11 
       (.CI(\rgf_c0bus_wb_reg[15]_i_19_n_0 ),
        .CO({\rgf_c0bus_wb_reg[19]_i_11_n_0 ,\rgf_c0bus_wb_reg[19]_i_11_n_1 ,\rgf_c0bus_wb_reg[19]_i_11_n_2 ,\rgf_c0bus_wb_reg[19]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[19]_i_23_n_0 ,\rgf_c0bus_wb[19]_i_24_n_0 ,\rgf_c0bus_wb[19]_i_25_n_0 ,\rgf_c0bus_wb[19]_i_26_n_0 }),
        .O({\rgf_c0bus_wb_reg[19]_i_11_n_4 ,\rgf_c0bus_wb_reg[19]_i_11_n_5 ,\alu0/art/add/tout [18],\rgf_c0bus_wb_reg[19]_i_11_n_7 }),
        .S({\rgf_c0bus_wb[19]_i_27_n_0 ,\art/add/rgf_c0bus_wb[19]_i_28_n_0 ,\art/add/rgf_c0bus_wb[19]_i_29_n_0 ,\art/add/rgf_c0bus_wb[19]_i_30_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[23]_i_24 
       (.CI(\rgf_c0bus_wb_reg[19]_i_11_n_0 ),
        .CO({\rgf_c0bus_wb_reg[23]_i_24_n_0 ,\rgf_c0bus_wb_reg[23]_i_24_n_1 ,\rgf_c0bus_wb_reg[23]_i_24_n_2 ,\rgf_c0bus_wb_reg[23]_i_24_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[23]_i_32_n_0 ,\rgf_c0bus_wb[23]_i_33_n_0 ,\rgf_c0bus_wb[23]_i_34_n_0 ,\rgf_c0bus_wb[23]_i_35_n_0 }),
        .O({\rgf_c0bus_wb_reg[23]_i_24_n_4 ,\rgf_c0bus_wb_reg[23]_i_24_n_5 ,\rgf_c0bus_wb_reg[23]_i_24_n_6 ,\rgf_c0bus_wb_reg[23]_i_24_n_7 }),
        .S({\rgf_c0bus_wb[23]_i_36_n_0 ,\rgf_c0bus_wb[23]_i_37_n_0 ,\art/add/rgf_c0bus_wb[23]_i_38_n_0 ,\art/add/rgf_c0bus_wb[23]_i_39_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[27]_i_23 
       (.CI(\rgf_c0bus_wb_reg[23]_i_24_n_0 ),
        .CO({\rgf_c0bus_wb_reg[27]_i_23_n_0 ,\rgf_c0bus_wb_reg[27]_i_23_n_1 ,\rgf_c0bus_wb_reg[27]_i_23_n_2 ,\rgf_c0bus_wb_reg[27]_i_23_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[27]_i_36_n_0 ,\rgf_c0bus_wb[27]_i_37_n_0 ,\rgf_c0bus_wb[27]_i_38_n_0 ,\rgf_c0bus_wb[27]_i_39_n_0 }),
        .O({\rgf_c0bus_wb_reg[27]_i_23_n_4 ,\rgf_c0bus_wb_reg[27]_i_23_n_5 ,\rgf_c0bus_wb_reg[27]_i_23_n_6 ,\rgf_c0bus_wb_reg[27]_i_23_n_7 }),
        .S({\art/add/rgf_c0bus_wb[27]_i_40_n_0 ,\art/add/rgf_c0bus_wb[27]_i_41_n_0 ,\rgf_c0bus_wb[27]_i_42_n_0 ,\rgf_c0bus_wb[27]_i_43_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[29]_i_11 
       (.CI(\rgf_c0bus_wb_reg[27]_i_23_n_0 ),
        .CO({\rgf_c0bus_wb_reg[29]_i_11_n_0 ,\rgf_c0bus_wb_reg[29]_i_11_n_1 ,\rgf_c0bus_wb_reg[29]_i_11_n_2 ,\rgf_c0bus_wb_reg[29]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c0bus_wb[29]_i_24_n_0 ,\rgf_c0bus_wb[29]_i_25_n_0 ,\rgf_c0bus_wb[29]_i_26_n_0 ,\rgf_c0bus_wb[29]_i_27_n_0 }),
        .O({\rgf_c0bus_wb_reg[29]_i_11_n_4 ,\rgf_c0bus_wb_reg[29]_i_11_n_5 ,\rgf_c0bus_wb_reg[29]_i_11_n_6 ,\rgf_c0bus_wb_reg[29]_i_11_n_7 }),
        .S({\rgf_c0bus_wb[29]_i_28_n_0 ,\art/add/rgf_c0bus_wb[29]_i_29_n_0 ,\art/add/rgf_c0bus_wb[29]_i_30_n_0 ,\rgf_c0bus_wb[29]_i_31_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[3]_i_11 
       (.CI(\<const0> ),
        .CO({\rgf_c0bus_wb_reg[3]_i_11_n_0 ,\rgf_c0bus_wb_reg[3]_i_11_n_1 ,\rgf_c0bus_wb_reg[3]_i_11_n_2 ,\rgf_c0bus_wb_reg[3]_i_11_n_3 }),
        .CYINIT(\rgf_c0bus_wb[3]_i_22_n_0 ),
        .DI(a0bus_0[3:0]),
        .O({\rgf_c0bus_wb_reg[3]_i_11_n_4 ,\rgf_c0bus_wb_reg[3]_i_11_n_5 ,\rgf_c0bus_wb_reg[3]_i_11_n_6 ,\rgf_c0bus_wb_reg[3]_i_11_n_7 }),
        .S({\art/add/rgf_c0bus_wb[3]_i_23_n_0 ,\art/add/rgf_c0bus_wb[3]_i_24_n_0 ,\art/add/rgf_c0bus_wb[3]_i_25_n_0 ,\art/add/rgf_c0bus_wb[3]_i_26_n_0 }));
  CARRY4 \rgf_c0bus_wb_reg[7]_i_12 
       (.CI(\rgf_c0bus_wb_reg[3]_i_11_n_0 ),
        .CO({\rgf_c0bus_wb_reg[7]_i_12_n_0 ,\rgf_c0bus_wb_reg[7]_i_12_n_1 ,\rgf_c0bus_wb_reg[7]_i_12_n_2 ,\rgf_c0bus_wb_reg[7]_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a0bus_0[7:4]),
        .O({\rgf_c0bus_wb_reg[7]_i_12_n_4 ,\rgf_c0bus_wb_reg[7]_i_12_n_5 ,\rgf_c0bus_wb_reg[7]_i_12_n_6 ,\rgf_c0bus_wb_reg[7]_i_12_n_7 }),
        .S({\art/add/rgf_c0bus_wb[7]_i_30_n_0 ,\art/add/rgf_c0bus_wb[7]_i_31_n_0 ,\art/add/rgf_c0bus_wb[7]_i_32_n_0 ,\art/add/rgf_c0bus_wb[7]_i_33_n_0 }));
  MUXF7 \rgf_c0bus_wb_reg[8]_i_19 
       (.I0(\rgf_c0bus_wb[8]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[8]_i_26_n_0 ),
        .O(\rgf_c0bus_wb_reg[8]_i_19_n_0 ),
        .S(\niss_dsp_a0[32]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[0]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_2_n_0 ),
        .I2(bdatr[0]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_4_n_0 ),
        .O(c1bus[0]));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[0]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[0]_i_11 
       (.I0(\rgf_c1bus_wb[16]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h008DFFFF008D008D)) 
    \rgf_c1bus_wb[0]_i_12 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I3(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000A033)) 
    \rgf_c1bus_wb[0]_i_13 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hE0EEE000EEEEEEEE)) 
    \rgf_c1bus_wb[0]_i_14 
       (.I0(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000B8FFB8)) 
    \rgf_c1bus_wb[0]_i_15 
       (.I0(\rgf_c1bus_wb[16]_i_37_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_21_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[0]_i_16 
       (.I0(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h444FFFFF)) 
    \rgf_c1bus_wb[0]_i_17 
       (.I0(\rgf_c1bus_wb[16]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[0]_i_18 
       (.I0(a1bus_0[24]),
        .I1(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I2(a1bus_0[0]),
        .O(\rgf_c1bus_wb[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[0]_i_19 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[8]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[0]),
        .O(\rgf_c1bus_wb[0]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[0]_i_2 
       (.I0(bdatr[0]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[8]),
        .O(\rgf_c1bus_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hC0AEC0EE00EA00AA)) 
    \rgf_c1bus_wb[0]_i_20 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(acmd1[0]),
        .I5(dctl_sign_f_i_2_n_0),
        .O(\rgf_c1bus_wb[0]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[0]_i_21 
       (.I0(acmd1[3]),
        .I1(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[0]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[0]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [0]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[0]),
        .I4(\rgf_c1bus_wb[0]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF4447)) 
    \rgf_c1bus_wb[0]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[0]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hAABA)) 
    \rgf_c1bus_wb[0]_i_6 
       (.I0(\rgf_c1bus_wb[0]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_14_n_0 ),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[0]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hBBFB)) 
    \rgf_c1bus_wb[0]_i_7 
       (.I0(\rgf_c1bus_wb[0]_i_15_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[0]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[0]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[0]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_7 ),
        .I2(\alu1/div/rem [0]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [0]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[0]_i_9 
       (.I0(\rgf_c1bus_wb[0]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[0]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[0]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[10]_i_1 
       (.I0(\rgf_c1bus_wb[10]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[10]),
        .O(c1bus[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[10]_i_10 
       (.I0(\rgf_c1bus_wb[10]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[10]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[10]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[10]),
        .O(\rgf_c1bus_wb[10]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c1bus_wb[10]_i_12 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(a1bus_0[10]),
        .I4(acmd1[3]),
        .I5(b1bus_0[10]),
        .O(\rgf_c1bus_wb[10]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[10]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[10]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[10]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[10]_i_14 
       (.I0(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[10]_i_15 
       (.I0(\rgf_c1bus_wb[26]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h3500350F35003500)) 
    \rgf_c1bus_wb[10]_i_16 
       (.I0(\rgf_c1bus_wb[10]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[10]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h3120333333333333)) 
    \rgf_c1bus_wb[10]_i_18 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[26]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c1bus_wb[10]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[10]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [10]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[10]),
        .I4(\rgf_c1bus_wb[10]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[10]_i_20 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c1bus_wb[10]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h47FF)) 
    \rgf_c1bus_wb[10]_i_22 
       (.I0(\rgf_c1bus_wb[10]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c1bus_wb[10]_i_23 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[10]),
        .I2(b1bus_0[10]),
        .I3(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I4(acmd1[3]),
        .I5(a1bus_0[18]),
        .O(\rgf_c1bus_wb[10]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hB1FFB1AAB155B100)) 
    \rgf_c1bus_wb[10]_i_24 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h1BBB)) 
    \rgf_c1bus_wb[10]_i_25 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[10]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[10]_i_27 
       (.I0(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[10]_i_28 
       (.I0(acmd1[3]),
        .I1(a1bus_0[9]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[10]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[10]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[10]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFCFC055555555)) 
    \rgf_c1bus_wb[10]_i_30 
       (.I0(\rgf_c1bus_wb[10]_i_31_n_0 ),
        .I1(\mul_a[16]_i_1__0_n_0 ),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul_a_i [17]),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[10]_i_31 
       (.I0(\rgf/a1bus_out/rgf_c1bus_wb[10]_i_32_n_0 ),
        .I1(\rgf/a1bus_out/rgf_c1bus_wb[10]_i_33_n_0 ),
        .I2(\rgf/a1bus_out/badr[14]_INST_0_i_6_n_0 ),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[10]_i_35 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf/sreg/sr [14]),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_14_n_0 ),
        .O(\rgf/a1bus_sr [14]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_37 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [14]),
        .O(\rgf_c1bus_wb[10]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_38 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr06 [14]),
        .O(\rgf_c1bus_wb[10]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_39 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [14]),
        .O(\rgf_c1bus_wb[10]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[10]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_5 ),
        .I2(\alu1/div/rem [10]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [10]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[10]_i_40 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [14]),
        .O(\rgf_c1bus_wb[10]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[10]_i_5 
       (.I0(\rgf_c1bus_wb[10]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[10]_i_12_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[10]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[10]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA00EF00EF00)) 
    \rgf_c1bus_wb[10]_i_7 
       (.I0(\rgf_c1bus_wb[10]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEE00F0)) 
    \rgf_c1bus_wb[10]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_17_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c1bus_wb[10]_i_9 
       (.I0(acmd1[3]),
        .I1(a1bus_0[9]),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[10]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[11]_i_1 
       (.I0(\rgf_c1bus_wb[11]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[11]),
        .O(c1bus[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[11]_i_11 
       (.I0(\rgf_c1bus_wb[11]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[11]_i_12 
       (.I0(acmd1[3]),
        .I1(b1bus_0[11]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[11]),
        .O(\rgf_c1bus_wb[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c1bus_wb[11]_i_13 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(a1bus_0[11]),
        .I4(acmd1[3]),
        .I5(b1bus_0[11]),
        .O(\rgf_c1bus_wb[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[11]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[11]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[11]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[11]_i_15 
       (.I0(\rgf_c1bus_wb[11]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0010F010)) 
    \rgf_c1bus_wb[11]_i_16 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[11]_i_17 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[11]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0B0B0F00)) 
    \rgf_c1bus_wb[11]_i_18 
       (.I0(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[28]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c1bus_wb[11]_i_19 
       (.I0(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[11]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [11]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[11]),
        .I4(\rgf_c1bus_wb[11]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEF0FE)) 
    \rgf_c1bus_wb[11]_i_20 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[11]_i_21 
       (.I0(acmd1[3]),
        .I1(a1bus_0[10]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[11]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h1B001B000000FF00)) 
    \rgf_c1bus_wb[11]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_37_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[11]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h00001B00FF001B00)) 
    \rgf_c1bus_wb[11]_i_24 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[11]_i_25 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[11]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c1bus_wb[11]_i_30 
       (.I0(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[11]),
        .I2(b1bus_0[11]),
        .I3(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I4(acmd1[3]),
        .I5(a1bus_0[19]),
        .O(\rgf_c1bus_wb[11]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hCFC05F5FCFC05050)) 
    \rgf_c1bus_wb[11]_i_31 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_37_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_41_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[11]_i_32 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[11]_i_33 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h303F5050303F5F5F)) 
    \rgf_c1bus_wb[11]_i_34 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(\rgf/sreg/sr [6]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[11]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[11]_i_35 
       (.I0(\rgf_c1bus_wb[15]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[11]_i_36 
       (.I0(acmd1[3]),
        .I1(a1bus_0[10]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[11]_i_37 
       (.I0(\alu1/mul_a_i [17]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [18]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[11]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_4 ),
        .I2(\alu1/div/rem [11]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [11]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[11]_i_5 
       (.I0(\rgf_c1bus_wb[11]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_12_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[11]_i_13_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[11]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c1bus_wb[11]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c1bus_wb[11]_i_7 
       (.I0(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_19_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[11]_i_8 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[11]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_22_n_0 ),
        .I4(\rgf_c1bus_wb[11]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[11]_i_9 
       (.I0(\rgf_c1bus_wb[11]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_25_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[12]_i_1 
       (.I0(\rgf_c1bus_wb[12]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[12]),
        .O(c1bus[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[12]_i_10 
       (.I0(\rgf_c1bus_wb[12]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[12]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[12]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[12]),
        .O(\rgf_c1bus_wb[12]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \rgf_c1bus_wb[12]_i_12 
       (.I0(a1bus_0[4]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(a1bus_0[12]),
        .I4(acmd1[3]),
        .I5(b1bus_0[12]),
        .O(\rgf_c1bus_wb[12]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[12]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[12]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[12]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[12]_i_14 
       (.I0(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[12]_i_15 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[12]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00EF00EF00FF0000)) 
    \rgf_c1bus_wb[12]_i_16 
       (.I0(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[29]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[12]_i_17 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h4700FFFF47004700)) 
    \rgf_c1bus_wb[12]_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[12]_i_19 
       (.I0(acmd1[3]),
        .I1(a1bus_0[11]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[12]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[12]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [12]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[12]),
        .I4(\rgf_c1bus_wb[12]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c1bus_wb[12]_i_20 
       (.I0(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[12]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[12]_i_22 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[12]_i_23 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h55FF3C0055003C00)) 
    \rgf_c1bus_wb[12]_i_24 
       (.I0(\bdatw[12]_INST_0_i_4_n_0 ),
        .I1(a1bus_0[12]),
        .I2(b1bus_0[12]),
        .I3(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I4(acmd1[3]),
        .I5(a1bus_0[20]),
        .O(\rgf_c1bus_wb[12]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hCFC05F5FCFC05050)) 
    \rgf_c1bus_wb[12]_i_25 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE4EEE444)) 
    \rgf_c1bus_wb[12]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[12]_i_27 
       (.I0(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[12]_i_28 
       (.I0(acmd1[3]),
        .I1(a1bus_0[11]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_29 
       (.I0(a1bus_0[15]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[12]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[12]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[12]_i_30 
       (.I0(a1bus_0[0]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[12]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[12]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_7 ),
        .I2(\alu1/div/rem [12]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [12]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[12]_i_5 
       (.I0(\rgf_c1bus_wb[12]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[12]_i_12_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[12]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c1bus_wb[12]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c1bus_wb[12]_i_7 
       (.I0(\rgf_c1bus_wb[12]_i_16_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[12]_i_8 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[12]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[12]_i_9 
       (.I0(\rgf_c1bus_wb[12]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[12]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_23_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[13]_i_1 
       (.I0(\rgf_c1bus_wb[13]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[13]),
        .O(c1bus[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[13]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[13]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[13]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[13]_i_12 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[13]),
        .I4(a1bus_0[13]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[13]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[13]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[13]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[13]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[13]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[13]_i_15 
       (.I0(\rgf_c1bus_wb[13]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[13]_i_16 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[13]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c1bus_wb[13]_i_17 
       (.I0(\rgf_c1bus_wb[29]_i_46_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[30]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c1bus_wb[13]_i_18 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h4F444FFF44444444)) 
    \rgf_c1bus_wb[13]_i_19 
       (.I0(\rgf_c1bus_wb[30]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[13]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [13]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[13]),
        .I4(\rgf_c1bus_wb[13]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[13]_i_20 
       (.I0(acmd1[3]),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[13]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c1bus_wb[13]_i_21 
       (.I0(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[13]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[13]_i_23 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[13]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[13]_i_24 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hA3FFA30FA30FA3FF)) 
    \rgf_c1bus_wb[13]_i_25 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[21]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .I4(a1bus_0[13]),
        .I5(b1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hEEE4)) 
    \rgf_c1bus_wb[13]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[13]_i_27 
       (.I0(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[13]_i_28 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hE4EEE444)) 
    \rgf_c1bus_wb[13]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[13]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[13]_i_30 
       (.I0(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[13]_i_31 
       (.I0(acmd1[3]),
        .I1(a1bus_0[12]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[13]_i_32 
       (.I0(a1bus_0[15]),
        .I1(\alu1/asr0 ),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[14]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[13]),
        .O(\rgf_c1bus_wb[13]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_33 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[15]),
        .O(\rgf_c1bus_wb[13]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_34 
       (.I0(a1bus_0[15]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[13]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[13]_i_35 
       (.I0(a1bus_0[13]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[14]),
        .O(\rgf_c1bus_wb[13]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[13]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_6 ),
        .I2(\alu1/div/quo [13]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\alu1/div/rem [13]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[13]_i_5 
       (.I0(\rgf_c1bus_wb[13]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[13]_i_12_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[13]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hA8AA)) 
    \rgf_c1bus_wb[13]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFF1D)) 
    \rgf_c1bus_wb[13]_i_7 
       (.I0(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[13]_i_8 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[13]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[13]_i_9 
       (.I0(\rgf_c1bus_wb[13]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_24_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[13]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[14]_i_1 
       (.I0(\rgf_c1bus_wb[14]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[14]),
        .O(c1bus[14]));
  LUT6 #(
    .INIT(64'h5FC050C000000000)) 
    \rgf_c1bus_wb[14]_i_10 
       (.I0(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[22]),
        .I2(acmd1[3]),
        .I3(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_25_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[14]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[14]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[14]_i_12 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[14]),
        .I4(a1bus_0[14]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[14]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[14]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[14]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[14]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[14]_i_14 
       (.I0(\rgf_c1bus_wb[16]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[14]_i_15 
       (.I0(\rgf_c1bus_wb[30]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[14]_i_16 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[14]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_45_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \rgf_c1bus_wb[14]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[14]_i_19 
       (.I0(acmd1[3]),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[14]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [14]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[14]),
        .I4(\rgf_c1bus_wb[14]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[14]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[14]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[14]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(acmd1[3]),
        .O(\rgf_c1bus_wb[14]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[14]_i_23 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0000757F)) 
    \rgf_c1bus_wb[14]_i_24 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_c1bus_wb[14]_i_25 
       (.I0(a1bus_0[14]),
        .I1(b1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h8BBB)) 
    \rgf_c1bus_wb[14]_i_26 
       (.I0(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_27 
       (.I0(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[14]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_29 
       (.I0(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[14]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[14]_i_30 
       (.I0(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \rgf_c1bus_wb[14]_i_31 
       (.I0(acmd1[3]),
        .I1(a1bus_0[13]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c1bus_wb[14]_i_32 
       (.I0(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I1(a1bus_0[15]),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(a1bus_0[14]),
        .O(\rgf_c1bus_wb[14]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h55577757)) 
    \rgf_c1bus_wb[14]_i_33 
       (.I0(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\alu1/mul_a_i [17]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\mul_a[16]_i_1__0_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h303F5050303F5F5F)) 
    \rgf_c1bus_wb[14]_i_34 
       (.I0(a1bus_0[0]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[14]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[14]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[14]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_5 ),
        .I2(\alu1/div/quo [14]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\alu1/div/rem [14]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[14]_i_5 
       (.I0(\rgf_c1bus_wb[14]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[14]_i_12_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[14]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[14]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[14]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'hFF27)) 
    \rgf_c1bus_wb[14]_i_7 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h7070707070707077)) 
    \rgf_c1bus_wb[14]_i_8 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[14]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[14]_i_9 
       (.I0(\rgf_c1bus_wb[14]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[14]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_24_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[14]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[15]_i_1 
       (.I0(\rgf_c1bus_wb[15]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[15]),
        .O(c1bus[15]));
  LUT6 #(
    .INIT(64'hFFFFFEFEFF00FEFE)) 
    \rgf_c1bus_wb[15]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_45_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h5544040404040404)) 
    \rgf_c1bus_wb[15]_i_11 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I3(acmd1[3]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[15]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hEAFFEAEAEAEAEAEA)) 
    \rgf_c1bus_wb[15]_i_13 
       (.I0(\rgf_c1bus_wb[31]_i_49_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I2(a1bus_0[15]),
        .I3(acmd1[3]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[15]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[15]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[15]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFB8FFFFFF00)) 
    \rgf_c1bus_wb[15]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0000F707)) 
    \rgf_c1bus_wb[15]_i_16 
       (.I0(\rgf_c1bus_wb[15]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I3(a1bus_0[31]),
        .I4(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_17 
       (.I0(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hF070)) 
    \rgf_c1bus_wb[15]_i_18 
       (.I0(acmd1[3]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[30]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hCCDDCFCFFFDDCFCF)) 
    \rgf_c1bus_wb[15]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_61_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[15]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [15]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[15]),
        .I4(\rgf_c1bus_wb[15]_i_6_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hE200)) 
    \rgf_c1bus_wb[15]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[15]_i_21 
       (.I0(acmd1[3]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[15]_i_22 
       (.I0(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_61_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[15]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_c1bus_wb[15]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .I1(\bdatw[12]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[15]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_24 
       (.I0(b1bus_0[15]),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[15]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFF66F0000066F000)) 
    \rgf_c1bus_wb[15]_i_25 
       (.I0(a1bus_0[15]),
        .I1(b1bus_0[15]),
        .I2(a1bus_0[23]),
        .I3(acmd1[3]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(b1bus_0[7]),
        .O(\rgf_c1bus_wb[15]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[15]_i_26 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[15]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \rgf_c1bus_wb[15]_i_27 
       (.I0(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I1(\alu1/mul_a_i [31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[15]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[15]_i_29 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[15]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_9_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c1bus_wb[15]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[15]_i_30 
       (.I0(\rgf_c1bus_wb[24]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[15]_i_31 
       (.I0(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[15]_i_32 
       (.I0(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[15]_i_33 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[15]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c1bus_wb[15]_i_4 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(acmd1[0]),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \rgf_c1bus_wb[15]_i_5 
       (.I0(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I1(\alu1/mul/mul_rslt ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[15]_i_6 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I2(\alu1/div/quo [15]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\alu1/div/rem [15]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hEFE0EFEFEFE0E0E0)) 
    \rgf_c1bus_wb[15]_i_7 
       (.I0(\rgf_c1bus_wb[15]_i_11_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_12_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[15]_i_13_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[15]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hAAAA8A88)) 
    \rgf_c1bus_wb[15]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hD000FFFFD000D000)) 
    \rgf_c1bus_wb[15]_i_9 
       (.I0(\rgf_c1bus_wb[15]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_17_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I4(\rgf_c1bus_wb[15]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[15]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[15]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[16]_i_1 
       (.I0(\rgf_c1bus_wb[16]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[16]),
        .O(c1bus[16]));
  LUT6 #(
    .INIT(64'h8A88AAAA8A888A88)) 
    \rgf_c1bus_wb[16]_i_10 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000FF1010)) 
    \rgf_c1bus_wb[16]_i_11 
       (.I0(\rgf_c1bus_wb[16]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_24_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[16]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h33220003)) 
    \rgf_c1bus_wb[16]_i_12 
       (.I0(\rgf_c1bus_wb[16]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_26_n_0 ),
        .I3(acmd1[3]),
        .I4(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0700FFFF0F0FFFFF)) 
    \rgf_c1bus_wb[16]_i_13 
       (.I0(acmd1[3]),
        .I1(a1bus_0[15]),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[16]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[16]_i_14 
       (.I0(a1bus_0[8]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[16]),
        .I4(a1bus_0[16]),
        .O(\rgf_c1bus_wb[16]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[16]_i_15 
       (.I0(a1bus_0[16]),
        .I1(b1bus_0[16]),
        .O(\rgf_c1bus_wb[16]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[16]_i_16 
       (.I0(a1bus_0[16]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h5151514040405140)) 
    \rgf_c1bus_wb[16]_i_17 
       (.I0(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\rgf_c1bus_wb[16]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[16]_i_18 
       (.I0(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[16]_i_19 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[16]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8F888)) 
    \rgf_c1bus_wb[16]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[16]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hDDC8DDDDDDC88888)) 
    \rgf_c1bus_wb[16]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[16]_i_21 
       (.I0(\rgf_c1bus_wb[16]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \rgf_c1bus_wb[16]_i_22 
       (.I0(acmd1[3]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[16]_i_23 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[16]_i_24 
       (.I0(\rgf_c1bus_wb[16]_i_35_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[16]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[16]_i_25 
       (.I0(\rgf_c1bus_wb[16]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c1bus_wb[16]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFF47)) 
    \rgf_c1bus_wb[16]_i_27 
       (.I0(\rgf_c1bus_wb[16]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_28 
       (.I0(\rgf_c1bus_wb[16]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_46_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_39_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_29 
       (.I0(\rgf_c1bus_wb[16]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[16]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[16]),
        .I2(\rgf_c1bus_wb[16]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19]_i_10_n_7 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c1bus_wb[16]_i_30 
       (.I0(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[16]_i_31 
       (.I0(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_32 
       (.I0(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000AACCAACC)) 
    \rgf_c1bus_wb[16]_i_33 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[16]_i_34 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[16]_i_35 
       (.I0(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[16]_i_36 
       (.I0(\rgf_c1bus_wb[24]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[16]_i_37 
       (.I0(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_38 
       (.I0(a1bus_0[29]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[30]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_39 
       (.I0(a1bus_0[25]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[26]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[16]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_40 
       (.I0(a1bus_0[21]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[22]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFDAAA8FFFCFFFC)) 
    \rgf_c1bus_wb[16]_i_41 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I2(\rgf/a1bus_out/rgf_c1bus_wb[19]_i_39_n_0 ),
        .I3(\rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ),
        .I4(a1bus_0[16]),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[16]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[16]_i_42 
       (.I0(\alu1/mul_a_i [18]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [19]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[16]_i_43 
       (.I0(a1bus_0[16]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[17]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[16]_i_5 
       (.I0(\rgf_c1bus_wb[16]_i_14_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[16]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c1bus_wb[16]_i_6 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[16]),
        .I2(a1bus_0[16]),
        .O(\rgf_c1bus_wb[16]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[16]_i_7 
       (.I0(a1bus_0[24]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[16]_i_8 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I3(a1bus_0[16]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[16]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[16]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [16]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo [16]),
        .O(\rgf_c1bus_wb[16]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[17]_i_1 
       (.I0(\rgf_c1bus_wb[17]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[17]),
        .O(c1bus[17]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[17]_i_10 
       (.I0(\rgf_c1bus_wb[17]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B800000000)) 
    \rgf_c1bus_wb[17]_i_11 
       (.I0(\rgf_c1bus_wb[17]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_21_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[17]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[17]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_24_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[17]_i_14 
       (.I0(a1bus_0[9]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[17]),
        .I4(a1bus_0[17]),
        .O(\rgf_c1bus_wb[17]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[17]_i_15 
       (.I0(a1bus_0[17]),
        .I1(b1bus_0[17]),
        .O(\rgf_c1bus_wb[17]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[17]_i_16 
       (.I0(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[17]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[17]_i_18 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\mul_a[16]_i_1__0_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[17]_i_19 
       (.I0(\rgf_c1bus_wb[25]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF888F8F8)) 
    \rgf_c1bus_wb[17]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[17]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[17]_i_20 
       (.I0(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[17]_i_21 
       (.I0(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[17]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFABFBFFFFFFFF)) 
    \rgf_c1bus_wb[17]_i_23 
       (.I0(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(a1bus_0[1]),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[17]_i_24 
       (.I0(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[17]_i_25 
       (.I0(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_44_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[17]_i_26 
       (.I0(\alu1/mul_a_i [19]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [20]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[17]_i_27 
       (.I0(a1bus_0[17]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[18]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[17]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[17]),
        .I2(\rgf_c1bus_wb[17]_i_9_n_0 ),
        .I3(\alu1/art/add/tout [18]),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[17]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[17]_i_5 
       (.I0(\rgf_c1bus_wb[17]_i_14_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[17]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[17]_i_6 
       (.I0(a1bus_0[25]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[17]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[17]),
        .I2(a1bus_0[17]),
        .O(\rgf_c1bus_wb[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[17]_i_8 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I3(a1bus_0[17]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[17]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[17]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo [17]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [17]),
        .O(\rgf_c1bus_wb[17]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[18]_i_1 
       (.I0(\rgf_c1bus_wb[18]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[18]),
        .O(c1bus[18]));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[18]_i_10 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [17]),
        .O(\rgf_c1bus_wb[18]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \rgf_c1bus_wb[18]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[18]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c1bus_wb[18]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[18]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[18]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[18]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[18]_i_17 
       (.I0(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[18]_i_18 
       (.I0(\rgf_c1bus_wb[26]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[18]_i_19 
       (.I0(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[18]_i_2 
       (.I0(\rgf_c1bus_wb[18]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(\rgf_c1bus_wb[18]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFAFCFA0C)) 
    \rgf_c1bus_wb[18]_i_20 
       (.I0(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[18]_i_21 
       (.I0(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[18]_i_22 
       (.I0(\rgf_c1bus_wb[18]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[18]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[18]_i_24 
       (.I0(a1bus_0[22]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[23]),
        .O(\rgf_c1bus_wb[18]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[18]_i_25 
       (.I0(a1bus_0[20]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[21]),
        .O(\rgf_c1bus_wb[18]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[18]_i_26 
       (.I0(a1bus_0[18]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[19]),
        .O(\rgf_c1bus_wb[18]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFABFBFFFFABFB)) 
    \rgf_c1bus_wb[18]_i_27 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(a1bus_0[1]),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(a1bus_0[2]),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[18]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[18]_i_28 
       (.I0(\alu1/mul_a_i [20]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [21]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[18]_i_29 
       (.I0(a1bus_0[18]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[19]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[18]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[18]),
        .I2(\rgf_c1bus_wb[18]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19]_i_10_n_5 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[18]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[18]_i_5 
       (.I0(a1bus_0[10]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[18]),
        .I4(a1bus_0[18]),
        .O(\rgf_c1bus_wb[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00BC008C00800080)) 
    \rgf_c1bus_wb[18]_i_6 
       (.I0(b1bus_0[15]),
        .I1(acmd1[3]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[4]),
        .I4(b1bus_0[18]),
        .I5(a1bus_0[18]),
        .O(\rgf_c1bus_wb[18]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h000DDDDD)) 
    \rgf_c1bus_wb[18]_i_7 
       (.I0(a1bus_0[26]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[18]),
        .I3(b1bus_0[18]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[18]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[18]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[18]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[18]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[18]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo [18]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [18]),
        .O(\rgf_c1bus_wb[18]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[19]_i_1 
       (.I0(\rgf_c1bus_wb[19]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[19]),
        .O(c1bus[19]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[19]_i_11 
       (.I0(\rgf_c1bus_wb[19]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[19]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c1bus_wb[19]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[19]_i_14 
       (.I0(\rgf_c1bus_wb[19]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hEEEEE000)) 
    \rgf_c1bus_wb[19]_i_15 
       (.I0(\rgf_c1bus_wb[19]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[19]_i_16 
       (.I0(a1bus_0[11]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[19]),
        .I4(a1bus_0[19]),
        .O(\rgf_c1bus_wb[19]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[19]_i_17 
       (.I0(a1bus_0[19]),
        .I1(b1bus_0[19]),
        .O(\rgf_c1bus_wb[19]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[19]_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[19]),
        .O(\rgf_c1bus_wb[19]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF888F8F8)) 
    \rgf_c1bus_wb[19]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[19]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[19]_i_20 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[18]),
        .O(\rgf_c1bus_wb[19]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[19]_i_21 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[17]),
        .O(\rgf_c1bus_wb[19]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0000FFFEFFFE)) 
    \rgf_c1bus_wb[19]_i_22 
       (.I0(\rgf/a1bus_out/badr[15]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [15]),
        .I2(\rgf/a1bus_out/rgf_c1bus_wb[19]_i_39_n_0 ),
        .I3(\rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ),
        .I4(a1bus_0[16]),
        .I5(\rgf/sreg/sr [8]),
        .O(\alu1/asr0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[19]_i_27 
       (.I0(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[19]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_37_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[19]_i_29 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [18]),
        .O(\rgf_c1bus_wb[19]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[19]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[19]),
        .I2(\rgf_c1bus_wb[19]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19]_i_10_n_4 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[19]_i_30 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[19]_i_31 
       (.I0(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[19]_i_32 
       (.I0(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[19]_i_33 
       (.I0(\rgf_c1bus_wb[23]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_c1bus_wb[19]_i_34 
       (.I0(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[19]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hE12D)) 
    \rgf_c1bus_wb[19]_i_40 
       (.I0(b1bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I3(b1bus_0[16]),
        .O(\alu1/art/add/p_0_in ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[19]_i_41 
       (.I0(a1bus_0[19]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[20]),
        .O(\rgf_c1bus_wb[19]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[19]_i_42 
       (.I0(\alu1/mul_a_i [21]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [22]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[19]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[19]_i_44 
       (.I0(a1bus_0[19]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[20]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[19]_i_45 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [15]),
        .O(\rgf_c1bus_wb[19]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[19]_i_46 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [15]),
        .O(\rgf_c1bus_wb[19]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[19]_i_5 
       (.I0(\rgf_c1bus_wb[19]_i_16_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[19]_i_6 
       (.I0(a1bus_0[27]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[19]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[19]),
        .I2(a1bus_0[19]),
        .O(\rgf_c1bus_wb[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[19]_i_8 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I3(a1bus_0[19]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[19]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[19]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [19]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo [19]),
        .O(\rgf_c1bus_wb[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[1]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_2_n_0 ),
        .I2(bdatr[1]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_4_n_0 ),
        .O(c1bus[1]));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[1]_i_10 
       (.I0(\rgf_c1bus_wb[17]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[1]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[1]_i_12 
       (.I0(\rgf_c1bus_wb[1]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[1]_i_13 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c1bus_wb[1]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_26_n_0 ),
        .I4(a1bus_0[0]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[1]_i_15 
       (.I0(\rgf_c1bus_wb[26]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_25_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_c1bus_wb[1]_i_16 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF44F444F444F4)) 
    \rgf_c1bus_wb[1]_i_17 
       (.I0(\rgf_c1bus_wb[17]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_16_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_c1bus_wb[1]_i_18 
       (.I0(\rgf_c1bus_wb[17]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[1]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[17]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[1]_i_2 
       (.I0(bdatr[1]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[9]),
        .O(\rgf_c1bus_wb[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[1]_i_20 
       (.I0(a1bus_0[25]),
        .I1(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I2(a1bus_0[1]),
        .O(\rgf_c1bus_wb[1]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c1bus_wb[1]_i_21 
       (.I0(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[1]),
        .I3(a1bus_0[9]),
        .I4(dctl_sign_f_i_2_n_0),
        .O(\rgf_c1bus_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[1]_i_22 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(a1bus_0[1]),
        .I3(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB1)) 
    \rgf_c1bus_wb[1]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[1]_i_24 
       (.I0(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[1]_i_25 
       (.I0(acmd1[3]),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[1]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[1]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [1]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[1]),
        .I4(\rgf_c1bus_wb[1]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[1]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[1]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[1]_i_6 
       (.I0(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_15_n_0 ),
        .I3(\bdatw[12]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_16_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h555555FF10FF10FF)) 
    \rgf_c1bus_wb[1]_i_7 
       (.I0(\rgf_c1bus_wb[1]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[1]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[1]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[1]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_6 ),
        .I2(\alu1/div/quo [1]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\alu1/div/rem [1]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[1]_i_9 
       (.I0(\rgf_c1bus_wb[1]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[1]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[1]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[20]_i_1 
       (.I0(\rgf_c1bus_wb[20]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[20]),
        .O(c1bus[20]));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[20]_i_10 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [19]),
        .O(\rgf_c1bus_wb[20]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \rgf_c1bus_wb[20]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[20]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[20]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h88FF808088FF80FF)) 
    \rgf_c1bus_wb[20]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[20]_i_15 
       (.I0(a1bus_0[12]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[20]),
        .I4(a1bus_0[20]),
        .O(\rgf_c1bus_wb[20]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[20]_i_16 
       (.I0(a1bus_0[20]),
        .I1(b1bus_0[20]),
        .O(\rgf_c1bus_wb[20]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[20]_i_17 
       (.I0(\rgf_c1bus_wb[29]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[20]_i_18 
       (.I0(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[20]_i_19 
       (.I0(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF888F8F8)) 
    \rgf_c1bus_wb[20]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[20]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[20]_i_20 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[20]_i_21 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \rgf_c1bus_wb[20]_i_22 
       (.I0(\rgf_c1bus_wb[29]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFB73FBFBFFFFFFFF)) 
    \rgf_c1bus_wb[20]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_25_n_0 ),
        .I4(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[20]_i_24 
       (.I0(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h5555555555555557)) 
    \rgf_c1bus_wb[20]_i_25 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(\rgf/a1bus_out/badr[0]_INST_0_i_6_n_0 ),
        .I2(\rgf/a1bus_b13 [0]),
        .I3(\rgf/a1bus_sr [0]),
        .I4(\rgf/a1bus_b02 [0]),
        .I5(\badr[0]_INST_0_i_3_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[20]_i_26 
       (.I0(\rgf_c1bus_wb[22]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\alu1/mul_a_i [20]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\alu1/mul_a_i [21]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[20]_i_27 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf/sreg/sr [0]),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_14_n_0 ),
        .O(\rgf/a1bus_sr [0]));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[20]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[20]),
        .I2(\rgf_c1bus_wb[20]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23]_i_11_n_7 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[20]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[20]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[20]_i_5 
       (.I0(\rgf_c1bus_wb[20]_i_15_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[20]_i_6 
       (.I0(a1bus_0[28]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \rgf_c1bus_wb[20]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[20]),
        .I2(a1bus_0[20]),
        .O(\rgf_c1bus_wb[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[20]_i_8 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I3(a1bus_0[20]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[20]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[20]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [20]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo [20]),
        .O(\rgf_c1bus_wb[20]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[21]_i_1 
       (.I0(\rgf_c1bus_wb[21]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[21]),
        .O(c1bus[21]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[21]_i_10 
       (.I0(\rgf_c1bus_wb[21]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[21]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEEEFEAAAAAAAA)) 
    \rgf_c1bus_wb[21]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[21]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[21]_i_14 
       (.I0(a1bus_0[13]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[21]),
        .I4(a1bus_0[21]),
        .O(\rgf_c1bus_wb[21]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[21]_i_15 
       (.I0(a1bus_0[21]),
        .I1(b1bus_0[21]),
        .O(\rgf_c1bus_wb[21]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[21]_i_16 
       (.I0(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[21]_i_17 
       (.I0(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[21]_i_18 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [20]),
        .O(\rgf_c1bus_wb[21]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[21]_i_19 
       (.I0(\rgf_c1bus_wb[25]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8F888)) 
    \rgf_c1bus_wb[21]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[21]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[21]_i_20 
       (.I0(\rgf_c1bus_wb[29]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFEAE)) 
    \rgf_c1bus_wb[21]_i_21 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[21]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFDA8FFFF)) 
    \rgf_c1bus_wb[21]_i_23 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[21]_i_24 
       (.I0(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[21]_i_25 
       (.I0(a1bus_0[25]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[26]),
        .O(\rgf_c1bus_wb[21]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[21]_i_26 
       (.I0(a1bus_0[23]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[24]),
        .O(\rgf_c1bus_wb[21]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[21]_i_27 
       (.I0(a1bus_0[21]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[22]),
        .O(\rgf_c1bus_wb[21]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[21]_i_28 
       (.I0(\rgf_c1bus_wb[23]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\alu1/mul_a_i [21]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\alu1/mul_a_i [22]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[21]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[21]),
        .I2(\rgf_c1bus_wb[21]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23]_i_11_n_6 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \rgf_c1bus_wb[21]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[21]_i_5 
       (.I0(\rgf_c1bus_wb[21]_i_14_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c1bus_wb[21]_i_6 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[21]),
        .I2(a1bus_0[21]),
        .O(\rgf_c1bus_wb[21]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[21]_i_7 
       (.I0(a1bus_0[29]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[21]_i_8 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I3(a1bus_0[21]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[21]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[21]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo [21]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [21]),
        .O(\rgf_c1bus_wb[21]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[22]_i_1 
       (.I0(\rgf_c1bus_wb[22]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[22]),
        .O(c1bus[22]));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[22]_i_10 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [21]),
        .O(\rgf_c1bus_wb[22]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \rgf_c1bus_wb[22]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[22]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[22]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[22]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \rgf_c1bus_wb[22]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[22]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[22]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[22]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[22]_i_18 
       (.I0(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_40_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFF00FEFE)) 
    \rgf_c1bus_wb[22]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[22]_i_2 
       (.I0(\rgf_c1bus_wb[22]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(\rgf_c1bus_wb[22]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \rgf_c1bus_wb[22]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[22]_i_21 
       (.I0(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[22]_i_22 
       (.I0(\alu1/mul_a_i [24]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [25]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[22]_i_23 
       (.I0(a1bus_0[22]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[23]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[22]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[22]),
        .I2(\rgf_c1bus_wb[22]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23]_i_11_n_5 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[22]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[22]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[22]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[22]_i_5 
       (.I0(a1bus_0[14]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[22]),
        .I4(a1bus_0[22]),
        .O(\rgf_c1bus_wb[22]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[22]_i_6 
       (.I0(b1bus_0[22]),
        .I1(a1bus_0[22]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[22]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h000DDDDD)) 
    \rgf_c1bus_wb[22]_i_7 
       (.I0(a1bus_0[30]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[22]),
        .I3(b1bus_0[22]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[22]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[22]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[22]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[22]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[22]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo [22]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [22]),
        .O(\rgf_c1bus_wb[22]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[23]_i_1 
       (.I0(\rgf_c1bus_wb[23]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[23]),
        .O(c1bus[23]));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[23]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo [23]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [23]),
        .O(\rgf_c1bus_wb[23]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0111011101115555)) 
    \rgf_c1bus_wb[23]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hCF88CF8F)) 
    \rgf_c1bus_wb[23]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFB8)) 
    \rgf_c1bus_wb[23]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[23]_i_15 
       (.I0(\rgf_c1bus_wb[23]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[23]_i_16 
       (.I0(a1bus_0[15]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[23]),
        .I4(a1bus_0[23]),
        .O(\rgf_c1bus_wb[23]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \rgf_c1bus_wb[23]_i_17 
       (.I0(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I1(acmd1[3]),
        .I2(acmd1[4]),
        .I3(b1bus_0[15]),
        .O(\rgf_c1bus_wb[23]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[23]_i_18 
       (.I0(a1bus_0[23]),
        .I1(b1bus_0[23]),
        .O(\rgf_c1bus_wb[23]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_19 
       (.I0(a1bus_0[23]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8F888)) 
    \rgf_c1bus_wb[23]_i_2 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[23]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_20 
       (.I0(acmd1[3]),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[23]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c1bus_wb[23]_i_21 
       (.I0(acmd1[4]),
        .I1(b1bus_0[7]),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[23]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_22 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[23]),
        .O(\rgf_c1bus_wb[23]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_23 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[22]),
        .O(\rgf_c1bus_wb[23]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_24 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[21]),
        .O(\rgf_c1bus_wb[23]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[23]_i_25 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[20]),
        .O(\rgf_c1bus_wb[23]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h2882)) 
    \rgf_c1bus_wb[23]_i_26 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[23]),
        .I2(b1bus_0[23]),
        .I3(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[23]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[23]),
        .I2(\rgf_c1bus_wb[23]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb_reg[23]_i_11_n_4 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[23]_i_30 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \rgf_c1bus_wb[23]_i_31 
       (.I0(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[23]_i_32 
       (.I0(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \rgf_c1bus_wb[23]_i_33 
       (.I0(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[23]_i_34 
       (.I0(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_41_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\alu1/mul_a_i [31]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[23]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_58_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[23]_i_36 
       (.I0(\rgf_c1bus_wb[23]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[23]_i_37 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [22]),
        .O(\rgf_c1bus_wb[23]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[23]_i_38 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[23]_i_39 
       (.I0(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[23]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_14_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[23]_i_40 
       (.I0(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[23]_i_41 
       (.I0(\alu1/mul_a_i [25]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [26]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[23]_i_42 
       (.I0(a1bus_0[23]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[24]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8B8BBB8)) 
    \rgf_c1bus_wb[23]_i_5 
       (.I0(\rgf_c1bus_wb[23]_i_16_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_18_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_6 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(acmd1[0]),
        .O(\rgf_c1bus_wb[23]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \rgf_c1bus_wb[23]_i_7 
       (.I0(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I1(b1bus_0[23]),
        .I2(a1bus_0[23]),
        .O(\rgf_c1bus_wb[23]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[23]_i_8 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \rgf_c1bus_wb[23]_i_9 
       (.I0(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I3(a1bus_0[23]),
        .I4(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[23]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[24]_i_1 
       (.I0(\rgf_c1bus_wb_reg[24]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[24]),
        .O(c1bus[24]));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[24]_i_10 
       (.I0(\rgf_c1bus_wb[24]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \rgf_c1bus_wb[24]_i_11 
       (.I0(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[24]_i_12 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[24]_i_13 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[24]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[24]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c1bus_wb[24]_i_14 
       (.I0(a1bus_0[24]),
        .I1(b1bus_0[24]),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[24]_i_15 
       (.I0(b1bus_0[24]),
        .I1(a1bus_0[24]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[24]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[24]_i_16 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[24]),
        .I4(a1bus_0[24]),
        .O(\rgf_c1bus_wb[24]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAACCAACCF0FFF000)) 
    \rgf_c1bus_wb[24]_i_17 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[24]_i_18 
       (.I0(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hF8F0)) 
    \rgf_c1bus_wb[24]_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[23]),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[24]_i_20 
       (.I0(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[24]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[24]_i_22 
       (.I0(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\alu1/mul_a_i [31]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[24]_i_23 
       (.I0(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000BBBBBBBB)) 
    \rgf_c1bus_wb[24]_i_24 
       (.I0(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[24]_i_25 
       (.I0(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[24]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_72_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[24]_i_27 
       (.I0(\rgf_c1bus_wb[30]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[24]_i_28 
       (.I0(\alu1/mul_a_i [26]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [27]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[24]_i_29 
       (.I0(a1bus_0[31]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[24]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[24]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[24]),
        .I2(\rgf_c1bus_wb[24]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27]_i_10_n_7 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[24]_i_30 
       (.I0(a1bus_0[29]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[28]),
        .O(\rgf_c1bus_wb[24]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[24]_i_31 
       (.I0(a1bus_0[26]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[27]),
        .O(\rgf_c1bus_wb[24]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[24]_i_32 
       (.I0(a1bus_0[25]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[24]),
        .O(\rgf_c1bus_wb[24]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c1bus_wb[24]_i_33 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[24]_i_34 
       (.I0(a1bus_0[24]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[25]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[24]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[24]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [24]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo [24]),
        .O(\rgf_c1bus_wb[24]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[24]_i_8 
       (.I0(\rgf_c1bus_wb[24]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[24]_i_9 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[24]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[25]_i_1 
       (.I0(\rgf_c1bus_wb[25]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[25]),
        .O(c1bus[25]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[25]_i_10 
       (.I0(\rgf_c1bus_wb[25]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[25]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[25]_i_12 
       (.I0(\rgf_c1bus_wb[25]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFE0E0E0)) 
    \rgf_c1bus_wb[25]_i_13 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[25]_i_14 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[25]_i_15 
       (.I0(a1bus_0[17]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[25]_i_16 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[25]_i_17 
       (.I0(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[25]_i_18 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [24]),
        .O(\rgf_c1bus_wb[25]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[25]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hAC00AC0FACF0ACFF)) 
    \rgf_c1bus_wb[25]_i_2 
       (.I0(\rgf_c1bus_wb[25]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_6_n_0 ),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(acmd1[0]),
        .I4(\rgf_c1bus_wb[25]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[25]_i_20 
       (.I0(\rgf_c1bus_wb[25]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[25]_i_21 
       (.I0(\rgf_c1bus_wb[29]_i_44_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\alu1/mul_a_i [31]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \rgf_c1bus_wb[25]_i_22 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFCFAFCFAFCFAFC0)) 
    \rgf_c1bus_wb[25]_i_23 
       (.I0(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[25]_i_24 
       (.I0(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_70_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[25]_i_25 
       (.I0(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[25]_i_26 
       (.I0(\rgf_c1bus_wb[30]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h303F5050303F5F5F)) 
    \rgf_c1bus_wb[25]_i_27 
       (.I0(a1bus_0[31]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[1]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[0]),
        .O(\rgf_c1bus_wb[25]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[25]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_76_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_77_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_71_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[25]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_46_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\alu1/mul_a_i [25]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\alu1/mul_a_i [26]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[25]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[25]),
        .I2(\rgf_c1bus_wb[25]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27]_i_10_n_6 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[25]_i_30 
       (.I0(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[25]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[25]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[25]_i_5 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[25]),
        .I4(a1bus_0[25]),
        .O(\rgf_c1bus_wb[25]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[25]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[25]),
        .I4(a1bus_0[25]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[25]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[25]_i_7 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[25]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[25]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0155)) 
    \rgf_c1bus_wb[25]_i_8 
       (.I0(\rgf_c1bus_wb[25]_i_15_n_0 ),
        .I1(a1bus_0[25]),
        .I2(b1bus_0[25]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[25]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[25]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [25]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo [25]),
        .O(\rgf_c1bus_wb[25]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[26]_i_1 
       (.I0(\rgf_c1bus_wb_reg[26]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[26]),
        .O(c1bus[26]));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[26]_i_10 
       (.I0(\rgf_c1bus_wb[26]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \rgf_c1bus_wb[26]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[26]_i_12 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[26]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[26]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFF22222)) 
    \rgf_c1bus_wb[26]_i_13 
       (.I0(a1bus_0[18]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[26]),
        .I3(b1bus_0[26]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[26]_i_14 
       (.I0(b1bus_0[26]),
        .I1(a1bus_0[26]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[26]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[26]_i_15 
       (.I0(a1bus_0[2]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[26]),
        .I4(a1bus_0[26]),
        .O(\rgf_c1bus_wb[26]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[26]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[26]_i_17 
       (.I0(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[26]_i_18 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [25]),
        .O(\rgf_c1bus_wb[26]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[26]_i_19 
       (.I0(\rgf_c1bus_wb[26]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_20 
       (.I0(\rgf_c1bus_wb[26]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_21 
       (.I0(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4FFE4FFE400)) 
    \rgf_c1bus_wb[26]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\alu1/mul_a_i [31]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hAFCFAFC0)) 
    \rgf_c1bus_wb[26]_i_23 
       (.I0(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCCCCCC480CCCC)) 
    \rgf_c1bus_wb[26]_i_24 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c1bus_wb[26]_i_25 
       (.I0(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_46_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[21]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_26 
       (.I0(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[26]_i_27 
       (.I0(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_50_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[26]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_74_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[26]_i_29 
       (.I0(\rgf_c1bus_wb[26]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\alu1/mul_a_i [26]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\alu1/mul_a_i [27]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[26]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[26]),
        .I2(\rgf_c1bus_wb[26]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27]_i_10_n_5 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFEF40)) 
    \rgf_c1bus_wb[26]_i_30 
       (.I0(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I1(\alu1/mul_a_i [30]),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(\alu1/mul_a_i [31]),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[26]_i_31 
       (.I0(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[26]_i_32 
       (.I0(a1bus_0[28]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[29]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[26]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_8_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[26]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[26]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [26]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo [26]),
        .O(\rgf_c1bus_wb[26]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[26]_i_8 
       (.I0(\rgf_c1bus_wb[26]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[26]_i_9 
       (.I0(\rgf_c1bus_wb[26]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_21_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[26]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[27]_i_1 
       (.I0(\rgf_c1bus_wb[27]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[27]),
        .O(c1bus[27]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[27]_i_11 
       (.I0(\rgf_c1bus_wb[27]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[27]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[27]_i_13 
       (.I0(\rgf_c1bus_wb[27]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \rgf_c1bus_wb[27]_i_14 
       (.I0(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFF0FEFEF0F0F0F0)) 
    \rgf_c1bus_wb[27]_i_15 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[27]_i_16 
       (.I0(a1bus_0[19]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_17 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[27]),
        .O(\rgf_c1bus_wb[27]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_18 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[26]),
        .O(\rgf_c1bus_wb[27]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[25]),
        .O(\rgf_c1bus_wb[27]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[27]_i_2 
       (.I0(\rgf_c1bus_wb[27]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(\rgf_c1bus_wb[27]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_20 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[24]),
        .O(\rgf_c1bus_wb[27]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[27]_i_25 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \rgf_c1bus_wb[27]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_37_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[27]_i_27 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [26]),
        .O(\rgf_c1bus_wb[27]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[27]_i_28 
       (.I0(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[27]_i_29 
       (.I0(\rgf_c1bus_wb[27]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[27]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[27]),
        .I2(\rgf_c1bus_wb[27]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[27]_i_10_n_4 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFEF40)) 
    \rgf_c1bus_wb[27]_i_30 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\alu1/mul_a_i [31]),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBFB0BFBFBFB0B0B0)) 
    \rgf_c1bus_wb[27]_i_31 
       (.I0(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I1(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[27]_i_32 
       (.I0(acmd1[0]),
        .I1(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c1bus_wb[27]_i_33 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I3(\bdatw[12]_INST_0_i_4_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[27]_i_34 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[0]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[3]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[2]),
        .O(\rgf_c1bus_wb[27]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF08080F)) 
    \rgf_c1bus_wb[27]_i_35 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_45_n_0 ),
        .I3(acmd1[0]),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[27]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_36 
       (.I0(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_37 
       (.I0(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_38 
       (.I0(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[27]_i_39 
       (.I0(\rgf_c1bus_wb[31]_i_77_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_71_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_72_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \rgf_c1bus_wb[27]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_12_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_13_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_14_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[27]_i_40 
       (.I0(\rgf_c1bus_wb[31]_i_75_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_76_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFB8FFFFFFB80000)) 
    \rgf_c1bus_wb[27]_i_41 
       (.I0(\alu1/mul_a_i [29]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\alu1/mul_a_i [30]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_41_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_c1bus_wb[27]_i_42 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .O(\rgf_c1bus_wb[27]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[27]_i_43 
       (.I0(a1bus_0[29]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[27]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[27]_i_44 
       (.I0(a1bus_0[27]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[28]),
        .O(\rgf_c1bus_wb[27]_i_44_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[27]_i_45 
       (.I0(acmd1[0]),
        .I1(a1bus_0[31]),
        .O(\rgf_c1bus_wb[27]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[27]_i_46 
       (.I0(a1bus_0[27]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[28]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[27]_i_5 
       (.I0(a1bus_0[3]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[27]),
        .I4(a1bus_0[27]),
        .O(\rgf_c1bus_wb[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[27]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[27]),
        .I4(a1bus_0[27]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[27]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0155)) 
    \rgf_c1bus_wb[27]_i_7 
       (.I0(\rgf_c1bus_wb[27]_i_16_n_0 ),
        .I1(a1bus_0[27]),
        .I2(b1bus_0[27]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[27]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[27]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[27]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[27]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[27]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo [27]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [27]),
        .O(\rgf_c1bus_wb[27]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[28]_i_1 
       (.I0(\rgf_c1bus_wb[28]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[28]),
        .O(c1bus[28]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[28]_i_10 
       (.I0(\rgf_c1bus_wb[28]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[28]_i_11 
       (.I0(\rgf_c1bus_wb[28]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[28]_i_12 
       (.I0(\rgf_c1bus_wb[28]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c1bus_wb[28]_i_13 
       (.I0(\rgf_c1bus_wb[28]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_23_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[28]_i_14 
       (.I0(a1bus_0[20]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[28]_i_15 
       (.I0(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[28]_i_16 
       (.I0(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[28]_i_17 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [27]),
        .O(\rgf_c1bus_wb[28]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hE4FFE4AAE455E400)) 
    \rgf_c1bus_wb[28]_i_18 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_32_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[28]_i_19 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[28]_i_2 
       (.I0(\rgf_c1bus_wb[28]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(\rgf_c1bus_wb[28]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[28]_i_20 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFEF40)) 
    \rgf_c1bus_wb[28]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\alu1/mul_a_i [31]),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[28]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFAAAAAAAA)) 
    \rgf_c1bus_wb[28]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_27_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hF011F0DD)) 
    \rgf_c1bus_wb[28]_i_24 
       (.I0(a1bus_0[16]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_46_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(a1bus_0[15]),
        .O(\rgf_c1bus_wb[28]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_25 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[14]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[11]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[12]),
        .O(\rgf_c1bus_wb[28]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h5050303F5F5F303F)) 
    \rgf_c1bus_wb[28]_i_26 
       (.I0(a1bus_0[1]),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[0]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[28]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_27 
       (.I0(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_28 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[10]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[7]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[8]),
        .O(\rgf_c1bus_wb[28]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_29 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[6]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[3]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[4]),
        .O(\rgf_c1bus_wb[28]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[28]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[28]),
        .I2(\rgf_c1bus_wb[28]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_i_11_n_7 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_30 
       (.I0(\rgf_c1bus_wb[30]_i_50_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_31 
       (.I0(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[28]_i_32 
       (.I0(\rgf_c1bus_wb[30]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h03CF444403CF7777)) 
    \rgf_c1bus_wb[28]_i_33 
       (.I0(a1bus_0[16]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[13]),
        .I3(a1bus_0[14]),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(a1bus_0[15]),
        .O(\rgf_c1bus_wb[28]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_34 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[4]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[3]),
        .O(\rgf_c1bus_wb[28]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c1bus_wb[28]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_74_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(a1bus_0[0]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[28]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_36 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[9]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[12]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[11]),
        .O(\rgf_c1bus_wb[28]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[28]_i_37 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[5]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[8]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[7]),
        .O(\rgf_c1bus_wb[28]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBB8BBB888)) 
    \rgf_c1bus_wb[28]_i_38 
       (.I0(\rgf_c1bus_wb[28]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\alu1/mul_a_i [28]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\alu1/mul_a_i [29]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFB800B8FFB8FFB8)) 
    \rgf_c1bus_wb[28]_i_39 
       (.I0(\rgf_c1bus_wb[28]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_25_n_0 ),
        .I5(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[28]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hB8FFB8FFB8FFB800)) 
    \rgf_c1bus_wb[28]_i_40 
       (.I0(a1bus_0[30]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_43_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[28]_i_41 
       (.I0(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_45_n_0 ),
        .I1(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_46_n_0 ),
        .I2(\rgf/a1bus_out/badr[2]_INST_0_i_6_n_0 ),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_47_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_48_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h01000100010001FF)) 
    \rgf_c1bus_wb[28]_i_42 
       (.I0(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_49_n_0 ),
        .I1(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_50_n_0 ),
        .I2(\rgf/a1bus_out/badr[4]_INST_0_i_6_n_0 ),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_51_n_0 ),
        .I5(\rgf/a1bus_out/rgf_c1bus_wb[28]_i_52_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[28]_i_5 
       (.I0(a1bus_0[4]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[28]),
        .I4(a1bus_0[28]),
        .O(\rgf_c1bus_wb[28]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_56 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf/sreg/sr [2]),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_14_n_0 ),
        .O(\rgf/a1bus_sr [2]));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[28]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[28]),
        .I4(a1bus_0[28]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[28]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_61 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf/sreg/sr [1]),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_14_n_0 ),
        .O(\rgf/a1bus_sr [1]));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_63 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf/sreg/sr [4]),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_14_n_0 ),
        .O(\rgf/a1bus_sr [4]));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[28]_i_68 
       (.I0(\badr[31]_INST_0_i_19_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\rgf/sreg/sr [3]),
        .I3(\badr[31]_INST_0_i_18_n_0 ),
        .I4(\badr[15]_INST_0_i_14_n_0 ),
        .O(\rgf/a1bus_sr [3]));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_69 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [15]),
        .O(\rgf_c1bus_wb[28]_i_69_n_0 ));
  LUT4 #(
    .INIT(16'h0155)) 
    \rgf_c1bus_wb[28]_i_7 
       (.I0(\rgf_c1bus_wb[28]_i_14_n_0 ),
        .I1(a1bus_0[28]),
        .I2(b1bus_0[28]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[28]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_70 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr06 [15]),
        .O(\rgf_c1bus_wb[28]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_71 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [15]),
        .O(\rgf_c1bus_wb[28]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_72 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr26 [15]),
        .O(\rgf_c1bus_wb[28]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_73 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [2]),
        .O(\rgf_c1bus_wb[28]_i_73_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_74 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr06 [2]),
        .O(\rgf_c1bus_wb[28]_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_75 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [2]),
        .O(\rgf_c1bus_wb[28]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_76 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [2]),
        .O(\rgf_c1bus_wb[28]_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_77 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [1]),
        .O(\rgf_c1bus_wb[28]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_78 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr06 [1]),
        .O(\rgf_c1bus_wb[28]_i_78_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_79 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [1]),
        .O(\rgf_c1bus_wb[28]_i_79_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[28]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[28]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[28]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_80 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [1]),
        .O(\rgf_c1bus_wb[28]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_81 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [1]),
        .O(\rgf_c1bus_wb[28]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_82 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr26 [1]),
        .O(\rgf_c1bus_wb[28]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_83 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [4]),
        .O(\rgf_c1bus_wb[28]_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_84 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr06 [4]),
        .O(\rgf_c1bus_wb[28]_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_85 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [4]),
        .O(\rgf_c1bus_wb[28]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_86 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [4]),
        .O(\rgf_c1bus_wb[28]_i_86_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_87 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [3]),
        .O(\rgf_c1bus_wb[28]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_88 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr06 [3]),
        .O(\rgf_c1bus_wb[28]_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_89 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [3]),
        .O(\rgf_c1bus_wb[28]_i_89_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[28]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo__0 [28]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [28]),
        .O(\rgf_c1bus_wb[28]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_90 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [3]),
        .O(\rgf_c1bus_wb[28]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_91 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr25 [3]),
        .O(\rgf_c1bus_wb[28]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[28]_i_92 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\badr[15]_INST_0_i_128_n_0 ),
        .I5(\rgf/bank13/gr26 [3]),
        .O(\rgf_c1bus_wb[28]_i_92_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[29]_i_1 
       (.I0(\rgf_c1bus_wb[29]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[29]),
        .O(c1bus[29]));
  LUT5 #(
    .INIT(32'hFFFF0047)) 
    \rgf_c1bus_wb[29]_i_10 
       (.I0(\rgf_c1bus_wb[29]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEEE222E200000000)) 
    \rgf_c1bus_wb[29]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_c1bus_wb[29]_i_12 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(acmd1[3]),
        .I2(acmd1[0]),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[29]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[29]_i_13 
       (.I0(\rgf_c1bus_wb[29]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c1bus_wb[29]_i_14 
       (.I0(\rgf_c1bus_wb[29]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[29]_i_15 
       (.I0(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I1(acmd1[3]),
        .I2(acmd1[4]),
        .O(\rgf_c1bus_wb[29]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[29]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I1(acmd1[3]),
        .O(\rgf_c1bus_wb[29]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[29]_i_17 
       (.I0(a1bus_0[21]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[29]_i_18 
       (.I0(\rgf_c1bus_wb[29]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[29]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA0C0AFC0A0CFAFCF)) 
    \rgf_c1bus_wb[29]_i_2 
       (.I0(\rgf_c1bus_wb[29]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_6_n_0 ),
        .I2(acmd1[0]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(\rgf_c1bus_wb[29]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_8_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[29]_i_20 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [28]),
        .O(\rgf_c1bus_wb[29]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \rgf_c1bus_wb[29]_i_21 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_35_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[29]_i_22 
       (.I0(\rgf_c1bus_wb[29]_i_37_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[29]_i_23 
       (.I0(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hEFEFEF40)) 
    \rgf_c1bus_wb[29]_i_24 
       (.I0(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\alu1/mul_a_i [31]),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[29]_i_25 
       (.I0(\rgf_c1bus_wb[29]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_45_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[29]_i_26 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_46_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[29]_i_27 
       (.I0(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_70_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h505F505F30303F3F)) 
    \rgf_c1bus_wb[29]_i_28 
       (.I0(a1bus_0[14]),
        .I1(a1bus_0[15]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[12]),
        .I4(a1bus_0[13]),
        .I5(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[29]_i_29 
       (.I0(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[29]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[29]),
        .I2(\rgf_c1bus_wb[29]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_i_11_n_6 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_30 
       (.I0(a1bus_0[2]),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[0]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[1]),
        .O(\rgf_c1bus_wb[29]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hD0FFD000)) 
    \rgf_c1bus_wb[29]_i_31 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_32 
       (.I0(a1bus_0[6]),
        .I1(a1bus_0[7]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[4]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[5]),
        .O(\rgf_c1bus_wb[29]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_33 
       (.I0(a1bus_0[10]),
        .I1(a1bus_0[11]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[8]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[9]),
        .O(\rgf_c1bus_wb[29]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[29]_i_34 
       (.I0(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_71_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_72_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[29]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_76_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_77_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \rgf_c1bus_wb[29]_i_36 
       (.I0(a1bus_0[15]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[14]),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_75_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[29]_i_37 
       (.I0(a1bus_0[31]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[29]_i_37_n_0 ));
  LUT5 #(
    .INIT(32'h0151FEAE)) 
    \rgf_c1bus_wb[29]_i_38 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(\bdatw[12]_INST_0_i_4_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[29]_i_39 
       (.I0(a1bus_0[1]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[0]),
        .O(\rgf_c1bus_wb[29]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \rgf_c1bus_wb[29]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_10_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_13_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_14_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_40 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[5]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[4]),
        .O(\rgf_c1bus_wb[29]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_41 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[6]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[9]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[8]),
        .O(\rgf_c1bus_wb[29]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[29]_i_42 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[10]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[13]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[12]),
        .O(\rgf_c1bus_wb[29]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c1bus_wb[29]_i_43 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I3(\bdatw[12]_INST_0_i_4_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFB8BBB888)) 
    \rgf_c1bus_wb[29]_i_44 
       (.I0(\alu1/mul_a_i [31]),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\alu1/mul_a_i [29]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\alu1/mul_a_i [30]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_c1bus_wb[29]_i_45 
       (.I0(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I1(a1bus_0[0]),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(a1bus_0[1]),
        .O(\rgf_c1bus_wb[29]_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFB8FFFF)) 
    \rgf_c1bus_wb[29]_i_46 
       (.I0(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_43_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[29]_i_5 
       (.I0(a1bus_0[5]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[29]),
        .I4(a1bus_0[29]),
        .O(\rgf_c1bus_wb[29]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0E0A080806020000)) 
    \rgf_c1bus_wb[29]_i_6 
       (.I0(acmd1[3]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(acmd1[4]),
        .I3(b1bus_0[29]),
        .I4(a1bus_0[29]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[29]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h001F)) 
    \rgf_c1bus_wb[29]_i_7 
       (.I0(a1bus_0[29]),
        .I1(b1bus_0[29]),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[29]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \rgf_c1bus_wb[29]_i_8 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[29]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\rgf_c1bus_wb[29]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[29]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [29]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo__0 [29]),
        .O(\rgf_c1bus_wb[29]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[2]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_2_n_0 ),
        .I2(bdatr[2]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_4_n_0 ),
        .O(c1bus[2]));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \rgf_c1bus_wb[2]_i_10 
       (.I0(\rgf_c1bus_wb[10]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[2]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[2]_i_12 
       (.I0(\rgf_c1bus_wb[10]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[2]_i_13 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c1bus_wb[2]_i_14 
       (.I0(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[11]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_29_n_0 ),
        .I4(a1bus_0[1]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hB8B8FF00FFFFFFFF)) 
    \rgf_c1bus_wb[2]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[2]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \rgf_c1bus_wb[2]_i_16 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h04C407C704C404C4)) 
    \rgf_c1bus_wb[2]_i_17 
       (.I0(\rgf_c1bus_wb[18]_i_18_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_31_n_0 ),
        .I4(\rgf_c1bus_wb[18]_i_22_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hCFCAC5C0FFFFFFFF)) 
    \rgf_c1bus_wb[2]_i_18 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[26]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_31_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[2]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_27_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[2]_i_2 
       (.I0(bdatr[2]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[10]),
        .O(\rgf_c1bus_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h505F30305F5F3F3F)) 
    \rgf_c1bus_wb[2]_i_20 
       (.I0(a1bus_0[26]),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I3(a1bus_0[10]),
        .I4(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[2]_i_21 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(a1bus_0[2]),
        .I3(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[2]_i_22 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[26]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[2]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[2]_i_24 
       (.I0(acmd1[3]),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[2]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h5C5F)) 
    \rgf_c1bus_wb[2]_i_25 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(a1bus_0[2]),
        .O(\rgf_c1bus_wb[2]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[2]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[2]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [2]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[2]),
        .I4(\rgf_c1bus_wb[2]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[2]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[2]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[2]_i_6 
       (.I0(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_15_n_0 ),
        .I3(\bdatw[12]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[2]_i_16_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h555555FF10FF10FF)) 
    \rgf_c1bus_wb[2]_i_7 
       (.I0(\rgf_c1bus_wb[2]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[2]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[2]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[2]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_5 ),
        .I2(\alu1/div/rem [2]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [2]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[2]_i_9 
       (.I0(\rgf_c1bus_wb[2]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[30]_i_1 
       (.I0(\rgf_c1bus_wb_reg[30]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[30]),
        .O(c1bus[30]));
  LUT6 #(
    .INIT(64'h0000015155550151)) 
    \rgf_c1bus_wb[30]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAAA)) 
    \rgf_c1bus_wb[30]_i_11 
       (.I0(\rgf_c1bus_wb[29]_i_12_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[30]_i_12 
       (.I0(\rgf_c1bus_wb[30]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \rgf_c1bus_wb[30]_i_13 
       (.I0(\rgf_c1bus_wb[30]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[30]_i_14 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[30]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[30]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFF22222)) 
    \rgf_c1bus_wb[30]_i_15 
       (.I0(a1bus_0[22]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(a1bus_0[30]),
        .I3(b1bus_0[30]),
        .I4(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000FC8000000C80)) 
    \rgf_c1bus_wb[30]_i_16 
       (.I0(b1bus_0[30]),
        .I1(a1bus_0[30]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(b1bus_0[15]),
        .O(\rgf_c1bus_wb[30]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h22F2F222)) 
    \rgf_c1bus_wb[30]_i_17 
       (.I0(a1bus_0[6]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(b1bus_0[30]),
        .I4(a1bus_0[30]),
        .O(\rgf_c1bus_wb[30]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[30]_i_18 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c1bus_wb[30]_i_19 
       (.I0(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_54_n_0 ),
        .I3(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I5(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \rgf_c1bus_wb[30]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_30_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \rgf_c1bus_wb[30]_i_21 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[30]_i_22 
       (.I0(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[30]_i_23 
       (.I0(\rgf_c1bus_wb[30]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_39_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_40_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \rgf_c1bus_wb[30]_i_24 
       (.I0(\rgf_c1bus_wb[30]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\alu1/mul_a_i [31]),
        .I3(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hEEFFE0FFA0FFA0FF)) 
    \rgf_c1bus_wb[30]_i_25 
       (.I0(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[30]_i_42_n_0 ),
        .I3(acmd1[0]),
        .I4(\rgf_c1bus_wb[30]_i_43_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \rgf_c1bus_wb[30]_i_26 
       (.I0(\rgf_c1bus_wb[30]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_44_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFEAA)) 
    \rgf_c1bus_wb[30]_i_27 
       (.I0(\rgf_c1bus_wb[27]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_45_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_28 
       (.I0(a1bus_0[7]),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[5]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[6]),
        .O(\rgf_c1bus_wb[30]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_29 
       (.I0(a1bus_0[11]),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[9]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[10]),
        .O(\rgf_c1bus_wb[30]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \rgf_c1bus_wb[30]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[30]),
        .I2(\rgf_c1bus_wb[30]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb_reg[31]_i_11_n_5 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \rgf_c1bus_wb[30]_i_30 
       (.I0(a1bus_0[0]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [6]),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_31 
       (.I0(a1bus_0[3]),
        .I1(a1bus_0[4]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[1]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[2]),
        .O(\rgf_c1bus_wb[30]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h1D001DCC1D331DFF)) 
    \rgf_c1bus_wb[30]_i_32 
       (.I0(a1bus_0[16]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(a1bus_0[13]),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[30]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[30]_i_33 
       (.I0(\rgf_c1bus_wb[19]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_46_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_34 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[7]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[10]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[9]),
        .O(\rgf_c1bus_wb[30]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h5050303F5F5F303F)) 
    \rgf_c1bus_wb[30]_i_35 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[11]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[13]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[30]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_36 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[6]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[5]),
        .O(\rgf_c1bus_wb[30]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[30]_i_37 
       (.I0(a1bus_0[0]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[2]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[1]),
        .O(\rgf_c1bus_wb[30]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \rgf_c1bus_wb[30]_i_38 
       (.I0(\rgf_c1bus_wb[30]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_49_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_50_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \rgf_c1bus_wb[30]_i_39 
       (.I0(a1bus_0[16]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[15]),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_51_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h00A800A800A8AAAA)) 
    \rgf_c1bus_wb[30]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_11_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[30]_i_40 
       (.I0(\rgf_c1bus_wb[30]_i_52_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_53_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFF1000)) 
    \rgf_c1bus_wb[30]_i_41 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\alu1/mul_a_i [30]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(\alu1/mul_a_i [31]),
        .I5(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_41_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[30]_i_42 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBBBB8)) 
    \rgf_c1bus_wb[30]_i_43 
       (.I0(a1bus_0[31]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf/a1bus_out/badr[15]_INST_0_i_3_n_0 ),
        .I3(\rgf/a1bus_b02 [15]),
        .I4(\rgf/a1bus_out/rgf_c1bus_wb[19]_i_39_n_0 ),
        .I5(\rgf/a1bus_out/badr[15]_INST_0_i_7_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_43_n_0 ));
  LUT5 #(
    .INIT(32'h47CC47FF)) 
    \rgf_c1bus_wb[30]_i_44 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(a1bus_0[2]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(a1bus_0[1]),
        .O(\rgf_c1bus_wb[30]_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_c1bus_wb[30]_i_45 
       (.I0(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_46 
       (.I0(a1bus_0[17]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[18]),
        .O(\rgf_c1bus_wb[30]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_47 
       (.I0(a1bus_0[28]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[27]),
        .O(\rgf_c1bus_wb[30]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[30]_i_48 
       (.I0(a1bus_0[29]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[30]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_49 
       (.I0(a1bus_0[24]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[23]),
        .O(\rgf_c1bus_wb[30]_i_49_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[30]_i_50 
       (.I0(a1bus_0[26]),
        .I1(a1bus_0[25]),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_50_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[30]_i_51 
       (.I0(a1bus_0[18]),
        .I1(a1bus_0[17]),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_51_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_52 
       (.I0(a1bus_0[20]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[19]),
        .O(\rgf_c1bus_wb[30]_i_52_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[30]_i_53 
       (.I0(a1bus_0[22]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[21]),
        .O(\rgf_c1bus_wb[30]_i_53_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[30]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I1(\alu1/div/quo__0 [30]),
        .I2(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I3(\alu1/div/rem [30]),
        .O(\rgf_c1bus_wb[30]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[30]_i_8 
       (.I0(acmd1[4]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .O(\rgf_c1bus_wb[30]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[30]_i_9 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [29]),
        .O(\rgf_c1bus_wb[30]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \rgf_c1bus_wb[31]_i_1 
       (.I0(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(bdatr[31]),
        .O(c1bus[31]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[31]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_c1bus_wb[31]_i_12 
       (.I0(a1bus_0[31]),
        .I1(acmd1[0]),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[31]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \rgf_c1bus_wb[31]_i_13 
       (.I0(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I1(\alu1/mul_a_i [30]),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[31]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \rgf_c1bus_wb[31]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_37_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFF4FFF4)) 
    \rgf_c1bus_wb[31]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_40_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_41_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_44_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_45_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_46_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h00308B00)) 
    \rgf_c1bus_wb[31]_i_17 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[31]),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .O(\rgf_c1bus_wb[31]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFFE0)) 
    \rgf_c1bus_wb[31]_i_18 
       (.I0(a1bus_0[31]),
        .I1(b1bus_0[31]),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hDFC0D5C055005500)) 
    \rgf_c1bus_wb[31]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(b1bus_0[15]),
        .I2(acmd1[3]),
        .I3(a1bus_0[31]),
        .I4(b1bus_0[31]),
        .I5(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'hAEEA)) 
    \rgf_c1bus_wb[31]_i_20 
       (.I0(\rgf_c1bus_wb[31]_i_49_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I2(b1bus_0[31]),
        .I3(a1bus_0[31]),
        .O(\rgf_c1bus_wb[31]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \rgf_c1bus_wb[31]_i_21 
       (.I0(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I1(acmd1[3]),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(div_crdy1),
        .I4(acmd1[4]),
        .I5(acmd1[0]),
        .O(\rgf_c1bus_wb[31]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rgf_c1bus_wb[31]_i_22 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(acmd1[3]),
        .I3(div_crdy1),
        .O(\rgf_c1bus_wb[31]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFDFFFDFFFD)) 
    \rgf_c1bus_wb[31]_i_23 
       (.I0(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I1(acmd1[4]),
        .I2(acmd1[3]),
        .I3(acmd1[0]),
        .I4(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_c1bus_wb[31]_i_24 
       (.I0(acmd1[3]),
        .I1(acmd1[0]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[4]),
        .O(\rgf_c1bus_wb[31]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_25 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[31]),
        .O(\rgf_c1bus_wb[31]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_26 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[30]),
        .O(\rgf_c1bus_wb[31]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_27 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[29]),
        .O(\rgf_c1bus_wb[31]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_28 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[28]),
        .O(\rgf_c1bus_wb[31]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hF4FFF4F4F4F4F4F4)) 
    \rgf_c1bus_wb[31]_i_3 
       (.I0(\rgf_c1bus_wb[31]_i_8_n_0 ),
        .I1(niss_dsp_c1[31]),
        .I2(\rgf_c1bus_wb[31]_i_9_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I4(\rgf_c1bus_wb_reg[31]_i_11_n_4 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[31]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \rgf_c1bus_wb[31]_i_33 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I3(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_34 
       (.I0(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[31]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hAAA9A9A9A9A9A9A9)) 
    \rgf_c1bus_wb[31]_i_36 
       (.I0(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_53_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_54_n_0 ),
        .I3(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I4(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I5(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_36_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_37 
       (.I0(\rgf_c1bus_wb[31]_i_55_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_56_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h04F8)) 
    \rgf_c1bus_wb[31]_i_38 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .I3(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \rgf_c1bus_wb[31]_i_39 
       (.I0(\rgf_c1bus_wb[31]_i_58_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_60_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF8A)) 
    \rgf_c1bus_wb[31]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_14_n_0 ),
        .I3(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_15_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFF8F)) 
    \rgf_c1bus_wb[31]_i_40 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(acmd1[0]),
        .I3(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_40_n_0 ));
  LUT3 #(
    .INIT(8'hAB)) 
    \rgf_c1bus_wb[31]_i_41 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .I2(\alu1/mul_a_i [31]),
        .O(\rgf_c1bus_wb[31]_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFF4FCF4F)) 
    \rgf_c1bus_wb[31]_i_42 
       (.I0(\rgf/sreg/sr [8]),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I3(acmd1[0]),
        .I4(dctl_sign_f_i_2_n_0),
        .O(\rgf_c1bus_wb[31]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h00000000BBBBFFFB)) 
    \rgf_c1bus_wb[31]_i_43 
       (.I0(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[31]_i_61_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_30_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_62_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_c1bus_wb[31]_i_44 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_45 
       (.I0(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_65_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_46 
       (.I0(\rgf_c1bus_wb[31]_i_66_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_67_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[31]_i_47 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_47_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[31]_i_48 
       (.I0(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I1(acmd1[4]),
        .O(\rgf_c1bus_wb[31]_i_48_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[31]_i_49 
       (.I0(a1bus_0[7]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_49_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[31]_i_5 
       (.I0(\mem/read_cyc [2]),
        .I1(\mem/read_cyc [1]),
        .I2(\mem/read_cyc [3]),
        .O(\rgf_c1bus_wb[31]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_50 
       (.I0(a1bus_0[12]),
        .I1(a1bus_0[13]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[10]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[11]),
        .O(\rgf_c1bus_wb[31]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h5555556A6A6A556A)) 
    \rgf_c1bus_wb[31]_i_51 
       (.I0(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I3(\bdatw[12]_INST_0_i_4_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_52 
       (.I0(a1bus_0[8]),
        .I1(a1bus_0[9]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[6]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[7]),
        .O(\rgf_c1bus_wb[31]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \rgf_c1bus_wb[31]_i_53 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf/b1bus_out/rgf_c1bus_wb[31]_i_68_n_0 ),
        .I2(\rgf/b1bus_out/niss_dsp_b1[5]_INST_0_i_5_n_0 ),
        .I3(p_2_in4_in[5]),
        .I4(\niss_dsp_b1[5]_INST_0_i_3_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_2_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \rgf_c1bus_wb[31]_i_54 
       (.I0(p_2_in4_in[4]),
        .I1(\rgf/b1bus_out/bdatw[12]_INST_0_i_15_n_0 ),
        .I2(\rgf/b1bus_b02 [4]),
        .I3(\rgf/b1bus_out/bdatw[12]_INST_0_i_12_n_0 ),
        .I4(\bdatw[12]_INST_0_i_11_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[31]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_55 
       (.I0(a1bus_0[4]),
        .I1(a1bus_0[5]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[2]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[3]),
        .O(\rgf_c1bus_wb[31]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h5F5030305F503F30)) 
    \rgf_c1bus_wb[31]_i_56 
       (.I0(a1bus_0[0]),
        .I1(a1bus_0[1]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[27]_i_42_n_0 ),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[31]_i_56_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_c1bus_wb[31]_i_57 
       (.I0(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I3(\niss_dsp_b1[2]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_57_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[31]_i_58 
       (.I0(\rgf_c1bus_wb[18]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_58_n_0 ));
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \rgf_c1bus_wb[31]_i_59 
       (.I0(\rgf_c1bus_wb[31]_i_70_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I2(a1bus_0[14]),
        .I3(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I4(a1bus_0[15]),
        .O(\rgf_c1bus_wb[31]_i_59_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_60 
       (.I0(\rgf_c1bus_wb[24]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_31_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[24]_i_32_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[18]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_60_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_c1bus_wb[31]_i_61 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[24]_i_33_n_0 ),
        .I2(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_61_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \rgf_c1bus_wb[31]_i_62 
       (.I0(acmd1[0]),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[31]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_63 
       (.I0(a1bus_0[9]),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[11]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[10]),
        .O(\rgf_c1bus_wb[31]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_64 
       (.I0(a1bus_0[13]),
        .I1(a1bus_0[12]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[15]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[14]),
        .O(\rgf_c1bus_wb[31]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h505F3030505F3F3F)) 
    \rgf_c1bus_wb[31]_i_65 
       (.I0(a1bus_0[5]),
        .I1(a1bus_0[4]),
        .I2(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I3(a1bus_0[7]),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(a1bus_0[6]),
        .O(\rgf_c1bus_wb[31]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_66 
       (.I0(\rgf_c1bus_wb[31]_i_71_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_72_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_73_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_74_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[31]_i_67 
       (.I0(\rgf_c1bus_wb[31]_i_75_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_76_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_77_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_78_n_0 ),
        .O(\rgf_c1bus_wb[31]_i_67_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \rgf_c1bus_wb[31]_i_70 
       (.I0(a1bus_0[17]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[16]),
        .O(\rgf_c1bus_wb[31]_i_70_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_71 
       (.I0(a1bus_0[25]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[24]),
        .O(\rgf_c1bus_wb[31]_i_71_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_72 
       (.I0(a1bus_0[27]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[26]),
        .O(\rgf_c1bus_wb[31]_i_72_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_73 
       (.I0(a1bus_0[29]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[28]),
        .O(\rgf_c1bus_wb[31]_i_73_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_74 
       (.I0(a1bus_0[31]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[30]),
        .O(\rgf_c1bus_wb[31]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_75 
       (.I0(a1bus_0[17]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[16]),
        .O(\rgf_c1bus_wb[31]_i_75_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_76 
       (.I0(a1bus_0[19]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[18]),
        .O(\rgf_c1bus_wb[31]_i_76_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_77 
       (.I0(a1bus_0[21]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[20]),
        .O(\rgf_c1bus_wb[31]_i_77_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[31]_i_78 
       (.I0(a1bus_0[23]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[22]),
        .O(\rgf_c1bus_wb[31]_i_78_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_c1bus_wb[31]_i_8 
       (.I0(\alu1/mul/mul_rslt ),
        .I1(\niss_dsp_a1[15]_INST_0_i_1_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_83 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr23 [5]),
        .O(\rgf_c1bus_wb[31]_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_85 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[2]),
        .I3(\niss_dsp_b1[5]_INST_0_i_60_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr21 [5]),
        .O(\rgf_c1bus_wb[31]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \rgf_c1bus_wb[31]_i_87 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr07 [4]),
        .O(\rgf_c1bus_wb[31]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_88 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\rgf/bank_sel [0]),
        .I5(\rgf/bank02/gr05 [4]),
        .O(\rgf_c1bus_wb[31]_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0002000000000000)) 
    \rgf_c1bus_wb[31]_i_89 
       (.I0(ctl_selb1_rn[2]),
        .I1(ctl_selb1_0[2]),
        .I2(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I3(\bdatw[15]_INST_0_i_64_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr27 [4]),
        .O(\rgf_c1bus_wb[31]_i_89_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[31]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I1(\alu1/div/rem [31]),
        .I2(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I3(\alu1/div/quo__0 [31]),
        .O(\rgf_c1bus_wb[31]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_c1bus_wb[31]_i_90 
       (.I0(ctl_selb1_0[2]),
        .I1(\niss_dsp_b1[5]_INST_0_i_58_n_0 ),
        .I2(ctl_selb1_rn[1]),
        .I3(\niss_dsp_b1[2]_INST_0_i_27_n_0 ),
        .I4(\badr[13]_INST_0_i_46_n_0 ),
        .I5(\rgf/bank02/gr25 [4]),
        .O(\rgf_c1bus_wb[31]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[3]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_2_n_0 ),
        .I2(bdatr[3]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_4_n_0 ),
        .O(c1bus[3]));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[3]_i_10 
       (.I0(\rgf_c1bus_wb[19]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[3]_i_11 
       (.I0(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[3]_i_12 
       (.I0(\rgf_c1bus_wb[3]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \rgf_c1bus_wb[3]_i_13 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_18_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hD080FFFFD080D080)) 
    \rgf_c1bus_wb[3]_i_14 
       (.I0(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_35_n_0 ),
        .I4(a1bus_0[2]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hE4E4FF00FFFFFFFF)) 
    \rgf_c1bus_wb[3]_i_15 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[3]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \rgf_c1bus_wb[3]_i_16 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h4070437340704070)) 
    \rgf_c1bus_wb[3]_i_17 
       (.I0(\rgf_c1bus_wb[20]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[19]_i_30_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_34_n_0 ),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hB8FF)) 
    \rgf_c1bus_wb[3]_i_18 
       (.I0(\rgf_c1bus_wb[19]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[27]_i_31_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[3]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[3]_i_2 
       (.I0(bdatr[3]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[11]),
        .O(\rgf_c1bus_wb[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0043CC4C3373FF7F)) 
    \rgf_c1bus_wb[3]_i_21 
       (.I0(a1bus_0[27]),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I4(a1bus_0[3]),
        .I5(\rgf_c1bus_wb[3]_i_31_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[3]_i_22 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(a1bus_0[3]),
        .I3(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB1)) 
    \rgf_c1bus_wb[3]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \rgf_c1bus_wb[3]_i_24 
       (.I0(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[3]_i_25 
       (.I0(acmd1[3]),
        .I1(a1bus_0[2]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[3]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h000000F0FFFFFFDD)) 
    \rgf_c1bus_wb[3]_i_26 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .I5(\rgf/sreg/sr [6]),
        .O(\rgf_c1bus_wb[3]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[3]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_7_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0DDD)) 
    \rgf_c1bus_wb[3]_i_31 
       (.I0(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I1(a1bus_0[11]),
        .I2(\niss_dsp_b1[3]_INST_0_i_1_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[3]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [3]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[3]),
        .I4(\rgf_c1bus_wb[3]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[3]_i_5 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_11_n_0 ),
        .I5(\rgf_c1bus_wb[3]_i_12_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF220F22)) 
    \rgf_c1bus_wb[3]_i_6 
       (.I0(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_15_n_0 ),
        .I3(\bdatw[12]_INST_0_i_4_n_0 ),
        .I4(\rgf_c1bus_wb[3]_i_16_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h555555FF10FF10FF)) 
    \rgf_c1bus_wb[3]_i_7 
       (.I0(\rgf_c1bus_wb[3]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_13_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[3]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[3]_i_8 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[3]_i_20_n_4 ),
        .I2(\alu1/div/rem [3]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [3]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \rgf_c1bus_wb[3]_i_9 
       (.I0(\rgf_c1bus_wb[3]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I2(\rgf_c1bus_wb[3]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[3]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[4]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_2_n_0 ),
        .I2(bdatr[4]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_4_n_0 ),
        .O(c1bus[4]));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[4]_i_10 
       (.I0(\rgf_c1bus_wb[4]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_21_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[4]_i_11 
       (.I0(\rgf_c1bus_wb[20]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h004080C000400040)) 
    \rgf_c1bus_wb[4]_i_12 
       (.I0(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[20]_i_25_n_0 ),
        .I5(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF2E002E)) 
    \rgf_c1bus_wb[4]_i_13 
       (.I0(\rgf_c1bus_wb[4]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(a1bus_0[31]),
        .I5(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_c1bus_wb[4]_i_14 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[4]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[4]_i_15 
       (.I0(\rgf_c1bus_wb[20]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_20_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[4]_i_16 
       (.I0(\rgf_c1bus_wb[21]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_22_n_0 ),
        .I3(acmd1[3]),
        .O(\rgf_c1bus_wb[4]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[4]_i_17 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[20]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[4]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[29]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h222AAA2A)) 
    \rgf_c1bus_wb[4]_i_19 
       (.I0(\rgf_c1bus_wb[4]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_27_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[4]_i_2 
       (.I0(bdatr[4]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[12]),
        .O(\rgf_c1bus_wb[4]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[4]_i_20 
       (.I0(a1bus_0[28]),
        .I1(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I2(a1bus_0[4]),
        .O(\rgf_c1bus_wb[4]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[4]_i_21 
       (.I0(\bdatw[12]_INST_0_i_4_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[12]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[4]),
        .O(\rgf_c1bus_wb[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hC000FFFFC0006C00)) 
    \rgf_c1bus_wb[4]_i_22 
       (.I0(acmd1[0]),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(a1bus_0[4]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB1)) 
    \rgf_c1bus_wb[4]_i_23 
       (.I0(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B8FFFFFFFF)) 
    \rgf_c1bus_wb[4]_i_24 
       (.I0(\rgf_c1bus_wb[4]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_42_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[28]_i_41_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[4]_i_25 
       (.I0(acmd1[3]),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[4]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h008F)) 
    \rgf_c1bus_wb[4]_i_26 
       (.I0(acmd1[3]),
        .I1(a1bus_0[3]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0001FFFFFFFFFFFF)) 
    \rgf_c1bus_wb[4]_i_27 
       (.I0(\badr[0]_INST_0_i_3_n_0 ),
        .I1(\rgf/a1bus_b02 [0]),
        .I2(\rgf/a1bus_out/rgf_c1bus_wb[4]_i_28_n_0 ),
        .I3(\rgf/a1bus_out/badr[0]_INST_0_i_6_n_0 ),
        .I4(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I5(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \rgf_c1bus_wb[4]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[4]_i_30 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_14_n_0 ),
        .I2(\badr[15]_INST_0_i_15_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr05 [0]),
        .O(\rgf_c1bus_wb[4]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \rgf_c1bus_wb[4]_i_31 
       (.I0(\badr[31]_INST_0_i_67_n_0 ),
        .I1(\badr[15]_INST_0_i_15_n_0 ),
        .I2(\badr[15]_INST_0_i_14_n_0 ),
        .I3(\badr[31]_INST_0_i_19_n_0 ),
        .I4(\grn[15]_i_4__7_n_0 ),
        .I5(\rgf/bank13/gr06 [0]),
        .O(\rgf_c1bus_wb[4]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[4]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [4]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[4]),
        .I4(\rgf_c1bus_wb[4]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \rgf_c1bus_wb[4]_i_5 
       (.I0(acmd1[0]),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(acmd1[3]),
        .O(\rgf_c1bus_wb[4]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FF47)) 
    \rgf_c1bus_wb[4]_i_6 
       (.I0(a1bus_0[31]),
        .I1(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_11_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[4]_i_12_n_0 ),
        .I5(\rgf_c1bus_wb[4]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDD00CF00CF00)) 
    \rgf_c1bus_wb[4]_i_7 
       (.I0(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_17_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[4]_i_8 
       (.I0(\rgf_c1bus_wb[4]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[4]_i_16_n_0 ),
        .I3(\rgf_c1bus_wb[4]_i_19_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[4]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_7 ),
        .I2(\alu1/div/rem [4]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [4]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[5]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_2_n_0 ),
        .I2(bdatr[5]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_4_n_0 ),
        .O(c1bus[5]));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[5]_i_10 
       (.I0(\rgf_c1bus_wb[5]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[5]_i_11 
       (.I0(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[21]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[5]_i_12 
       (.I0(\rgf_c1bus_wb[21]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2222222230333000)) 
    \rgf_c1bus_wb[5]_i_13 
       (.I0(\rgf_c1bus_wb[5]_i_26_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[5]_i_14 
       (.I0(\rgf_c1bus_wb[21]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[5]_i_15 
       (.I0(acmd1[3]),
        .I1(a1bus_0[4]),
        .O(\rgf_c1bus_wb[5]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c1bus_wb[5]_i_16 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[5]_i_17 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[5]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[14]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[13]_i_29_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFDFFFCFF)) 
    \rgf_c1bus_wb[5]_i_19 
       (.I0(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_40_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_45_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_2 
       (.I0(bdatr[5]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[13]),
        .O(\rgf_c1bus_wb[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h08AA2AAA)) 
    \rgf_c1bus_wb[5]_i_20 
       (.I0(\rgf_c1bus_wb[5]_i_27_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[5]_i_21 
       (.I0(a1bus_0[29]),
        .I1(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I2(a1bus_0[5]),
        .O(\rgf_c1bus_wb[5]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[5]_i_22 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[13]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[5]),
        .O(\rgf_c1bus_wb[5]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h8800FFFF88006A00)) 
    \rgf_c1bus_wb[5]_i_23 
       (.I0(dctl_sign_f_i_2_n_0),
        .I1(a1bus_0[5]),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h3F305F5F3F305050)) 
    \rgf_c1bus_wb[5]_i_24 
       (.I0(\rgf_c1bus_wb[30]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_25 
       (.I0(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[5]_i_26 
       (.I0(\rgf_c1bus_wb[21]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[5]_i_27 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_15_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[5]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[5]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[5]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[5]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [5]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[5]),
        .I4(\rgf_c1bus_wb[5]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[5]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[5]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hCDCDCDFD)) 
    \rgf_c1bus_wb[5]_i_6 
       (.I0(\rgf_c1bus_wb[5]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_14_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c1bus_wb[5]_i_7 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c1bus_wb[5]_i_16_n_0 ),
        .I5(\rgf_c1bus_wb[5]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[5]_i_8 
       (.I0(\rgf_c1bus_wb[5]_i_18_n_0 ),
        .I1(\rgf_c1bus_wb[5]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[5]_i_20_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[5]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_6 ),
        .I2(\alu1/div/rem [5]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [5]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[6]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I2(bdatr[6]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_4_n_0 ),
        .O(c1bus[6]));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[6]_i_10 
       (.I0(\rgf_c1bus_wb[6]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_22_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[6]_i_11 
       (.I0(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_24_n_0 ),
        .I4(\rgf_c1bus_wb[22]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[6]_i_12 
       (.I0(\rgf_c1bus_wb[22]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2222222230333000)) 
    \rgf_c1bus_wb[6]_i_13 
       (.I0(\rgf_c1bus_wb[22]_i_19_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_25_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \rgf_c1bus_wb[6]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[22]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_c1bus_wb[6]_i_15 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[6]_i_16 
       (.I0(acmd1[3]),
        .I1(a1bus_0[5]),
        .O(\rgf_c1bus_wb[6]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \rgf_c1bus_wb[6]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[6]_i_18 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[22]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c1bus_wb[6]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_63_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_64_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[14]_i_28_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[6]_i_2 
       (.I0(bdatr[6]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[14]),
        .O(\rgf_c1bus_wb[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h08AA2AAA)) 
    \rgf_c1bus_wb[6]_i_20 
       (.I0(\rgf_c1bus_wb[6]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_35_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[14]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[6]_i_21 
       (.I0(a1bus_0[30]),
        .I1(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I2(a1bus_0[6]),
        .O(\rgf_c1bus_wb[6]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8B8)) 
    \rgf_c1bus_wb[6]_i_22 
       (.I0(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[6]),
        .I3(a1bus_0[14]),
        .I4(dctl_sign_f_i_2_n_0),
        .O(\rgf_c1bus_wb[6]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hC0BEC0EE00AA00AA)) 
    \rgf_c1bus_wb[6]_i_23 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(a1bus_0[6]),
        .I3(\niss_dsp_b1[6]_INST_0_i_1_n_0 ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \rgf_c1bus_wb[6]_i_24 
       (.I0(\rgf_c1bus_wb[31]_i_50_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_52_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[18]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[6]_i_25 
       (.I0(\rgf_c1bus_wb[31]_i_58_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_59_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[6]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[6]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[6]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_6_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_7_n_0 ),
        .I4(\rgf_c1bus_wb[6]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[6]_i_4 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [6]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[6]),
        .I4(\rgf_c1bus_wb[6]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[6]_i_5 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_11_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_12_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[6]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hCDFD)) 
    \rgf_c1bus_wb[6]_i_6 
       (.I0(\rgf_c1bus_wb[6]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_14_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c1bus_wb[6]_i_7 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c1bus_wb[6]_i_17_n_0 ),
        .I5(\rgf_c1bus_wb[6]_i_18_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[6]_i_8 
       (.I0(\rgf_c1bus_wb[6]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[6]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_13_n_0 ),
        .I3(\rgf_c1bus_wb[6]_i_20_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[6]_i_9 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_5 ),
        .I2(\alu1/div/rem [6]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [6]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \rgf_c1bus_wb[7]_i_1 
       (.I0(\rgf_c1bus_wb[7]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_3_n_0 ),
        .I2(bdatr[7]),
        .I3(\rgf_c1bus_wb[31]_i_5_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_5_n_0 ),
        .O(c1bus[7]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[7]_i_10 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_4 ),
        .I2(\alu1/div/rem [7]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [7]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \rgf_c1bus_wb[7]_i_11 
       (.I0(\rgf_c1bus_wb[7]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_27_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h00E2)) 
    \rgf_c1bus_wb[7]_i_12 
       (.I0(\rgf_c1bus_wb[7]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(a1bus_0[31]),
        .I3(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[7]_i_13 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_34_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[7]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h2230)) 
    \rgf_c1bus_wb[7]_i_14 
       (.I0(\rgf_c1bus_wb[23]_i_33_n_0 ),
        .I1(acmd1[3]),
        .I2(\rgf_c1bus_wb[24]_i_17_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[7]_i_15 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(acmd1[3]),
        .O(\rgf_c1bus_wb[7]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_c1bus_wb[7]_i_16 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_16_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[7]_i_17 
       (.I0(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_c1bus_wb[7]_i_18 
       (.I0(acmd1[3]),
        .I1(a1bus_0[6]),
        .O(\rgf_c1bus_wb[7]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[7]_i_19 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \rgf_c1bus_wb[7]_i_2 
       (.I0(\mem/read_cyc [1]),
        .I1(\mem/read_cyc [2]),
        .I2(\mem/read_cyc [3]),
        .O(\rgf_c1bus_wb[7]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \rgf_c1bus_wb[7]_i_20 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_36_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00004700FF004700)) 
    \rgf_c1bus_wb[7]_i_21 
       (.I0(\rgf_c1bus_wb[28]_i_36_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[11]_i_34_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hAA2A222A)) 
    \rgf_c1bus_wb[7]_i_22 
       (.I0(\rgf_c1bus_wb[7]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_32_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \rgf_c1bus_wb[7]_i_24 
       (.I0(a1bus_0[31]),
        .I1(\niss_dsp_a1[15]_INST_0_i_3_n_0 ),
        .I2(a1bus_0[7]),
        .O(\rgf_c1bus_wb[7]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c1bus_wb[7]_i_25 
       (.I0(acmd1[0]),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \rgf_c1bus_wb[7]_i_26 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[15]),
        .I3(dctl_sign_f_i_2_n_0),
        .I4(a1bus_0[7]),
        .O(\rgf_c1bus_wb[7]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \rgf_c1bus_wb[7]_i_27 
       (.I0(\rgf_c1bus_wb[7]_i_35_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(b1bus_0[7]),
        .I3(a1bus_0[7]),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \rgf_c1bus_wb[7]_i_28 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[19]_i_42_n_0 ),
        .I4(\rgf_c1bus_wb[27]_i_33_n_0 ),
        .I5(\rgf_c1bus_wb[11]_i_37_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \rgf_c1bus_wb[7]_i_29 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_18_n_0 ),
        .I2(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[7]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[7]_i_3 
       (.I0(bdatr[7]),
        .I1(\mem/read_cyc [0]),
        .I2(bdatr[15]),
        .O(\rgf_c1bus_wb[7]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \rgf_c1bus_wb[7]_i_30 
       (.I0(\rgf_c1bus_wb[28]_i_25_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_28_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_c1bus_wb[7]_i_35 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I2(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_c1bus_wb[7]_i_4 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[7]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[7]_i_5 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [7]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[7]),
        .I4(\rgf_c1bus_wb[7]_i_10_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A888888AAAAAAAA)) 
    \rgf_c1bus_wb[7]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_12_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_39_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF30FF7575)) 
    \rgf_c1bus_wb[7]_i_7 
       (.I0(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_21_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_15_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I4(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_17_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h10FF10FF10FF55FF)) 
    \rgf_c1bus_wb[7]_i_8 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c1bus_wb[7]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[7]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44FF50FF444450FF)) 
    \rgf_c1bus_wb[7]_i_9 
       (.I0(\rgf_c1bus_wb[7]_i_21_n_0 ),
        .I1(\rgf_c1bus_wb[7]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[7]_i_14_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_22_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[8]_i_1 
       (.I0(\rgf_c1bus_wb[8]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[8]),
        .O(c1bus[8]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[8]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[8]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[8]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[8]),
        .O(\rgf_c1bus_wb[8]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[8]_i_12 
       (.I0(a1bus_0[0]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[8]),
        .I4(a1bus_0[8]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[8]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[8]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[8]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[8]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4F444F4F4F444444)) 
    \rgf_c1bus_wb[8]_i_14 
       (.I0(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .I2(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I3(a1bus_0[31]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_23_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h8BBB8B88)) 
    \rgf_c1bus_wb[8]_i_15 
       (.I0(\rgf_c1bus_wb[24]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_24_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_25_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0004F00400F4F0F4)) 
    \rgf_c1bus_wb[8]_i_16 
       (.I0(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[24]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[8]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0B0F)) 
    \rgf_c1bus_wb[8]_i_18 
       (.I0(\rgf_c1bus_wb[24]_i_23_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \rgf_c1bus_wb[8]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_18_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_16_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[8]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [8]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[8]),
        .I4(\rgf_c1bus_wb[8]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047000000FF00)) 
    \rgf_c1bus_wb[8]_i_20 
       (.I0(\rgf_c1bus_wb[28]_i_34_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_37_n_0 ),
        .I3(acmd1[3]),
        .I4(\rgf_c1bus_wb[8]_i_27_n_0 ),
        .I5(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0047FF47FFFFFFFF)) 
    \rgf_c1bus_wb[8]_i_21 
       (.I0(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_26_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_24_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hA3FFA30FA30FA3FF)) 
    \rgf_c1bus_wb[8]_i_22 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[16]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .I4(a1bus_0[8]),
        .I5(b1bus_0[8]),
        .O(\rgf_c1bus_wb[8]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h5F503F3F5F503030)) 
    \rgf_c1bus_wb[8]_i_23 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[8]_i_24 
       (.I0(\rgf_c1bus_wb[29]_i_28_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_33_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_c1bus_wb[8]_i_25 
       (.I0(\rgf_c1bus_wb[20]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[29]_i_43_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_42_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[8]_i_26 
       (.I0(acmd1[3]),
        .I1(a1bus_0[7]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[8]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[8]_i_27 
       (.I0(\rgf_c1bus_wb[29]_i_42_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[12]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[12]_i_30_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[8]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[8]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_7 ),
        .I2(\alu1/div/quo [8]),
        .I3(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .I4(\alu1/div/rem [8]),
        .I5(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[8]_i_5 
       (.I0(\rgf_c1bus_wb[8]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[8]_i_12_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[8]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h8A8A8A8888888A88)) 
    \rgf_c1bus_wb[8]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_15_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[8]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA00EF00EF00)) 
    \rgf_c1bus_wb[8]_i_7 
       (.I0(\rgf_c1bus_wb[8]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEE00F0)) 
    \rgf_c1bus_wb[8]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_24_n_0 ),
        .I2(\rgf_c1bus_wb[8]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[8]_i_17_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c1bus_wb[8]_i_9 
       (.I0(acmd1[3]),
        .I1(a1bus_0[7]),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[8]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEEEEEEEEEEEEE)) 
    \rgf_c1bus_wb[9]_i_1 
       (.I0(\rgf_c1bus_wb[9]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_3_n_0 ),
        .I2(\mem/read_cyc [2]),
        .I3(\mem/read_cyc [1]),
        .I4(\mem/read_cyc [3]),
        .I5(bdatr[9]),
        .O(c1bus[9]));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_c1bus_wb[9]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \rgf_c1bus_wb[9]_i_11 
       (.I0(acmd1[3]),
        .I1(b1bus_0[9]),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I4(a1bus_0[9]),
        .O(\rgf_c1bus_wb[9]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \rgf_c1bus_wb[9]_i_12 
       (.I0(a1bus_0[1]),
        .I1(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_48_n_0 ),
        .I3(b1bus_0[9]),
        .I4(a1bus_0[9]),
        .I5(acmd1[3]),
        .O(\rgf_c1bus_wb[9]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \rgf_c1bus_wb[9]_i_13 
       (.I0(\rgf_c1bus_wb[23]_i_21_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(b1bus_0[9]),
        .I3(\niss_dsp_a1[32]_INST_0_i_3_n_0 ),
        .I4(a1bus_0[9]),
        .I5(\rgf_c1bus_wb[23]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \rgf_c1bus_wb[9]_i_14 
       (.I0(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_23_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_47_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \rgf_c1bus_wb[9]_i_15 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_21_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_34_n_0 ),
        .I5(a1bus_0[31]),
        .O(\rgf_c1bus_wb[9]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0004F00400F4F0F4)) 
    \rgf_c1bus_wb[9]_i_16 
       (.I0(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I1(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[26]_i_19_n_0 ),
        .I5(\rgf_c1bus_wb[25]_i_19_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_c1bus_wb[9]_i_17 
       (.I0(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_16_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \rgf_c1bus_wb[9]_i_18 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[25]_i_22_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \rgf_c1bus_wb[9]_i_19 
       (.I0(\rgf_c1bus_wb[14]_i_22_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_16_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_17_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_24_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \rgf_c1bus_wb[9]_i_2 
       (.I0(\rgf_c1bus_wb[15]_i_4_n_0 ),
        .I1(\alu1/mul/mulh [9]),
        .I2(\rgf_c1bus_wb[15]_i_5_n_0 ),
        .I3(niss_dsp_c1[9]),
        .I4(\rgf_c1bus_wb[9]_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_5_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \rgf_c1bus_wb[9]_i_20 
       (.I0(acmd1[3]),
        .I1(\rgf_c1bus_wb[9]_i_25_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0047FF47FFFFFFFF)) 
    \rgf_c1bus_wb[9]_i_21 
       (.I0(\rgf_c1bus_wb[29]_i_32_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_30_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_26_n_0 ),
        .I5(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hA3FFA30FA30FA3FF)) 
    \rgf_c1bus_wb[9]_i_22 
       (.I0(\niss_dsp_b1[1]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[17]),
        .I2(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I3(acmd1[3]),
        .I4(a1bus_0[9]),
        .I5(b1bus_0[9]),
        .O(\rgf_c1bus_wb[9]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hCFC05F5FCFC05050)) 
    \rgf_c1bus_wb[9]_i_23 
       (.I0(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_32_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_19_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_28_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I5(\rgf_c1bus_wb[17]_i_26_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \rgf_c1bus_wb[9]_i_24 
       (.I0(acmd1[3]),
        .I1(a1bus_0[8]),
        .I2(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .O(\rgf_c1bus_wb[9]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \rgf_c1bus_wb[9]_i_25 
       (.I0(\rgf_c1bus_wb[30]_i_35_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_33_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[29]_i_39_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hE4EEE444)) 
    \rgf_c1bus_wb[9]_i_26 
       (.I0(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_29_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_34_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\rgf_c1bus_wb[13]_i_35_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \rgf_c1bus_wb[9]_i_3 
       (.I0(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[9]_i_9_n_0 ),
        .I5(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_c1bus_wb[9]_i_4 
       (.I0(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_6 ),
        .I2(\alu1/div/rem [9]),
        .I3(\rgf_c1bus_wb[31]_i_21_n_0 ),
        .I4(\alu1/div/quo [9]),
        .I5(\rgf_c1bus_wb[31]_i_22_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \rgf_c1bus_wb[9]_i_5 
       (.I0(\rgf_c1bus_wb[9]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_11_n_0 ),
        .I2(acmd1[0]),
        .I3(\rgf_c1bus_wb[9]_i_12_n_0 ),
        .I4(dctl_sign_f_i_2_n_0),
        .I5(\rgf_c1bus_wb[9]_i_13_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \rgf_c1bus_wb[9]_i_6 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_14_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_15_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAA00EF00EF00)) 
    \rgf_c1bus_wb[9]_i_7 
       (.I0(\rgf_c1bus_wb[9]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_19_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEE00F0)) 
    \rgf_c1bus_wb[9]_i_8 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\rgf_c1bus_wb[25]_i_23_n_0 ),
        .I2(\rgf_c1bus_wb[9]_i_18_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_17_n_0 ),
        .I4(\bdatw[12]_INST_0_i_4_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_20_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF07FF00FF0FFF0F)) 
    \rgf_c1bus_wb[9]_i_9 
       (.I0(acmd1[3]),
        .I1(a1bus_0[8]),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I5(\rgf_c1bus_wb[9]_i_21_n_0 ),
        .O(\rgf_c1bus_wb[9]_i_9_n_0 ));
  CARRY4 \rgf_c1bus_wb_reg[11]_i_10 
       (.CI(\rgf_c1bus_wb_reg[7]_i_23_n_0 ),
        .CO({\rgf_c1bus_wb_reg[11]_i_10_n_0 ,\rgf_c1bus_wb_reg[11]_i_10_n_1 ,\rgf_c1bus_wb_reg[11]_i_10_n_2 ,\rgf_c1bus_wb_reg[11]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a1bus_0[11:8]),
        .O({\rgf_c1bus_wb_reg[11]_i_10_n_4 ,\rgf_c1bus_wb_reg[11]_i_10_n_5 ,\rgf_c1bus_wb_reg[11]_i_10_n_6 ,\rgf_c1bus_wb_reg[11]_i_10_n_7 }),
        .S({\art/add/rgf_c1bus_wb[11]_i_26_n_0 ,\art/add/rgf_c1bus_wb[11]_i_27_n_0 ,\art/add/rgf_c1bus_wb[11]_i_28_n_0 ,\art/add/rgf_c1bus_wb[11]_i_29_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[19]_i_10 
       (.CI(\rgf_c1bus_wb_reg[19]_i_18_n_0 ),
        .CO({\rgf_c1bus_wb_reg[19]_i_10_n_0 ,\rgf_c1bus_wb_reg[19]_i_10_n_1 ,\rgf_c1bus_wb_reg[19]_i_10_n_2 ,\rgf_c1bus_wb_reg[19]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[19]_i_19_n_0 ,\rgf_c1bus_wb[19]_i_20_n_0 ,\rgf_c1bus_wb[19]_i_21_n_0 ,\alu1/asr0 }),
        .O({\rgf_c1bus_wb_reg[19]_i_10_n_4 ,\rgf_c1bus_wb_reg[19]_i_10_n_5 ,\alu1/art/add/tout [18],\rgf_c1bus_wb_reg[19]_i_10_n_7 }),
        .S({\art/add/rgf_c1bus_wb[19]_i_23_n_0 ,\art/add/rgf_c1bus_wb[19]_i_24_n_0 ,\art/add/rgf_c1bus_wb[19]_i_25_n_0 ,\art/add/rgf_c1bus_wb[19]_i_26_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[19]_i_18 
       (.CI(\rgf_c1bus_wb_reg[11]_i_10_n_0 ),
        .CO({\rgf_c1bus_wb_reg[19]_i_18_n_0 ,\rgf_c1bus_wb_reg[19]_i_18_n_1 ,\rgf_c1bus_wb_reg[19]_i_18_n_2 ,\rgf_c1bus_wb_reg[19]_i_18_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a1bus_0[15:12]),
        .O({\rgf_c1bus_wb_reg[19]_i_18_n_4 ,\rgf_c1bus_wb_reg[19]_i_18_n_5 ,\rgf_c1bus_wb_reg[19]_i_18_n_6 ,\rgf_c1bus_wb_reg[19]_i_18_n_7 }),
        .S({\art/add/rgf_c1bus_wb[19]_i_35_n_0 ,\art/add/rgf_c1bus_wb[19]_i_36_n_0 ,\art/add/rgf_c1bus_wb[19]_i_37_n_0 ,\art/add/rgf_c1bus_wb[19]_i_38_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[23]_i_11 
       (.CI(\rgf_c1bus_wb_reg[19]_i_10_n_0 ),
        .CO({\rgf_c1bus_wb_reg[23]_i_11_n_0 ,\rgf_c1bus_wb_reg[23]_i_11_n_1 ,\rgf_c1bus_wb_reg[23]_i_11_n_2 ,\rgf_c1bus_wb_reg[23]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[23]_i_22_n_0 ,\rgf_c1bus_wb[23]_i_23_n_0 ,\rgf_c1bus_wb[23]_i_24_n_0 ,\rgf_c1bus_wb[23]_i_25_n_0 }),
        .O({\rgf_c1bus_wb_reg[23]_i_11_n_4 ,\rgf_c1bus_wb_reg[23]_i_11_n_5 ,\rgf_c1bus_wb_reg[23]_i_11_n_6 ,\rgf_c1bus_wb_reg[23]_i_11_n_7 }),
        .S({\rgf_c1bus_wb[23]_i_26_n_0 ,\art/add/rgf_c1bus_wb[23]_i_27_n_0 ,\art/add/rgf_c1bus_wb[23]_i_28_n_0 ,\art/add/rgf_c1bus_wb[23]_i_29_n_0 }));
  MUXF8 \rgf_c1bus_wb_reg[24]_i_2 
       (.I0(\rgf_c1bus_wb_reg[24]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[24]_i_6_n_0 ),
        .O(\rgf_c1bus_wb_reg[24]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[24]_i_5 
       (.I0(\rgf_c1bus_wb[24]_i_13_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_14_n_0 ),
        .O(\rgf_c1bus_wb_reg[24]_i_5_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  MUXF7 \rgf_c1bus_wb_reg[24]_i_6 
       (.I0(\rgf_c1bus_wb[24]_i_15_n_0 ),
        .I1(\rgf_c1bus_wb[24]_i_16_n_0 ),
        .O(\rgf_c1bus_wb_reg[24]_i_6_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  MUXF8 \rgf_c1bus_wb_reg[26]_i_2 
       (.I0(\rgf_c1bus_wb_reg[26]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[26]_i_6_n_0 ),
        .O(\rgf_c1bus_wb_reg[26]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[26]_i_5 
       (.I0(\rgf_c1bus_wb[26]_i_12_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_13_n_0 ),
        .O(\rgf_c1bus_wb_reg[26]_i_5_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  MUXF7 \rgf_c1bus_wb_reg[26]_i_6 
       (.I0(\rgf_c1bus_wb[26]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_15_n_0 ),
        .O(\rgf_c1bus_wb_reg[26]_i_6_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  CARRY4 \rgf_c1bus_wb_reg[27]_i_10 
       (.CI(\rgf_c1bus_wb_reg[23]_i_11_n_0 ),
        .CO({\rgf_c1bus_wb_reg[27]_i_10_n_0 ,\rgf_c1bus_wb_reg[27]_i_10_n_1 ,\rgf_c1bus_wb_reg[27]_i_10_n_2 ,\rgf_c1bus_wb_reg[27]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[27]_i_17_n_0 ,\rgf_c1bus_wb[27]_i_18_n_0 ,\rgf_c1bus_wb[27]_i_19_n_0 ,\rgf_c1bus_wb[27]_i_20_n_0 }),
        .O({\rgf_c1bus_wb_reg[27]_i_10_n_4 ,\rgf_c1bus_wb_reg[27]_i_10_n_5 ,\rgf_c1bus_wb_reg[27]_i_10_n_6 ,\rgf_c1bus_wb_reg[27]_i_10_n_7 }),
        .S({\art/add/rgf_c1bus_wb[27]_i_21_n_0 ,\art/add/rgf_c1bus_wb[27]_i_22_n_0 ,\art/add/rgf_c1bus_wb[27]_i_23_n_0 ,\art/add/rgf_c1bus_wb[27]_i_24_n_0 }));
  MUXF8 \rgf_c1bus_wb_reg[30]_i_2 
       (.I0(\rgf_c1bus_wb_reg[30]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb_reg[30]_i_6_n_0 ),
        .O(\rgf_c1bus_wb_reg[30]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[30]_i_5 
       (.I0(\rgf_c1bus_wb[30]_i_14_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_15_n_0 ),
        .O(\rgf_c1bus_wb_reg[30]_i_5_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  MUXF7 \rgf_c1bus_wb_reg[30]_i_6 
       (.I0(\rgf_c1bus_wb[30]_i_16_n_0 ),
        .I1(\rgf_c1bus_wb[30]_i_17_n_0 ),
        .O(\rgf_c1bus_wb_reg[30]_i_6_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  CARRY4 \rgf_c1bus_wb_reg[31]_i_11 
       (.CI(\rgf_c1bus_wb_reg[27]_i_10_n_0 ),
        .CO({\rgf_c1bus_wb_reg[31]_i_11_n_0 ,\rgf_c1bus_wb_reg[31]_i_11_n_1 ,\rgf_c1bus_wb_reg[31]_i_11_n_2 ,\rgf_c1bus_wb_reg[31]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rgf_c1bus_wb[31]_i_25_n_0 ,\rgf_c1bus_wb[31]_i_26_n_0 ,\rgf_c1bus_wb[31]_i_27_n_0 ,\rgf_c1bus_wb[31]_i_28_n_0 }),
        .O({\rgf_c1bus_wb_reg[31]_i_11_n_4 ,\rgf_c1bus_wb_reg[31]_i_11_n_5 ,\rgf_c1bus_wb_reg[31]_i_11_n_6 ,\rgf_c1bus_wb_reg[31]_i_11_n_7 }),
        .S({\art/add/rgf_c1bus_wb[31]_i_29_n_0 ,\art/add/rgf_c1bus_wb[31]_i_30_n_0 ,\art/add/rgf_c1bus_wb[31]_i_31_n_0 ,\art/add/rgf_c1bus_wb[31]_i_32_n_0 }));
  MUXF8 \rgf_c1bus_wb_reg[31]_i_2 
       (.I0(\rgf_c1bus_wb_reg[31]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb_reg[31]_i_7_n_0 ),
        .O(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .S(acmd1[0]));
  MUXF7 \rgf_c1bus_wb_reg[31]_i_6 
       (.I0(\rgf_c1bus_wb[31]_i_17_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_18_n_0 ),
        .O(\rgf_c1bus_wb_reg[31]_i_6_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  MUXF7 \rgf_c1bus_wb_reg[31]_i_7 
       (.I0(\rgf_c1bus_wb[31]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_20_n_0 ),
        .O(\rgf_c1bus_wb_reg[31]_i_7_n_0 ),
        .S(dctl_sign_f_i_2_n_0));
  CARRY4 \rgf_c1bus_wb_reg[3]_i_20 
       (.CI(\<const0> ),
        .CO({\rgf_c1bus_wb_reg[3]_i_20_n_0 ,\rgf_c1bus_wb_reg[3]_i_20_n_1 ,\rgf_c1bus_wb_reg[3]_i_20_n_2 ,\rgf_c1bus_wb_reg[3]_i_20_n_3 }),
        .CYINIT(\rgf_c1bus_wb[3]_i_26_n_0 ),
        .DI(a1bus_0[3:0]),
        .O({\rgf_c1bus_wb_reg[3]_i_20_n_4 ,\rgf_c1bus_wb_reg[3]_i_20_n_5 ,\rgf_c1bus_wb_reg[3]_i_20_n_6 ,\rgf_c1bus_wb_reg[3]_i_20_n_7 }),
        .S({\art/add/rgf_c1bus_wb[3]_i_27_n_0 ,\art/add/rgf_c1bus_wb[3]_i_28_n_0 ,\art/add/rgf_c1bus_wb[3]_i_29_n_0 ,\art/add/rgf_c1bus_wb[3]_i_30_n_0 }));
  CARRY4 \rgf_c1bus_wb_reg[7]_i_23 
       (.CI(\rgf_c1bus_wb_reg[3]_i_20_n_0 ),
        .CO({\rgf_c1bus_wb_reg[7]_i_23_n_0 ,\rgf_c1bus_wb_reg[7]_i_23_n_1 ,\rgf_c1bus_wb_reg[7]_i_23_n_2 ,\rgf_c1bus_wb_reg[7]_i_23_n_3 }),
        .CYINIT(\<const0> ),
        .DI(a1bus_0[7:4]),
        .O({\rgf_c1bus_wb_reg[7]_i_23_n_4 ,\rgf_c1bus_wb_reg[7]_i_23_n_5 ,\rgf_c1bus_wb_reg[7]_i_23_n_6 ,\rgf_c1bus_wb_reg[7]_i_23_n_7 }),
        .S({\art/add/rgf_c1bus_wb[7]_i_31_n_0 ,\art/add/rgf_c1bus_wb[7]_i_32_n_0 ,\art/add/rgf_c1bus_wb[7]_i_33_n_0 ,\art/add/rgf_c1bus_wb[7]_i_34_n_0 }));
  LUT6 #(
    .INIT(64'hDDDDDDD0DDDDDDDD)) 
    \rgf_selc0_rn_wb[0]_i_1 
       (.I0(stat[2]),
        .I1(\rgf_selc0_rn_wb[0]_i_2_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_3_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_4_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_5_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_6_n_0 ),
        .O(ctl_selc0_rn));
  LUT6 #(
    .INIT(64'h0000000040000000)) 
    \rgf_selc0_rn_wb[0]_i_10 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [13]),
        .I4(stat[0]),
        .I5(stat[1]),
        .O(\rgf_selc0_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h11110000FFF10000)) 
    \rgf_selc0_rn_wb[0]_i_11 
       (.I0(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I4(\fch/ir0 [3]),
        .I5(\rgf_selc0_rn_wb[0]_i_18_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFF70FFFF)) 
    \rgf_selc0_rn_wb[0]_i_12 
       (.I0(crdy),
        .I1(div_crdy0),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hABBBBBBBAAAAAAAA)) 
    \rgf_selc0_rn_wb[0]_i_13 
       (.I0(\ccmd[4]_INST_0_i_2_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_19_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_20_n_0 ),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [0]),
        .I5(\rgf_selc0_rn_wb[0]_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00FF00E0000000E0)) 
    \rgf_selc0_rn_wb[0]_i_14 
       (.I0(\rgf_selc0_rn_wb[0]_i_22_n_0 ),
        .I1(\fch/ir0 [13]),
        .I2(\rgf_selc0_rn_wb[0]_i_23_n_0 ),
        .I3(\fch/ir0 [15]),
        .I4(\fch/ir0 [14]),
        .I5(\bdatw[31]_INST_0_i_77_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h000D0D0D000D000D)) 
    \rgf_selc0_rn_wb[0]_i_15 
       (.I0(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_24_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_25_n_0 ),
        .I3(\fch/ir0 [3]),
        .I4(\rgf_selc0_rn_wb[0]_i_26_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h000000005555FFDF)) 
    \rgf_selc0_rn_wb[0]_i_16 
       (.I0(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .I2(\ccmd[2]_INST_0_i_12_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_28_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_29_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_30_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc0_rn_wb[0]_i_17 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [10]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[0]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \rgf_selc0_rn_wb[0]_i_18 
       (.I0(\fch/ir0 [7]),
        .I1(div_crdy0),
        .I2(crdy),
        .O(\rgf_selc0_rn_wb[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \rgf_selc0_rn_wb[0]_i_19 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .O(\rgf_selc0_rn_wb[0]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc0_rn_wb[0]_i_2 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\fch/ir0 [15]),
        .I3(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_selc0_rn_wb[0]_i_20 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(brdy),
        .I3(\fch/ir0 [7]),
        .O(\rgf_selc0_rn_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hDDDFDFFFDFFFDFFF)) 
    \rgf_selc0_rn_wb[0]_i_21 
       (.I0(\fch/ir0 [3]),
        .I1(\rgf_selc0_rn_wb[0]_i_31_n_0 ),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [4]),
        .I4(brdy),
        .I5(\fch/ir0 [0]),
        .O(\rgf_selc0_rn_wb[0]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h9A)) 
    \rgf_selc0_rn_wb[0]_i_22 
       (.I0(\fch/ir0 [11]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir0 [12]),
        .O(\rgf_selc0_rn_wb[0]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hB847FFFF)) 
    \rgf_selc0_rn_wb[0]_i_23 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir0 [12]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [13]),
        .O(\rgf_selc0_rn_wb[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hFF5577FCF7DFFFFD)) 
    \rgf_selc0_rn_wb[0]_i_24 
       (.I0(\fch/ir0 [0]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [7]),
        .O(\rgf_selc0_rn_wb[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0007000000000000)) 
    \rgf_selc0_rn_wb[0]_i_25 
       (.I0(\fch/ir0 [8]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [3]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h00000000C0000404)) 
    \rgf_selc0_rn_wb[0]_i_26 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [11]),
        .O(\rgf_selc0_rn_wb[0]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'h5515)) 
    \rgf_selc0_rn_wb[0]_i_27 
       (.I0(\fch/ir0 [8]),
        .I1(brdy),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .O(\rgf_selc0_rn_wb[0]_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hABFB)) 
    \rgf_selc0_rn_wb[0]_i_28 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [0]),
        .O(\rgf_selc0_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hB0B0A0A030FF0000)) 
    \rgf_selc0_rn_wb[0]_i_29 
       (.I0(\rgf_selc0_rn_wb[0]_i_32_n_0 ),
        .I1(\ccmd[1]_INST_0_i_13_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_20_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_17_n_0 ),
        .I4(\fch/ir0 [0]),
        .I5(\fch/ir0 [3]),
        .O(\rgf_selc0_rn_wb[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \rgf_selc0_rn_wb[0]_i_3 
       (.I0(\rgf_selc0_rn_wb[0]_i_8_n_0 ),
        .I1(\ccmd[1]_INST_0_i_6_n_0 ),
        .I2(\rgf_selc0_rn_wb[0]_i_9_n_0 ),
        .I3(brdy),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [1]),
        .O(\rgf_selc0_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0045000000000000)) 
    \rgf_selc0_rn_wb[0]_i_30 
       (.I0(\fch/ir0 [14]),
        .I1(brdy),
        .I2(\fch/ir0 [1]),
        .I3(\badr[31]_INST_0_i_133_n_0 ),
        .I4(\fadr[15]_INST_0_i_12_n_0 ),
        .I5(\stat[0]_i_7__0_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[0]_i_31 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .O(\rgf_selc0_rn_wb[0]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_selc0_rn_wb[0]_i_32 
       (.I0(brdy),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [6]),
        .O(\rgf_selc0_rn_wb[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h88A8AAAA88888888)) 
    \rgf_selc0_rn_wb[0]_i_4 
       (.I0(\rgf_selc0_rn_wb[0]_i_10_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_11_n_0 ),
        .I2(\fch/ir0 [3]),
        .I3(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc0_rn_wb[0]_i_13_n_0 ),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h8A888A888A88AAAA)) 
    \rgf_selc0_rn_wb[0]_i_5 
       (.I0(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_14_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\ccmd[3]_INST_0_i_3_n_0 ),
        .I5(\rgf_selc0_rn_wb[0]_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h3333313333333111)) 
    \rgf_selc0_rn_wb[0]_i_6 
       (.I0(stat[1]),
        .I1(stat[2]),
        .I2(\rgf_selc0_rn_wb[0]_i_7_n_0 ),
        .I3(stat[0]),
        .I4(\fch/ir0 [15]),
        .I5(\rgf_selc0_rn_wb[0]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \rgf_selc0_rn_wb[0]_i_7 
       (.I0(\stat[2]_i_8__0_n_0 ),
        .I1(\fadr[15]_INST_0_i_12_n_0 ),
        .I2(\fch/ir0 [1]),
        .I3(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [6]),
        .O(\rgf_selc0_rn_wb[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \rgf_selc0_rn_wb[0]_i_8 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(\rgf_selc0_rn_wb[0]_i_17_n_0 ),
        .O(\rgf_selc0_rn_wb[0]_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \rgf_selc0_rn_wb[0]_i_9 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [0]),
        .O(\rgf_selc0_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4544555545444544)) 
    \rgf_selc0_rn_wb[1]_i_1 
       (.I0(stat[2]),
        .I1(\rgf_selc0_rn_wb[1]_i_2_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_3_n_0 ),
        .I3(\ccmd[1]_INST_0_i_6_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_4_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h1010000010FF0000)) 
    \rgf_selc0_rn_wb[1]_i_10 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\rgf_selc0_rn_wb[1]_i_18_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I4(\fch/ir0 [4]),
        .I5(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFFFFFAAAAFFFF)) 
    \rgf_selc0_rn_wb[1]_i_11 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0202020202028A02)) 
    \rgf_selc0_rn_wb[1]_i_12 
       (.I0(\stat[2]_i_8__0_n_0 ),
        .I1(brdy),
        .I2(\rgf_selc0_rn_wb[1]_i_19_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_20_n_0 ),
        .I4(\fch/ir0 [6]),
        .I5(\bdatw[8]_INST_0_i_21_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hC000040400000000)) 
    \rgf_selc0_rn_wb[1]_i_13 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_selc0_rn_wb[1]_i_21_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [4]),
        .O(\rgf_selc0_rn_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00103010)) 
    \rgf_selc0_rn_wb[1]_i_14 
       (.I0(\rgf_selc0_rn_wb[1]_i_22_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [7]),
        .I4(\rgf_selc0_rn_wb[1]_i_23_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_24_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc0_rn_wb[1]_i_15 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [7]),
        .I2(brdy),
        .O(\rgf_selc0_rn_wb[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[1]_i_16 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .O(\rgf_selc0_rn_wb[1]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[1]_i_17 
       (.I0(\fch/ir0 [6]),
        .I1(brdy),
        .O(\rgf_selc0_rn_wb[1]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \rgf_selc0_rn_wb[1]_i_18 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [11]),
        .O(\rgf_selc0_rn_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    \rgf_selc0_rn_wb[1]_i_19 
       (.I0(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [1]),
        .O(\rgf_selc0_rn_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h1111111011101110)) 
    \rgf_selc0_rn_wb[1]_i_2 
       (.I0(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I1(\ccmd[3]_INST_0_i_3_n_0 ),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_6_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_8_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \rgf_selc0_rn_wb[1]_i_20 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[1]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_rn_wb[1]_i_21 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .O(\rgf_selc0_rn_wb[1]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hF7FFFF7B)) 
    \rgf_selc0_rn_wb[1]_i_22 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [4]),
        .O(\rgf_selc0_rn_wb[1]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hBF77)) 
    \rgf_selc0_rn_wb[1]_i_23 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0007000003FF0000)) 
    \rgf_selc0_rn_wb[1]_i_24 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [10]),
        .O(\rgf_selc0_rn_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h000000005D5D555D)) 
    \rgf_selc0_rn_wb[1]_i_3 
       (.I0(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_9_n_0 ),
        .I2(\rgf_selc0_rn_wb[1]_i_10_n_0 ),
        .I3(\fch/ir0 [4]),
        .I4(\rgf_selc0_rn_wb[1]_i_11_n_0 ),
        .I5(\rgf_selc0_rn_wb[1]_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0D0DDDDDDD0DD)) 
    \rgf_selc0_rn_wb[1]_i_4 
       (.I0(\fch/ir0 [9]),
        .I1(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I2(\ccmd[3]_INST_0_i_3_n_0 ),
        .I3(\rgf_selc0_rn_wb[1]_i_13_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\rgf_selc0_rn_wb[1]_i_14_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc0_rn_wb[1]_i_5 
       (.I0(stat[0]),
        .I1(stat[1]),
        .O(\rgf_selc0_rn_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000000C000A0A)) 
    \rgf_selc0_rn_wb[1]_i_6 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [8]),
        .I3(\rgf_selc0_rn_wb[1]_i_15_n_0 ),
        .I4(\fch/ir0 [9]),
        .I5(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000040F0F0F0F0)) 
    \rgf_selc0_rn_wb[1]_i_7 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [3]),
        .I4(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I5(\fch/ir0 [9]),
        .O(\rgf_selc0_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF00400000004000)) 
    \rgf_selc0_rn_wb[1]_i_8 
       (.I0(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I1(\fch/ir0 [4]),
        .I2(\ccmd[3]_INST_0_i_15_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [1]),
        .O(\rgf_selc0_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF700F7F7FFFFFFFF)) 
    \rgf_selc0_rn_wb[1]_i_9 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [3]),
        .I2(\rgf_selc0_rn_wb[2]_i_13_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I4(\fch/ir0 [4]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \rgf_selc0_rn_wb[2]_i_1 
       (.I0(stat[2]),
        .I1(\rgf_selc0_rn_wb[2]_i_2_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_3_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_4_n_0 ),
        .I4(\fch/ir0 [10]),
        .I5(\rgf_selc0_rn_wb[2]_i_5_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hE33FFF1EFFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_10 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [2]),
        .O(\rgf_selc0_rn_wb[2]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \rgf_selc0_rn_wb[2]_i_11 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    \rgf_selc0_rn_wb[2]_i_12 
       (.I0(\rgf_selc0_rn_wb[2]_i_23_n_0 ),
        .I1(\ccmd[3]_INST_0_i_7_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_24_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .I4(\fch/ir0 [8]),
        .I5(\fch/ir0 [7]),
        .O(\rgf_selc0_rn_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFEFFFBFFFBFFF)) 
    \rgf_selc0_rn_wb[2]_i_13 
       (.I0(\ccmd[4]_INST_0_i_2_n_0 ),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [6]),
        .I3(brdy),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [4]),
        .O(\rgf_selc0_rn_wb[2]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h9FFF9FBF)) 
    \rgf_selc0_rn_wb[2]_i_14 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .O(\rgf_selc0_rn_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \rgf_selc0_rn_wb[2]_i_15 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [7]),
        .I5(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h77775777FFFFDFFF)) 
    \rgf_selc0_rn_wb[2]_i_16 
       (.I0(\rgf_selc0_rn_wb[2]_i_26_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [5]),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(\fch/ir0 [2]),
        .O(\rgf_selc0_rn_wb[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_17 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\ccmd[4]_INST_0_i_2_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [10]),
        .I5(\rgf_selc0_wb[1]_i_3_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h00008B8800000000)) 
    \rgf_selc0_rn_wb[2]_i_18 
       (.I0(\rgf_selc0_rn_wb[2]_i_27_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\rgf_selc0_rn_wb[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h000000003EFFFEFF)) 
    \rgf_selc0_rn_wb[2]_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [5]),
        .I4(\fch/ir0 [6]),
        .I5(\fch/ir0 [9]),
        .O(\rgf_selc0_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h000000DD000F0000)) 
    \rgf_selc0_rn_wb[2]_i_2 
       (.I0(\rgf_selc0_rn_wb[2]_i_6_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_7_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_8_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(stat[1]),
        .I5(stat[0]),
        .O(\rgf_selc0_rn_wb[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00202222)) 
    \rgf_selc0_rn_wb[2]_i_20 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .O(\rgf_selc0_rn_wb[2]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFDFDFDDD)) 
    \rgf_selc0_rn_wb[2]_i_21 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [8]),
        .O(\rgf_selc0_rn_wb[2]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFECCFFCF)) 
    \rgf_selc0_rn_wb[2]_i_22 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [5]),
        .O(\rgf_selc0_rn_wb[2]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_selc0_rn_wb[2]_i_23 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [2]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [3]),
        .O(\rgf_selc0_rn_wb[2]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc0_rn_wb[2]_i_24 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [14]),
        .O(\rgf_selc0_rn_wb[2]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[2]_i_25 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [9]),
        .O(\rgf_selc0_rn_wb[2]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc0_rn_wb[2]_i_26 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [11]),
        .O(\rgf_selc0_rn_wb[2]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc0_rn_wb[2]_i_27 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [6]),
        .I4(brdy),
        .O(\rgf_selc0_rn_wb[2]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4044404055555555)) 
    \rgf_selc0_rn_wb[2]_i_3 
       (.I0(\fch/ir0 [15]),
        .I1(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_9_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_10_n_0 ),
        .I4(\rgf_selc0_rn_wb[2]_i_11_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \rgf_selc0_rn_wb[2]_i_4 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .O(\rgf_selc0_rn_wb[2]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_rn_wb[2]_i_5 
       (.I0(stat[1]),
        .I1(stat[0]),
        .O(\rgf_selc0_rn_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF700F7F7FFFFFFFF)) 
    \rgf_selc0_rn_wb[2]_i_6 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [2]),
        .I2(\rgf_selc0_rn_wb[2]_i_13_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_12_n_0 ),
        .I4(\fch/ir0 [5]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF50705050)) 
    \rgf_selc0_rn_wb[2]_i_7 
       (.I0(\rgf_selc0_rn_wb[1]_i_11_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_14_n_0 ),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [6]),
        .I4(brdy),
        .I5(\rgf_selc0_rn_wb[2]_i_15_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000000022222022)) 
    \rgf_selc0_rn_wb[2]_i_8 
       (.I0(\rgf_selc0_rn_wb[2]_i_16_n_0 ),
        .I1(\ccmd[4]_INST_0_i_1_n_0 ),
        .I2(\rgf_selc0_rn_wb[2]_i_17_n_0 ),
        .I3(\fch/ir0 [2]),
        .I4(\fch/ir0 [3]),
        .I5(\rgf_selc0_rn_wb[2]_i_18_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \rgf_selc0_rn_wb[2]_i_9 
       (.I0(\rgf_selc0_rn_wb[2]_i_19_n_0 ),
        .I1(\rgf_selc0_rn_wb[2]_i_20_n_0 ),
        .I2(\fch/ir0 [5]),
        .I3(\rgf_selc0_rn_wb[2]_i_21_n_0 ),
        .I4(\ccmd[2]_INST_0_i_12_n_0 ),
        .I5(\rgf_selc0_rn_wb[2]_i_22_n_0 ),
        .O(\rgf_selc0_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    rgf_selc0_stat_i_1
       (.I0(fch_term),
        .I1(rst_n),
        .O(rgf_selc0_stat_i_1_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc0_stat_i_2
       (.I0(ctl_selc0[1]),
        .I1(ctl_selc0[0]),
        .O(rgf_selc0_stat_i_2_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc0_stat_i_3
       (.I0(fch_wrbufn0),
        .O(\rgf/rctl/p_2_in ));
  LUT5 #(
    .INIT(32'hFFFFE200)) 
    rgf_selc0_stat_i_4
       (.I0(\fch/ir0_id_fl [20]),
        .I1(\fch/fch_term_fl ),
        .I2(\ir0_id_fl[20]_i_2_n_0 ),
        .I3(\fch/rst_n_fl ),
        .I4(\fch/fch_irq_req_fl ),
        .O(fch_wrbufn0));
  LUT6 #(
    .INIT(64'hFFFFFFFF282A8A2A)) 
    \rgf_selc0_wb[0]_i_1 
       (.I0(\rgf_selc0_wb[0]_i_2_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [13]),
        .I5(\rgf_selc0_wb[0]_i_3_n_0 ),
        .O(ctl_selc0[0]));
  LUT6 #(
    .INIT(64'h00000000A80AA8AA)) 
    \rgf_selc0_wb[0]_i_10 
       (.I0(\rgf_selc0_wb[0]_i_13_n_0 ),
        .I1(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [9]),
        .I4(\ccmd[2]_INST_0_i_10_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_14_n_0 ),
        .O(\rgf_selc0_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF9F9FFF7FBFBFBBE)) 
    \rgf_selc0_wb[0]_i_11 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [6]),
        .I2(stat[1]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [4]),
        .O(\rgf_selc0_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF00FF80FF008080)) 
    \rgf_selc0_wb[0]_i_12 
       (.I0(\fch/ir0 [6]),
        .I1(\ccmd[3]_INST_0_i_15_n_0 ),
        .I2(\ccmd[2]_INST_0_i_16_n_0 ),
        .I3(\rgf_selc0_rn_wb[2]_i_26_n_0 ),
        .I4(stat[1]),
        .I5(\rgf_selc0_wb[1]_i_25_n_0 ),
        .O(\rgf_selc0_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF2AFFAAFFFFFFFF)) 
    \rgf_selc0_wb[0]_i_13 
       (.I0(\fch/ir0 [9]),
        .I1(\rgf_selc0_wb[0]_i_15_n_0 ),
        .I2(\rgf_selc0_wb[0]_i_16_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [4]),
        .I5(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0080000000000000)) 
    \rgf_selc0_wb[0]_i_14 
       (.I0(\ccmd[0]_INST_0_i_14_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_17_n_0 ),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [7]),
        .I5(brdy),
        .O(\rgf_selc0_wb[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[0]_i_15 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [5]),
        .O(\rgf_selc0_wb[0]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_wb[0]_i_16 
       (.I0(\fch/ir0 [3]),
        .I1(brdy),
        .O(\rgf_selc0_wb[0]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_wb[0]_i_17 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [3]),
        .O(\rgf_selc0_wb[0]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \rgf_selc0_wb[0]_i_2 
       (.I0(stat[2]),
        .I1(stat[0]),
        .I2(stat[1]),
        .I3(\fch/ir0 [15]),
        .O(\rgf_selc0_wb[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000E00)) 
    \rgf_selc0_wb[0]_i_3 
       (.I0(\rgf_selc0_wb[0]_i_4_n_0 ),
        .I1(stat[0]),
        .I2(\rgf_selc0_wb[0]_i_5_n_0 ),
        .I3(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I4(stat[2]),
        .I5(\fch/ir0 [15]),
        .O(\rgf_selc0_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8888B888BBBBBBBB)) 
    \rgf_selc0_wb[0]_i_4 
       (.I0(\rgf_selc0_wb[0]_i_6_n_0 ),
        .I1(\rgf_selc0_wb[0]_i_7_n_0 ),
        .I2(stat[1]),
        .I3(\fch/ir0 [10]),
        .I4(\rgf_selc0_wb[0]_i_8_n_0 ),
        .I5(\rgf_selc0_wb[0]_i_9_n_0 ),
        .O(\rgf_selc0_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0D0F0F0F0D000)) 
    \rgf_selc0_wb[0]_i_5 
       (.I0(\fch/ir0 [8]),
        .I1(\rgf_selc0_wb[0]_i_10_n_0 ),
        .I2(stat[0]),
        .I3(\fch/ir0 [11]),
        .I4(stat[1]),
        .I5(\rgf_selc0_wb[1]_i_17_n_0 ),
        .O(\rgf_selc0_wb[0]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4000)) 
    \rgf_selc0_wb[0]_i_6 
       (.I0(\rgf_selc0_wb[0]_i_11_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [10]),
        .I4(\rgf_selc0_wb[0]_i_12_n_0 ),
        .O(\rgf_selc0_wb[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hF0F000D0)) 
    \rgf_selc0_wb[0]_i_7 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hEFFF8AAAFFFFDFFF)) 
    \rgf_selc0_wb[0]_i_8 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(brdy),
        .I4(\fch/ir0 [9]),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\rgf_selc0_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFCC0FFFB)) 
    \rgf_selc0_wb[0]_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [11]),
        .I5(stat[1]),
        .O(\rgf_selc0_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h1111111F11111111)) 
    \rgf_selc0_wb[1]_i_1 
       (.I0(\rgf_selc0_wb[1]_i_2_n_0 ),
        .I1(stat[2]),
        .I2(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(\rgf_selc0_wb[1]_i_4_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_5_n_0 ),
        .O(ctl_selc0[1]));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_10 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[1]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_wb[1]_i_11 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [8]),
        .O(\rgf_selc0_wb[1]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc0_wb[1]_i_12 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [12]),
        .O(\rgf_selc0_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF000E0F0E)) 
    \rgf_selc0_wb[1]_i_13 
       (.I0(\fch/ir0 [15]),
        .I1(\rgf_selc0_wb[1]_i_22_n_0 ),
        .I2(stat[0]),
        .I3(\fch/ir0 [12]),
        .I4(\rgf_selc0_wb[1]_i_23_n_0 ),
        .I5(\fch/ir0 [14]),
        .O(\rgf_selc0_wb[1]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h1FFF9BBB)) 
    \rgf_selc0_wb[1]_i_14 
       (.I0(\fch/ir0 [1]),
        .I1(\fch/ir0 [3]),
        .I2(stat[0]),
        .I3(brdy),
        .I4(\fch/ir0 [0]),
        .O(\rgf_selc0_wb[1]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \rgf_selc0_wb[1]_i_15 
       (.I0(\fch/ir0 [6]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hD7)) 
    \rgf_selc0_wb[1]_i_16 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .O(\rgf_selc0_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFB3B)) 
    \rgf_selc0_wb[1]_i_17 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_24_n_0 ),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\rgf_selc0_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h5151510055555555)) 
    \rgf_selc0_wb[1]_i_18 
       (.I0(stat[0]),
        .I1(\rgf_selc0_wb[1]_i_25_n_0 ),
        .I2(\ccmd[1]_INST_0_i_13_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(\fch/ir0 [10]),
        .O(\rgf_selc0_wb[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBBAAAAAAAAA)) 
    \rgf_selc0_wb[1]_i_19 
       (.I0(\rgf_selc0_wb[1]_i_26_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [10]),
        .I5(\rgf_selc0_wb[1]_i_28_n_0 ),
        .O(\rgf_selc0_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EFEFFFEF)) 
    \rgf_selc0_wb[1]_i_2 
       (.I0(\fch/ir0 [11]),
        .I1(stat[1]),
        .I2(\rgf_selc0_wb[1]_i_6_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_7_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_8_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_9_n_0 ),
        .O(\rgf_selc0_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF440044F0)) 
    \rgf_selc0_wb[1]_i_20 
       (.I0(\rgf_selc0_wb[1]_i_29_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .I4(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I5(\ccmd[2]_INST_0_i_17_n_0 ),
        .O(\rgf_selc0_wb[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFABAAAAAAAA)) 
    \rgf_selc0_wb[1]_i_21 
       (.I0(\rgf_selc0_wb[1]_i_30_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_31_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_32_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\rgf_selc0_wb[1]_i_33_n_0 ),
        .O(\rgf_selc0_wb[1]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc0_wb[1]_i_22 
       (.I0(\fch/ir0 [13]),
        .I1(\rgf/sreg/sr [6]),
        .O(\rgf_selc0_wb[1]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_selc0_wb[1]_i_23 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir0 [13]),
        .I2(\rgf/sreg/sr [4]),
        .O(\rgf_selc0_wb[1]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h40444444)) 
    \rgf_selc0_wb[1]_i_24 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [9]),
        .I3(crdy),
        .I4(div_crdy0),
        .O(\rgf_selc0_wb[1]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc0_wb[1]_i_25 
       (.I0(\fch/ir0 [7]),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf_selc0_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFE2FF)) 
    \rgf_selc0_wb[1]_i_26 
       (.I0(\rgf_selc0_wb[1]_i_34_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\rgf_selc0_wb[1]_i_35_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [15]),
        .I5(stat[1]),
        .O(\rgf_selc0_wb[1]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \rgf_selc0_wb[1]_i_27 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(stat[0]),
        .I3(\fch/ir0 [12]),
        .O(\rgf_selc0_wb[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h55555555FC000000)) 
    \rgf_selc0_wb[1]_i_28 
       (.I0(\rgf_selc0_wb[1]_i_36_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [9]),
        .O(\rgf_selc0_wb[1]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h7F7C377FFFFF37FF)) 
    \rgf_selc0_wb[1]_i_29 
       (.I0(brdy),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [5]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [9]),
        .O(\rgf_selc0_wb[1]_i_29_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_3 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [5]),
        .O(\rgf_selc0_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0002020002020202)) 
    \rgf_selc0_wb[1]_i_30 
       (.I0(\fch/ir0 [15]),
        .I1(stat[1]),
        .I2(stat[0]),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [14]),
        .I5(\fch/ir0 [13]),
        .O(\rgf_selc0_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDFDFDFD)) 
    \rgf_selc0_wb[1]_i_31 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [9]),
        .I3(brdy),
        .I4(\bbus_o[5]_INST_0_i_25_n_0 ),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\rgf_selc0_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \rgf_selc0_wb[1]_i_32 
       (.I0(\fch/ir0 [12]),
        .I1(\rgf_selc0_wb[1]_i_37_n_0 ),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [7]),
        .I4(\rgf_selc0_wb[1]_i_38_n_0 ),
        .I5(\fch_irq_lev[1]_i_3_n_0 ),
        .O(\rgf_selc0_wb[1]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000004044444444)) 
    \rgf_selc0_wb[1]_i_33 
       (.I0(\fch/ir0 [15]),
        .I1(stat[1]),
        .I2(\rgf_selc0_rn_wb[1]_i_7_n_0 ),
        .I3(\rgf_selc0_rn_wb[0]_i_27_n_0 ),
        .I4(\rgf_selc0_wb[1]_i_27_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\rgf_selc0_wb[1]_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF530)) 
    \rgf_selc0_wb[1]_i_34 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [14]),
        .O(\rgf_selc0_wb[1]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h510B015B)) 
    \rgf_selc0_wb[1]_i_35 
       (.I0(\fch/ir0 [13]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir0 [14]),
        .I3(\rgf/sreg/sr [7]),
        .I4(\rgf/sreg/sr [5]),
        .O(\rgf_selc0_wb[1]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h2020A0882820A0A2)) 
    \rgf_selc0_wb[1]_i_36 
       (.I0(\rgf_selc0_wb[1]_i_39_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [3]),
        .O(\rgf_selc0_wb[1]_i_36_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc0_wb[1]_i_37 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [2]),
        .O(\rgf_selc0_wb[1]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h00002F0000000000)) 
    \rgf_selc0_wb[1]_i_38 
       (.I0(brdy),
        .I1(stat[0]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [8]),
        .I5(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .O(\rgf_selc0_wb[1]_i_38_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc0_wb[1]_i_39 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .O(\rgf_selc0_wb[1]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    \rgf_selc0_wb[1]_i_4 
       (.I0(stat[1]),
        .I1(\fch/ir0 [9]),
        .I2(\rgf_selc0_wb[1]_i_10_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_11_n_0 ),
        .I4(\fch/ir0 [1]),
        .I5(stat[2]),
        .O(\rgf_selc0_wb[1]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc0_wb[1]_i_5 
       (.I0(\fch/ir0 [2]),
        .I1(stat[0]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [3]),
        .I4(\rgf_selc0_wb[1]_i_12_n_0 ),
        .O(\rgf_selc0_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAE)) 
    \rgf_selc0_wb[1]_i_6 
       (.I0(\rgf_selc0_wb[1]_i_13_n_0 ),
        .I1(\stat[0]_i_8__0_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_14_n_0 ),
        .I3(\fch/ir0 [12]),
        .I4(\fch/ir0 [15]),
        .I5(\fch/ir0 [13]),
        .O(\rgf_selc0_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEF0)) 
    \rgf_selc0_wb[1]_i_7 
       (.I0(\rgf_selc0_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc0_wb[1]_i_16_n_0 ),
        .I2(\rgf_selc0_wb[1]_i_17_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_18_n_0 ),
        .I4(\fch/ir0 [15]),
        .I5(\ccmd[0]_INST_0_i_20_n_0 ),
        .O(\rgf_selc0_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000087FFFFFFFF)) 
    \rgf_selc0_wb[1]_i_8 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir0 [12]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir0 [13]),
        .I4(stat[0]),
        .I5(\fch/ir0 [14]),
        .O(\rgf_selc0_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40005555)) 
    \rgf_selc0_wb[1]_i_9 
       (.I0(\rgf_selc0_wb[1]_i_19_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\bbus_o[5]_INST_0_i_9_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_20_n_0 ),
        .I4(stat[0]),
        .I5(\rgf_selc0_wb[1]_i_21_n_0 ),
        .O(\rgf_selc0_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h4044404075757575)) 
    \rgf_selc1_rn_wb[0]_i_1 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\rgf_selc1_rn_wb[0]_i_2_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_3_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_4_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_5_n_0 ),
        .O(ctl_selc1_rn));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \rgf_selc1_rn_wb[0]_i_10 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [0]),
        .O(\rgf_selc1_rn_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F2F200F2)) 
    \rgf_selc1_rn_wb[0]_i_11 
       (.I0(\rgf_selc1_rn_wb[0]_i_18_n_0 ),
        .I1(\bdatw[31]_INST_0_i_110_n_0 ),
        .I2(\badr[15]_INST_0_i_51_n_0 ),
        .I3(\fch/ir1 [8]),
        .I4(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFBEFFFF)) 
    \rgf_selc1_rn_wb[0]_i_12 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [3]),
        .I3(\rgf_selc1_rn_wb[1]_i_14_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_20_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8A888A888A88AAAA)) 
    \rgf_selc1_rn_wb[0]_i_13 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_21_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_22_n_0 ),
        .I3(\rgf_selc1_rn_wb[0]_i_23_n_0 ),
        .I4(\rgf_selc1_rn_wb[0]_i_24_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_25_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_14 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_15 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h440F000000000000)) 
    \rgf_selc1_rn_wb[0]_i_16 
       (.I0(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_26_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [0]),
        .O(\rgf_selc1_rn_wb[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00F7FFF7FFF7FFF7)) 
    \rgf_selc1_rn_wb[0]_i_17 
       (.I0(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [0]),
        .I5(\rgf_selc1_rn_wb[2]_i_25_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAFEAAFEAAAA)) 
    \rgf_selc1_rn_wb[0]_i_18 
       (.I0(\rgf_selc1_wb[1]_i_38_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_28_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\rgf_selc1_rn_wb[0]_i_29_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_30_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h88884444CC0C00C0)) 
    \rgf_selc1_rn_wb[0]_i_19 
       (.I0(\rgf_selc1_rn_wb[0]_i_31_n_0 ),
        .I1(\bdatw[31]_INST_0_i_44_n_0 ),
        .I2(\fch/ir1 [12]),
        .I3(\rgf/sreg/sr [4]),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [13]),
        .O(\rgf_selc1_rn_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \rgf_selc1_rn_wb[0]_i_2 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\niss_dsp_b1[1]_INST_0_i_8_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \rgf_selc1_rn_wb[0]_i_20 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [4]),
        .O(\rgf_selc1_rn_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \rgf_selc1_rn_wb[0]_i_21 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [6]),
        .O(\rgf_selc1_rn_wb[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h33FFF7FFFFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_22 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [10]),
        .I2(\rgf_selc1_rn_wb[1]_i_23_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[0]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0E0AFFFF)) 
    \rgf_selc1_rn_wb[0]_i_23 
       (.I0(\rgf_selc1_rn_wb[0]_i_33_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_34_n_0 ),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [9]),
        .I5(\rgf_selc1_rn_wb[0]_i_35_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hF500FD00FF000000)) 
    \rgf_selc1_rn_wb[0]_i_24 
       (.I0(\rgf_selc1_rn_wb[0]_i_27_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF0075FFFF7777)) 
    \rgf_selc1_rn_wb[0]_i_25 
       (.I0(\fch/ir1 [3]),
        .I1(div_crdy1),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [11]),
        .I5(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_25_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_26 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[0]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[0]_i_27 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [3]),
        .O(\rgf_selc1_rn_wb[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF3FFFEEFF)) 
    \rgf_selc1_rn_wb[0]_i_28 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [7]),
        .I5(dctl_sign_f_i_4_n_0),
        .O(\rgf_selc1_rn_wb[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00004400C400CC00)) 
    \rgf_selc1_rn_wb[0]_i_29 
       (.I0(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hA2AAAAAAA2AAA2AA)) 
    \rgf_selc1_rn_wb[0]_i_3 
       (.I0(\rgf_selc1_rn_wb[0]_i_8_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_9_n_0 ),
        .I2(\rgf_selc1_rn_wb[0]_i_10_n_0 ),
        .I3(\niss_dsp_b1[0]_INST_0_i_8_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\fch/ir1 [1]),
        .O(\rgf_selc1_rn_wb[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF5F5DFF75FFCFFFD)) 
    \rgf_selc1_rn_wb[0]_i_30 
       (.I0(\fch/ir1 [0]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [6]),
        .O(\rgf_selc1_rn_wb[0]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'hCA)) 
    \rgf_selc1_rn_wb[0]_i_31 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [12]),
        .O(\rgf_selc1_rn_wb[0]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_rn_wb[0]_i_32 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[0]_i_32_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[0]_i_33 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .O(\rgf_selc1_rn_wb[0]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h7777FF7F)) 
    \rgf_selc1_rn_wb[0]_i_34 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [5]),
        .O(\rgf_selc1_rn_wb[0]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \rgf_selc1_rn_wb[0]_i_35 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [4]),
        .O(\rgf_selc1_rn_wb[0]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_rn_wb[0]_i_4 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .O(\rgf_selc1_rn_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h000000000D000D0D)) 
    \rgf_selc1_rn_wb[0]_i_5 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_11_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\rgf_selc1_rn_wb[0]_i_12_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\rgf_selc1_rn_wb[0]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \rgf_selc1_rn_wb[0]_i_6 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [5]),
        .O(\rgf_selc1_rn_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \rgf_selc1_rn_wb[0]_i_7 
       (.I0(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_15_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [14]),
        .O(\rgf_selc1_rn_wb[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h55554155FFFFFFFF)) 
    \rgf_selc1_rn_wb[0]_i_8 
       (.I0(\rgf_selc1_rn_wb[0]_i_16_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [10]),
        .I4(\rgf_selc1_rn_wb[0]_i_17_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_4_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \rgf_selc1_rn_wb[0]_i_9 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [14]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [9]),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h1055101055555555)) 
    \rgf_selc1_rn_wb[1]_i_1 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\rgf_selc1_rn_wb[1]_i_2_n_0 ),
        .I2(\bcmd[2]_INST_0_i_5_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_3_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_5_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[1]_i_10 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [1]),
        .O(\rgf_selc1_rn_wb[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAABAAAAAA)) 
    \rgf_selc1_rn_wb[1]_i_11 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [10]),
        .I5(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[1]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \rgf_selc1_rn_wb[1]_i_12 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[1]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \rgf_selc1_rn_wb[1]_i_13 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [4]),
        .O(\rgf_selc1_rn_wb[1]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_selc1_rn_wb[1]_i_14 
       (.I0(\fch/ir1 [15]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .O(\rgf_selc1_rn_wb[1]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_15 
       (.I0(brdy),
        .I1(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    \rgf_selc1_rn_wb[1]_i_16 
       (.I0(\fch/ir1 [6]),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_19_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_20_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_21_n_0 ),
        .I5(\bcmd[1]_INST_0_i_21_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5DDDDDD)) 
    \rgf_selc1_rn_wb[1]_i_17 
       (.I0(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_22_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_23_n_0 ),
        .I3(\fch/ir1 [4]),
        .I4(\rgf_selc1_rn_wb[1]_i_24_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_25_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0EFE0EFE0EFE0)) 
    \rgf_selc1_rn_wb[1]_i_18 
       (.I0(\rgf_selc1_rn_wb[1]_i_26_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_27_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\rgf_selc1_rn_wb[1]_i_28_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[1]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc1_rn_wb[1]_i_19 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [2]),
        .O(\rgf_selc1_rn_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hD0D0D0DDDDDDD0DD)) 
    \rgf_selc1_rn_wb[1]_i_2 
       (.I0(\fch/ir1 [9]),
        .I1(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_6_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_7_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\rgf_selc1_rn_wb[1]_i_8_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[1]_i_20 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[1]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc1_rn_wb[1]_i_21 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [13]),
        .O(\rgf_selc1_rn_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFFFFFFFFFF)) 
    \rgf_selc1_rn_wb[1]_i_22 
       (.I0(\fch/ir1 [3]),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\bdatw[31]_INST_0_i_151_n_0 ),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [8]),
        .I5(ctl_fetch1_fl_i_30_n_0),
        .O(\rgf_selc1_rn_wb[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_23 
       (.I0(\fch/ir1 [7]),
        .I1(div_crdy1),
        .O(\rgf_selc1_rn_wb[1]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_24 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[1]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF040404)) 
    \rgf_selc1_rn_wb[1]_i_25 
       (.I0(\rgf_selc1_rn_wb[1]_i_29_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_30_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_5_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_31_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0280000200000000)) 
    \rgf_selc1_rn_wb[1]_i_26 
       (.I0(\bcmd[2]_INST_0_i_2_n_0 ),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [1]),
        .O(\rgf_selc1_rn_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0808800000000000)) 
    \rgf_selc1_rn_wb[1]_i_27 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [1]),
        .O(\rgf_selc1_rn_wb[1]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[1]_i_28 
       (.I0(\fch/ir1 [4]),
        .I1(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[1]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \rgf_selc1_rn_wb[1]_i_29 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [4]),
        .O(\rgf_selc1_rn_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h0000007500770077)) 
    \rgf_selc1_rn_wb[1]_i_3 
       (.I0(\rgf_selc1_rn_wb[1]_i_9_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_10_n_0 ),
        .I2(\fch/ir1 [9]),
        .I3(\rgf_selc1_rn_wb[1]_i_11_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_12_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \rgf_selc1_rn_wb[1]_i_30 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [10]),
        .I2(div_crdy1),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[1]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0000570000000000)) 
    \rgf_selc1_rn_wb[1]_i_31 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(dctl_sign_f_i_4_n_0),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [11]),
        .I5(div_crdy1),
        .O(\rgf_selc1_rn_wb[1]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h0400000000000000)) 
    \rgf_selc1_rn_wb[1]_i_4 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [13]),
        .O(\rgf_selc1_rn_wb[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAFEAAAAAAFEAAFE)) 
    \rgf_selc1_rn_wb[1]_i_5 
       (.I0(\rgf_selc1_rn_wb[1]_i_14_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_16_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_17_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_4_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \rgf_selc1_rn_wb[1]_i_6 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [15]),
        .O(\rgf_selc1_rn_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h5000010000000100)) 
    \rgf_selc1_rn_wb[1]_i_7 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [6]),
        .O(\rgf_selc1_rn_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88B888B888B8B8B8)) 
    \rgf_selc1_rn_wb[1]_i_8 
       (.I0(\rgf_selc1_rn_wb[1]_i_18_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0088808800880088)) 
    \rgf_selc1_rn_wb[1]_i_9 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .I5(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .O(\rgf_selc1_rn_wb[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5455545444444444)) 
    \rgf_selc1_rn_wb[2]_i_1 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\rgf_selc1_rn_wb[2]_i_2_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_3_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I4(\fch/ir1 [10]),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0B000000)) 
    \rgf_selc1_rn_wb[2]_i_10 
       (.I0(\bcmd[1]_INST_0_i_26_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [10]),
        .I4(\rgf_selc1_rn_wb[2]_i_23_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_24_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \rgf_selc1_rn_wb[2]_i_11 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFF5577FFF7DFFFFD)) 
    \rgf_selc1_rn_wb[2]_i_12 
       (.I0(\fch/ir1 [2]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \rgf_selc1_rn_wb[2]_i_13 
       (.I0(\rgf_selc1_rn_wb[0]_i_7_n_0 ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [2]),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_selc1_rn_wb[2]_i_14 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF0F0000080008000)) 
    \rgf_selc1_rn_wb[2]_i_15 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_25_n_0 ),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[2]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_rn_wb[2]_i_16 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[2]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_rn_wb[2]_i_17 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [4]),
        .O(\rgf_selc1_rn_wb[2]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \rgf_selc1_rn_wb[2]_i_18 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .O(\rgf_selc1_rn_wb[2]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[2]_i_19 
       (.I0(div_crdy1),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hF200FFFFF200F200)) 
    \rgf_selc1_rn_wb[2]_i_2 
       (.I0(\rgf_selc1_rn_wb[2]_i_5_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_7_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_8_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h55455555FFFFFFFF)) 
    \rgf_selc1_rn_wb[2]_i_20 
       (.I0(\rgf_selc1_rn_wb[2]_i_26_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [5]),
        .I3(\rgf_selc1_rn_wb[1]_i_23_n_0 ),
        .I4(\fch/ir1 [8]),
        .I5(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h004400000F440000)) 
    \rgf_selc1_rn_wb[2]_i_21 
       (.I0(\fch/ir1 [11]),
        .I1(div_crdy1),
        .I2(\rgf_selc1_rn_wb[2]_i_27_n_0 ),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[2]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hF2FF3FFF)) 
    \rgf_selc1_rn_wb[2]_i_22 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [10]),
        .O(\rgf_selc1_rn_wb[2]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA0000300)) 
    \rgf_selc1_rn_wb[2]_i_23 
       (.I0(\fch/ir1 [6]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [8]),
        .I5(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[2]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h44444C44FC44FC44)) 
    \rgf_selc1_rn_wb[2]_i_24 
       (.I0(\rgf_selc1_rn_wb[2]_i_28_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [7]),
        .I3(\rgf_selc1_rn_wb[2]_i_25_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[2]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \rgf_selc1_rn_wb[2]_i_25 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[2]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \rgf_selc1_rn_wb[2]_i_26 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\bdatw[31]_INST_0_i_151_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [2]),
        .I5(ctl_fetch1_fl_i_30_n_0),
        .O(\rgf_selc1_rn_wb[2]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFF4)) 
    \rgf_selc1_rn_wb[2]_i_27 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[2]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFDFDFDDD)) 
    \rgf_selc1_rn_wb[2]_i_28 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [8]),
        .O(\rgf_selc1_rn_wb[2]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h4040404455555555)) 
    \rgf_selc1_rn_wb[2]_i_3 
       (.I0(\fch/ir1 [15]),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_10_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_11_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_12_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_13_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \rgf_selc1_rn_wb[2]_i_4 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [12]),
        .O(\rgf_selc1_rn_wb[2]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_rn_wb[2]_i_5 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .O(\rgf_selc1_rn_wb[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFBFFFBFFF00FFBF)) 
    \rgf_selc1_rn_wb[2]_i_6 
       (.I0(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I1(\fch/ir1 [5]),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [2]),
        .I5(\fch/ir1 [9]),
        .O(\rgf_selc1_rn_wb[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAEAAA)) 
    \rgf_selc1_rn_wb[2]_i_7 
       (.I0(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_18_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .O(\rgf_selc1_rn_wb[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h2222220222222222)) 
    \rgf_selc1_rn_wb[2]_i_8 
       (.I0(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .I2(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [5]),
        .O(\rgf_selc1_rn_wb[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000800000)) 
    \rgf_selc1_rn_wb[2]_i_9 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [14]),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\fch/ir1 [15]),
        .O(\rgf_selc1_rn_wb[2]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    rgf_selc1_stat_i_1
       (.I0(ctl_selc1[1]),
        .I1(ctl_selc1[0]),
        .O(rgf_selc1_stat_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rgf_selc1_stat_i_2
       (.I0(fch_wrbufn1),
        .O(rgf_selc1_stat_i_2_n_0));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAFEAAAA)) 
    \rgf_selc1_wb[0]_i_1 
       (.I0(\rgf_selc1_wb[0]_i_2_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\rgf_selc1_wb[0]_i_3_n_0 ),
        .I3(\bcmd[3]_INST_0_i_4_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_5_n_0 ),
        .O(ctl_selc1[0]));
  LUT6 #(
    .INIT(64'hFFFFEFEEEFEFCFCF)) 
    \rgf_selc1_wb[0]_i_10 
       (.I0(\fch/ir1 [9]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [11]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [10]),
        .O(\rgf_selc1_wb[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h70FF50FFFFFF50FF)) 
    \rgf_selc1_wb[0]_i_11 
       (.I0(\bcmd[3]_INST_0_i_13_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_16_n_0 ),
        .I2(\fch/ir1 [10]),
        .I3(\rgf_selc1_wb[0]_i_17_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_18_n_0 ),
        .O(\rgf_selc1_wb[0]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h8080BF80B0B0BFBF)) 
    \rgf_selc1_wb[0]_i_12 
       (.I0(\rgf_selc1_wb[0]_i_19_n_0 ),
        .I1(\fch/ir1 [9]),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\fch/ir1 [7]),
        .I4(div_crdy1),
        .I5(\rgf_selc1_wb[1]_i_31_n_0 ),
        .O(\rgf_selc1_wb[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF0C0400FFFFFFFF)) 
    \rgf_selc1_wb[0]_i_13 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [5]),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [4]),
        .O(\rgf_selc1_wb[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFC000000FCFFF9FE)) 
    \rgf_selc1_wb[0]_i_14 
       (.I0(\fch/ir1 [3]),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [4]),
        .O(\rgf_selc1_wb[0]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFBBFFAAFFBBF0)) 
    \rgf_selc1_wb[0]_i_15 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I2(ctl_fetch1_fl_i_13_n_0),
        .I3(\fch/ir1 [11]),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\rgf_selc1_wb[0]_i_20_n_0 ),
        .O(\rgf_selc1_wb[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFCFFFFF7FFFFFFF)) 
    \rgf_selc1_wb[0]_i_16 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [4]),
        .O(\rgf_selc1_wb[0]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \rgf_selc1_wb[0]_i_17 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .I2(div_crdy1),
        .O(\rgf_selc1_wb[0]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \rgf_selc1_wb[0]_i_18 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [10]),
        .O(\rgf_selc1_wb[0]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFF5DFFFF)) 
    \rgf_selc1_wb[0]_i_19 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\rgf_selc1_wb[0]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h6D77000000000000)) 
    \rgf_selc1_wb[0]_i_2 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [15]),
        .I5(\rgf_selc1_wb[0]_i_6_n_0 ),
        .O(\rgf_selc1_wb[0]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \rgf_selc1_wb[0]_i_20 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h8888B888BBBBBBBB)) 
    \rgf_selc1_wb[0]_i_3 
       (.I0(\rgf_selc1_wb[0]_i_7_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_8_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\fch/ir1 [10]),
        .I4(\rgf_selc1_wb[0]_i_9_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_10_n_0 ),
        .O(\rgf_selc1_wb[0]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \rgf_selc1_wb[0]_i_4 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [12]),
        .O(\rgf_selc1_wb[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF0F070F0F0F07000)) 
    \rgf_selc1_wb[0]_i_5 
       (.I0(\fch/ir1 [8]),
        .I1(\rgf_selc1_wb[0]_i_11_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [11]),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\rgf_selc1_wb[0]_i_12_n_0 ),
        .O(\rgf_selc1_wb[0]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \rgf_selc1_wb[0]_i_6 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .O(\rgf_selc1_wb[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00008000FFFFFFFF)) 
    \rgf_selc1_wb[0]_i_7 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [10]),
        .I3(\rgf_selc1_wb[0]_i_13_n_0 ),
        .I4(\rgf_selc1_wb[0]_i_14_n_0 ),
        .I5(\rgf_selc1_wb[0]_i_15_n_0 ),
        .O(\rgf_selc1_wb[0]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hF000FB00)) 
    \rgf_selc1_wb[0]_i_8 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [10]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFBFFFBFFA2AAFFFF)) 
    \rgf_selc1_wb[0]_i_9 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\bcmd[2]_INST_0_i_6_n_0 ),
        .I5(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FDDD)) 
    \rgf_selc1_wb[1]_i_1 
       (.I0(\rgf_selc1_wb[1]_i_2_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_3_n_0 ),
        .I2(\rgf_selc1_wb_reg[1]_i_4_n_0 ),
        .I3(\rgf_selc1_wb[1]_i_5_n_0 ),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\rgf_selc1_wb[1]_i_6_n_0 ),
        .O(ctl_selc1[1]));
  LUT6 #(
    .INIT(64'h0000000000002A8A)) 
    \rgf_selc1_wb[1]_i_10 
       (.I0(\fch/ir1 [15]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [14]),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\rgf_selc1_wb[1]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_11 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [15]),
        .O(\rgf_selc1_wb[1]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0101010101000000)) 
    \rgf_selc1_wb[1]_i_12 
       (.I0(\rgf_selc1_wb[1]_i_28_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\bcmd[1]_INST_0_i_16_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I5(\fch/ir1 [8]),
        .O(\rgf_selc1_wb[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h2000202020002000)) 
    \rgf_selc1_wb[1]_i_13 
       (.I0(\fch/ir1 [12]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(ctl_fetch1_fl_i_16_n_0),
        .I3(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_30_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_31_n_0 ),
        .O(\rgf_selc1_wb[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000203030)) 
    \rgf_selc1_wb[1]_i_14 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_32_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\fch/ir1 [1]),
        .I5(\fch/ir1 [9]),
        .O(\rgf_selc1_wb[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hABBBABBBABBBAABA)) 
    \rgf_selc1_wb[1]_i_15 
       (.I0(\rgf_selc1_wb[1]_i_34_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\fch/ir1 [12]),
        .I3(\rgf_selc1_wb[1]_i_35_n_0 ),
        .I4(\bdatw[31]_INST_0_i_116_n_0 ),
        .I5(\fch/ir1 [15]),
        .O(\rgf_selc1_wb[1]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000047)) 
    \rgf_selc1_wb[1]_i_16 
       (.I0(\rgf_selc1_wb[0]_i_12_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_36_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_37_n_0 ),
        .I3(\fch/ir1 [15]),
        .I4(\rgf_selc1_wb[1]_i_38_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_39_n_0 ),
        .O(\rgf_selc1_wb[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \rgf_selc1_wb[1]_i_17 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [9]),
        .I2(\bdatw[31]_INST_0_i_44_n_0 ),
        .I3(\fch/ir1 [12]),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\rgf_selc1_rn_wb[0]_i_14_n_0 ),
        .O(\rgf_selc1_wb[1]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \rgf_selc1_wb[1]_i_18 
       (.I0(\fch/ir1 [1]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [13]),
        .O(\rgf_selc1_wb[1]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \rgf_selc1_wb[1]_i_19 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [4]),
        .O(\rgf_selc1_wb[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF7F00)) 
    \rgf_selc1_wb[1]_i_2 
       (.I0(\rgf_selc1_wb[1]_i_7_n_0 ),
        .I1(\rgf_selc1_wb[0]_i_4_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\rgf_selc1_wb[1]_i_8_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_9_n_0 ),
        .O(\rgf_selc1_wb[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4FCF5FFFDFDFF3FF)) 
    \rgf_selc1_wb[1]_i_20 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [5]),
        .O(\rgf_selc1_wb[1]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \rgf_selc1_wb[1]_i_21 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hF7F7F7F7FF7FF7FF)) 
    \rgf_selc1_wb[1]_i_22 
       (.I0(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I1(\bdatw[31]_INST_0_i_151_n_0 ),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \rgf_selc1_wb[1]_i_23 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [8]),
        .O(\rgf_selc1_wb[1]_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[1]_i_24 
       (.I0(\fch/ir1 [7]),
        .I1(\rgf/sreg/sr [8]),
        .O(\rgf_selc1_wb[1]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hFF01FFFF)) 
    \rgf_selc1_wb[1]_i_25 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [10]),
        .I2(\fch/ir1 [7]),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\rgf_selc1_wb[0]_i_4_n_0 ),
        .O(\rgf_selc1_wb[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0404000400000004)) 
    \rgf_selc1_wb[1]_i_26 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [8]),
        .I2(\stat[1]_i_22_n_0 ),
        .I3(\fch/ir1 [3]),
        .I4(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I5(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFABAFABAAAAAFAA)) 
    \rgf_selc1_wb[1]_i_27 
       (.I0(\rgf_selc1_wb[1]_i_40_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [14]),
        .I4(\rgf/sreg/sr [5]),
        .I5(\fch/ir1 [13]),
        .O(\rgf_selc1_wb[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFE0000FFFF0000)) 
    \rgf_selc1_wb[1]_i_28 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [5]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[1]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_29 
       (.I0(\fch/ir1 [7]),
        .I1(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[1]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hEEAEEEAEEEAEEAAA)) 
    \rgf_selc1_wb[1]_i_3 
       (.I0(\rgf_selc1_wb[1]_i_10_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_11_n_0 ),
        .I2(\fch/ir1 [11]),
        .I3(\rgf_selc1_wb[1]_i_12_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_13_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_14_n_0 ),
        .O(\rgf_selc1_wb[1]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hA2AA)) 
    \rgf_selc1_wb[1]_i_30 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\rgf_selc1_wb[1]_i_30_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rgf_selc1_wb[1]_i_31 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [8]),
        .O(\rgf_selc1_wb[1]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \rgf_selc1_wb[1]_i_32 
       (.I0(\bcmd[1]_INST_0_i_25_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [8]),
        .O(\rgf_selc1_wb[1]_i_32_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \rgf_selc1_wb[1]_i_33 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [6]),
        .O(\rgf_selc1_wb[1]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080A0B300)) 
    \rgf_selc1_wb[1]_i_34 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .I5(\rgf_selc1_wb[1]_i_41_n_0 ),
        .O(\rgf_selc1_wb[1]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \rgf_selc1_wb[1]_i_35 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\fch/ir1 [13]),
        .I2(\rgf/sreg/sr [4]),
        .O(\rgf_selc1_wb[1]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'hFFEFAAAAAAAAAAAA)) 
    \rgf_selc1_wb[1]_i_36 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [10]),
        .I5(\rgf_selc1_wb[1]_i_42_n_0 ),
        .O(\rgf_selc1_wb[1]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hF57FFFFF)) 
    \rgf_selc1_wb[1]_i_37 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .O(\rgf_selc1_wb[1]_i_37_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \rgf_selc1_wb[1]_i_38 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [13]),
        .O(\rgf_selc1_wb[1]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h10010101)) 
    \rgf_selc1_wb[1]_i_39 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [13]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir1 [12]),
        .I4(\rgf/sreg/sr [7]),
        .O(\rgf_selc1_wb[1]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \rgf_selc1_wb[1]_i_40 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [15]),
        .I2(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[1]_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \rgf_selc1_wb[1]_i_41 
       (.I0(\niss_dsp_a1[32]_INST_0_i_26_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [12]),
        .I4(\fch/ir1 [13]),
        .O(\rgf_selc1_wb[1]_i_41_n_0 ));
  LUT5 #(
    .INIT(32'h14001403)) 
    \rgf_selc1_wb[1]_i_42 
       (.I0(\bcmd[2]_INST_0_i_6_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [7]),
        .I4(\rgf/sreg/sr [8]),
        .O(\rgf_selc1_wb[1]_i_42_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \rgf_selc1_wb[1]_i_5 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\fch/ir1 [11]),
        .O(\rgf_selc1_wb[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020000000)) 
    \rgf_selc1_wb[1]_i_6 
       (.I0(\rgf_selc1_wb[1]_i_17_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_18_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [0]),
        .I4(\niss_dsp_b1[0]_INST_0_i_8_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_19_n_0 ),
        .O(\rgf_selc1_wb[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF4F0F4F0F4F0FFF0)) 
    \rgf_selc1_wb[1]_i_7 
       (.I0(\rgf_selc1_wb[1]_i_20_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\rgf_selc1_wb[1]_i_21_n_0 ),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [9]),
        .I5(\rgf_selc1_rn_wb[1]_i_23_n_0 ),
        .O(\rgf_selc1_wb[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000AA08)) 
    \rgf_selc1_wb[1]_i_8 
       (.I0(\rgf_selc1_wb[1]_i_22_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I2(\rgf_selc1_wb[1]_i_24_n_0 ),
        .I3(\fch/ir1 [9]),
        .I4(\rgf_selc1_wb[1]_i_25_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_26_n_0 ),
        .O(\rgf_selc1_wb[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF213F0000)) 
    \rgf_selc1_wb[1]_i_9 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir1 [13]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir1 [14]),
        .I4(\stat[2]_i_9_n_0 ),
        .I5(\rgf_selc1_wb[1]_i_27_n_0 ),
        .O(\rgf_selc1_wb[1]_i_9_n_0 ));
  MUXF7 \rgf_selc1_wb_reg[1]_i_4 
       (.I0(\rgf_selc1_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_16_n_0 ),
        .O(\rgf_selc1_wb_reg[1]_i_4_n_0 ),
        .S(\fch/ir1 [14]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[0]_i_1 
       (.I0(\sp[0]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [0]),
        .I4(\rgf/rgf_c1bus_0 [0]),
        .O(\sp[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \sp[0]_i_2 
       (.I0(\rgf/sptr/sp [0]),
        .I1(\sp[31]_i_8_n_0 ),
        .I2(\rgf/sptr/data2 [0]),
        .O(\sp[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[10]_i_1 
       (.I0(\sp[10]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [10]),
        .I4(\rgf/rgf_c1bus_0 [10]),
        .O(\sp[10]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[10]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [10]),
        .I2(\rgf/sptr/sp [10]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [10]),
        .O(\sp[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[11]_i_1 
       (.I0(\sp[11]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [11]),
        .I4(\rgf/rgf_c1bus_0 [11]),
        .O(\sp[11]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[11]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [11]),
        .I2(\rgf/sptr/sp [11]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [11]),
        .O(\sp[11]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[12]_i_1 
       (.I0(\sp[12]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [12]),
        .I4(\rgf/rgf_c1bus_0 [12]),
        .O(\sp[12]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[12]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [12]),
        .I2(\rgf/sptr/sp [12]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [12]),
        .O(\sp[12]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[13]_i_1 
       (.I0(\sp[13]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [13]),
        .I4(\rgf/rgf_c1bus_0 [13]),
        .O(\sp[13]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[13]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [13]),
        .I2(\rgf/sptr/sp [13]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [13]),
        .O(\sp[13]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[14]_i_1 
       (.I0(\sp[14]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [14]),
        .I4(\rgf/rgf_c1bus_0 [14]),
        .O(\sp[14]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[14]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [14]),
        .I2(\rgf/sptr/sp [14]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [14]),
        .O(\sp[14]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[15]_i_1 
       (.I0(\sp[15]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [15]),
        .I4(\rgf/rgf_c1bus_0 [15]),
        .O(\sp[15]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[15]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [15]),
        .I2(\rgf/sptr/sp [15]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [15]),
        .O(\sp[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[16]_i_1 
       (.I0(\sp[16]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [16]),
        .I4(\rgf/rgf_c1bus_0 [16]),
        .O(\sp[16]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[16]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [16]),
        .I2(\rgf/sptr/sp [16]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [16]),
        .O(\sp[16]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[16]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[16]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [16]),
        .O(\rgf/rgf_c0bus_0 [16]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[16]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[16]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [16]),
        .O(\rgf/rgf_c1bus_0 [16]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[17]_i_1 
       (.I0(\sp[17]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [17]),
        .I4(\rgf/rgf_c1bus_0 [17]),
        .O(\sp[17]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[17]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [17]),
        .I2(\rgf/sptr/sp [17]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [17]),
        .O(\sp[17]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[17]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[17]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [17]),
        .O(\rgf/rgf_c0bus_0 [17]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[17]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[17]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [17]),
        .O(\rgf/rgf_c1bus_0 [17]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[18]_i_1 
       (.I0(\sp[18]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [18]),
        .I4(\rgf/rgf_c1bus_0 [18]),
        .O(\sp[18]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[18]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [18]),
        .I2(\rgf/sptr/sp [18]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [18]),
        .O(\sp[18]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[18]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[18]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [18]),
        .O(\rgf/rgf_c0bus_0 [18]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[18]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[18]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [18]),
        .O(\rgf/rgf_c1bus_0 [18]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[19]_i_1 
       (.I0(\sp[19]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [19]),
        .I4(\rgf/rgf_c1bus_0 [19]),
        .O(\sp[19]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[19]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [19]),
        .I2(\rgf/sptr/sp [19]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [19]),
        .O(\sp[19]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[19]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[19]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [19]),
        .O(\rgf/rgf_c0bus_0 [19]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[19]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[19]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [19]),
        .O(\rgf/rgf_c1bus_0 [19]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[1]_i_1 
       (.I0(\sp[1]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [1]),
        .I4(\rgf/rgf_c1bus_0 [1]),
        .O(\sp[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[1]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [1]),
        .I2(\rgf/sptr/sp [1]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [1]),
        .O(\sp[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[20]_i_1 
       (.I0(\sp[20]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [20]),
        .I4(\rgf/rgf_c1bus_0 [20]),
        .O(\sp[20]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[20]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [20]),
        .I2(\rgf/sptr/sp [20]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [20]),
        .O(\sp[20]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[20]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[20]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [20]),
        .O(\rgf/rgf_c0bus_0 [20]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[20]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[20]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [20]),
        .O(\rgf/rgf_c1bus_0 [20]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[21]_i_1 
       (.I0(\sp[21]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [21]),
        .I4(\rgf/rgf_c1bus_0 [21]),
        .O(\sp[21]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[21]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [21]),
        .I2(\rgf/sptr/sp [21]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [21]),
        .O(\sp[21]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[21]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[21]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [21]),
        .O(\rgf/rgf_c0bus_0 [21]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[21]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[21]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [21]),
        .O(\rgf/rgf_c1bus_0 [21]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[22]_i_1 
       (.I0(\sp[22]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [22]),
        .I4(\rgf/rgf_c1bus_0 [22]),
        .O(\sp[22]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[22]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [22]),
        .I2(\rgf/sptr/sp [22]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [22]),
        .O(\sp[22]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[22]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[22]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [22]),
        .O(\rgf/rgf_c0bus_0 [22]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[22]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[22]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [22]),
        .O(\rgf/rgf_c1bus_0 [22]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[23]_i_1 
       (.I0(\sp[23]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [23]),
        .I4(\rgf/rgf_c1bus_0 [23]),
        .O(\sp[23]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[23]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [23]),
        .I2(\rgf/sptr/sp [23]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [23]),
        .O(\sp[23]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[23]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[23]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [23]),
        .O(\rgf/rgf_c0bus_0 [23]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[23]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[23]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [23]),
        .O(\rgf/rgf_c1bus_0 [23]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[24]_i_1 
       (.I0(\sp[24]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [24]),
        .I4(\rgf/rgf_c1bus_0 [24]),
        .O(\sp[24]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[24]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [24]),
        .I2(\rgf/sptr/sp [24]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [24]),
        .O(\sp[24]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[24]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[24]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [24]),
        .O(\rgf/rgf_c0bus_0 [24]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[24]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[24]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [24]),
        .O(\rgf/rgf_c1bus_0 [24]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[25]_i_1 
       (.I0(\sp[25]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [25]),
        .I4(\rgf/rgf_c1bus_0 [25]),
        .O(\sp[25]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[25]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [25]),
        .I2(\rgf/sptr/sp [25]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [25]),
        .O(\sp[25]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[25]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[25]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [25]),
        .O(\rgf/rgf_c0bus_0 [25]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[25]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[25]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [25]),
        .O(\rgf/rgf_c1bus_0 [25]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[26]_i_1 
       (.I0(\sp[26]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [26]),
        .I4(\rgf/rgf_c1bus_0 [26]),
        .O(\sp[26]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[26]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [26]),
        .I2(\rgf/sptr/sp [26]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [26]),
        .O(\sp[26]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[26]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[26]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [26]),
        .O(\rgf/rgf_c0bus_0 [26]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[26]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[26]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [26]),
        .O(\rgf/rgf_c1bus_0 [26]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[27]_i_1 
       (.I0(\sp[27]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [27]),
        .I4(\rgf/rgf_c1bus_0 [27]),
        .O(\sp[27]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[27]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [27]),
        .I2(\rgf/sptr/sp [27]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [27]),
        .O(\sp[27]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[27]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[27]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [27]),
        .O(\rgf/rgf_c0bus_0 [27]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[27]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[27]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [27]),
        .O(\rgf/rgf_c1bus_0 [27]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[28]_i_1 
       (.I0(\sp[28]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [28]),
        .I4(\rgf/rgf_c1bus_0 [28]),
        .O(\sp[28]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[28]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [28]),
        .I2(\rgf/sptr/sp [28]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [28]),
        .O(\sp[28]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[28]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[28]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [28]),
        .O(\rgf/rgf_c0bus_0 [28]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[28]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[28]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [28]),
        .O(\rgf/rgf_c1bus_0 [28]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[29]_i_1 
       (.I0(\sp[29]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [29]),
        .I4(\rgf/rgf_c1bus_0 [29]),
        .O(\sp[29]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[29]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [29]),
        .I2(\rgf/sptr/sp [29]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [29]),
        .O(\sp[29]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[29]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[29]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [29]),
        .O(\rgf/rgf_c0bus_0 [29]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[29]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[29]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [29]),
        .O(\rgf/rgf_c1bus_0 [29]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[2]_i_1 
       (.I0(\sp[2]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [2]),
        .I4(\rgf/rgf_c1bus_0 [2]),
        .O(\sp[2]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[2]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [2]),
        .I2(\rgf/sptr/sp [2]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [2]),
        .O(\sp[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[30]_i_1 
       (.I0(\sp[30]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [30]),
        .I4(\rgf/rgf_c1bus_0 [30]),
        .O(\sp[30]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[30]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [30]),
        .I2(\rgf/sptr/sp [30]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [30]),
        .O(\sp[30]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[30]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[30]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [30]),
        .O(\rgf/rgf_c0bus_0 [30]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[30]_i_4 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[30]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [30]),
        .O(\rgf/rgf_c1bus_0 [30]));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[31]_i_1 
       (.I0(\sp[31]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [31]),
        .I4(\rgf/rgf_c1bus_0 [31]),
        .O(\sp[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEEFFFF89)) 
    \sp[31]_i_10 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(fch_irq_req),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [12]),
        .I5(\sp[31]_i_18_n_0 ),
        .O(\sp[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFE5F)) 
    \sp[31]_i_11 
       (.I0(stat[1]),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [1]),
        .I5(\fch/ir0 [2]),
        .O(\sp[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h2204920022009200)) 
    \sp[31]_i_12 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [8]),
        .O(\sp[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFF45000000000000)) 
    \sp[31]_i_13 
       (.I0(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I1(\sp[31]_i_19_n_0 ),
        .I2(\sp[31]_i_20_n_0 ),
        .I3(\sp[31]_i_21_n_0 ),
        .I4(\sp[31]_i_22_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(ctl_sp_dec1));
  LUT6 #(
    .INIT(64'h0000000020000002)) 
    \sp[31]_i_14 
       (.I0(\sp_reg[31]_i_23_n_0 ),
        .I1(\sp[31]_i_24_n_0 ),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [13]),
        .I5(\bcmd[0]_INST_0_i_17_n_0 ),
        .O(ctl_sp_inc0));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sp[31]_i_15 
       (.I0(\bcmd[0]_INST_0_i_3_n_0 ),
        .I1(\fch/ir1 [15]),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .O(\sp[31]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7FFFFFFD)) 
    \sp[31]_i_16 
       (.I0(brdy),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [14]),
        .I5(\sp[31]_i_25_n_0 ),
        .O(\sp[31]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0002000200000002)) 
    \sp[31]_i_17 
       (.I0(\bcmd[0]_INST_0_i_18_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [5]),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [7]),
        .O(\sp[31]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF5FFFEFFF)) 
    \sp[31]_i_18 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [6]),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(brdy),
        .I4(\fch/ir0 [9]),
        .I5(\sp[31]_i_26_n_0 ),
        .O(\sp[31]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h2000)) 
    \sp[31]_i_19 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [7]),
        .O(\sp[31]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[31]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [31]),
        .I2(\rgf/sptr/sp [31]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [31]),
        .O(\sp[31]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFDFFFDFFFFFFFFDF)) 
    \sp[31]_i_20 
       (.I0(\sp[31]_i_27_n_0 ),
        .I1(\bdatw[9]_INST_0_i_10_n_0 ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [8]),
        .I5(\ctl1/stat_reg_n_0_[1] ),
        .O(\sp[31]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h22009200)) 
    \sp[31]_i_21 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [7]),
        .O(\sp[31]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011000076)) 
    \sp[31]_i_22 
       (.I0(\ctl1/stat_reg_n_0_[1] ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(fch_irq_req),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [12]),
        .I5(\sp[31]_i_28_n_0 ),
        .O(\sp[31]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAFFFFFFE)) 
    \sp[31]_i_24 
       (.I0(\sp[31]_i_31_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [9]),
        .I5(\stat[0]_i_10__1_n_0 ),
        .O(\sp[31]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h7FFFFFFF7FFFFFFE)) 
    \sp[31]_i_25 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [7]),
        .O(\sp[31]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h7EFFFFFFFFFFFF7E)) 
    \sp[31]_i_26 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [10]),
        .O(\sp[31]_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \sp[31]_i_27 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .O(\sp[31]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBBFE)) 
    \sp[31]_i_28 
       (.I0(\bcmd[3]_INST_0_i_4_n_0 ),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [9]),
        .I4(\sp[31]_i_32_n_0 ),
        .I5(\bcmd[0]_INST_0_i_2_n_0 ),
        .O(\sp[31]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000007410)) 
    \sp[31]_i_29 
       (.I0(stat[0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [1]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [2]),
        .I5(\fch/ir0 [6]),
        .O(\sp[31]_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[31]_i_3 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_11_n_0 ),
        .O(\rgf/c0bus_sel_cr [2]));
  LUT6 #(
    .INIT(64'h4044444400000000)) 
    \sp[31]_i_30 
       (.I0(stat[0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [5]),
        .I5(\fch/ir0 [6]),
        .O(\sp[31]_i_30_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \sp[31]_i_31 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [9]),
        .O(\sp[31]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \sp[31]_i_32 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [10]),
        .O(\sp[31]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \sp[31]_i_4 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\rgf/c1bus_sel_cr [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[31]_i_5 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[31]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [31]),
        .O(\rgf/rgf_c0bus_0 [31]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sp[31]_i_6 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(c1bus[31]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_c1bus_wb [31]),
        .O(\rgf/rgf_c1bus_0 [31]));
  LUT6 #(
    .INIT(64'hFFFFFFFF55550010)) 
    \sp[31]_i_7 
       (.I0(\sp[31]_i_10_n_0 ),
        .I1(\sp[31]_i_11_n_0 ),
        .I2(\ccmd[2]_INST_0_i_18_n_0 ),
        .I3(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I4(\sp[31]_i_12_n_0 ),
        .I5(ctl_sp_dec1),
        .O(\sp[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hABABABABAAABAAAA)) 
    \sp[31]_i_8 
       (.I0(ctl_sp_inc0),
        .I1(\sp[31]_i_15_n_0 ),
        .I2(\sp[31]_i_16_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\bcmd[0]_INST_0_i_14_n_0 ),
        .I5(\sp[31]_i_17_n_0 ),
        .O(\sp[31]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[3]_i_1 
       (.I0(\sp[3]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [3]),
        .I4(\rgf/rgf_c1bus_0 [3]),
        .O(\sp[3]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[3]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [3]),
        .I2(\rgf/sptr/sp [3]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [3]),
        .O(\sp[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \sp[3]_i_4 
       (.I0(\rgf/sptr/sp [2]),
        .I1(\rgf/sptr/ctl_sp_id4 ),
        .O(\sp[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \sp[3]_i_5 
       (.I0(\rgf/sptr/sp [1]),
        .I1(\rgf/sptr/ctl_sp_id4 ),
        .O(\sp[3]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[4]_i_1 
       (.I0(\sp[4]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [4]),
        .I4(\rgf/rgf_c1bus_0 [4]),
        .O(\sp[4]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[4]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [4]),
        .I2(\rgf/sptr/sp [4]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [4]),
        .O(\sp[4]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[5]_i_1 
       (.I0(\sp[5]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [5]),
        .I4(\rgf/rgf_c1bus_0 [5]),
        .O(\sp[5]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[5]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [5]),
        .I2(\rgf/sptr/sp [5]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [5]),
        .O(\sp[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[6]_i_1 
       (.I0(\sp[6]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [6]),
        .I4(\rgf/rgf_c1bus_0 [6]),
        .O(\sp[6]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[6]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [6]),
        .I2(\rgf/sptr/sp [6]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [6]),
        .O(\sp[6]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[7]_i_1 
       (.I0(\sp[7]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [7]),
        .I4(\rgf/rgf_c1bus_0 [7]),
        .O(\sp[7]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[7]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [7]),
        .I2(\rgf/sptr/sp [7]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [7]),
        .O(\sp[7]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[8]_i_1 
       (.I0(\sp[8]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [8]),
        .I4(\rgf/rgf_c1bus_0 [8]),
        .O(\sp[8]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[8]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [8]),
        .I2(\rgf/sptr/sp [8]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [8]),
        .O(\sp[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFEF20E02)) 
    \sp[9]_i_1 
       (.I0(\sp[9]_i_2_n_0 ),
        .I1(\rgf/c0bus_sel_cr [2]),
        .I2(\rgf/c1bus_sel_cr [2]),
        .I3(\rgf/rgf_c0bus_0 [9]),
        .I4(\rgf/rgf_c1bus_0 [9]),
        .O(\sp[9]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'hFFD800D8)) 
    \sp[9]_i_2 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\rgf/sptr/data3 [9]),
        .I2(\rgf/sptr/sp [9]),
        .I3(\sp[31]_i_8_n_0 ),
        .I4(\rgf/sptr/data2 [9]),
        .O(\sp[9]_i_2_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [11:8]),
        .S(\rgf/sptr/sp [11:8]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_3 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_3_n_0 ,\sp_reg[15]_i_3_n_1 ,\sp_reg[15]_i_3_n_2 ,\sp_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [15:12]),
        .S(\rgf/sptr/sp [15:12]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[19]_i_5 
       (.CI(\sp_reg[15]_i_3_n_0 ),
        .CO({\sp_reg[19]_i_5_n_0 ,\sp_reg[19]_i_5_n_1 ,\sp_reg[19]_i_5_n_2 ,\sp_reg[19]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [19:16]),
        .S(\rgf/sptr/sp [19:16]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[23]_i_5 
       (.CI(\sp_reg[19]_i_5_n_0 ),
        .CO({\sp_reg[23]_i_5_n_0 ,\sp_reg[23]_i_5_n_1 ,\sp_reg[23]_i_5_n_2 ,\sp_reg[23]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [23:20]),
        .S(\rgf/sptr/sp [23:20]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[27]_i_5 
       (.CI(\sp_reg[23]_i_5_n_0 ),
        .CO({\sp_reg[27]_i_5_n_0 ,\sp_reg[27]_i_5_n_1 ,\sp_reg[27]_i_5_n_2 ,\sp_reg[27]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [27:24]),
        .S(\rgf/sptr/sp [27:24]));
  MUXF7 \sp_reg[31]_i_23 
       (.I0(\sp[31]_i_29_n_0 ),
        .I1(\sp[31]_i_30_n_0 ),
        .O(\sp_reg[31]_i_23_n_0 ),
        .S(\stat[0]_i_26_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[31]_i_9 
       (.CI(\sp_reg[27]_i_5_n_0 ),
        .CO({\sp_reg[31]_i_9_n_1 ,\sp_reg[31]_i_9_n_2 ,\sp_reg[31]_i_9_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [31:28]),
        .S(\rgf/sptr/sp [31:28]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[3]_i_3 
       (.CI(\<const0> ),
        .CO({\sp_reg[3]_i_3_n_0 ,\sp_reg[3]_i_3_n_1 ,\sp_reg[3]_i_3_n_2 ,\sp_reg[3]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rgf/sptr/sp [2:1],\<const0> }),
        .O(\rgf/sptr/data2 [3:0]),
        .S({\rgf/sptr/sp [3],\sp[3]_i_4_n_0 ,\sp[3]_i_5_n_0 ,\rgf/sptr/sp [0]}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\sp_reg[3]_i_3_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(\rgf/sptr/data2 [7:4]),
        .S(\rgf/sptr/sp [7:4]));
  LUT6 #(
    .INIT(64'h8C8C808C8C808080)) 
    \sr[0]_i_1 
       (.I0(\sr[0]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\sr[11]_i_3_n_0 ),
        .I3(\sr[11]_i_4_n_0 ),
        .I4(\rgf/sreg/sr [0]),
        .I5(\rgf/rgf_c0bus_0 [0]),
        .O(\rgf/sreg/p_0_in__0 [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[0]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/sreg/sr [0]),
        .O(\sr[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[0]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[0]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [0]),
        .O(\rgf/rgf_c0bus_0 [0]));
  LUT6 #(
    .INIT(64'h8C8C808C8C808080)) 
    \sr[10]_i_1 
       (.I0(\sr[10]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\sr[11]_i_3_n_0 ),
        .I3(\sr[11]_i_4_n_0 ),
        .I4(\rgf/sreg/sr [10]),
        .I5(\rgf/rgf_c0bus_0 [10]),
        .O(\rgf/sreg/p_0_in__0 [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[10]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/sreg/sr [10]),
        .O(\sr[10]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[10]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[10]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [10]),
        .O(\rgf/rgf_c0bus_0 [10]));
  LUT6 #(
    .INIT(64'h8C8C808C8C808080)) 
    \sr[11]_i_1 
       (.I0(\sr[11]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\sr[11]_i_3_n_0 ),
        .I3(\sr[11]_i_4_n_0 ),
        .I4(\rgf/sreg/sr [11]),
        .I5(\rgf/rgf_c0bus_0 [11]),
        .O(\rgf/sreg/p_0_in__0 [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_10 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(ctl_selc1[0]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_wb [0]),
        .O(\rgf/rctl/rgf_selc1 [0]));
  LUT4 #(
    .INIT(16'h0001)) 
    \sr[11]_i_11 
       (.I0(\rgf/rctl/p_0_in [2]),
        .I1(\rgf/rctl/p_0_in [0]),
        .I2(\rgf/rctl/p_0_in [1]),
        .I3(\pc[15]_i_11_n_0 ),
        .O(\rgf/c0bus_sel_cr [0]));
  LUT6 #(
    .INIT(64'h00000000000055F7)) 
    \sr[11]_i_12 
       (.I0(\bcmd[2]_INST_0_i_5_n_0 ),
        .I1(\fch/ir1 [10]),
        .I2(\rgf_selc1_rn_wb[2]_i_4_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_3_n_0 ),
        .I4(\sr[11]_i_13_n_0 ),
        .I5(\sr[11]_i_14_n_0 ),
        .O(\sr[11]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA0200AAAAAAAA)) 
    \sr[11]_i_13 
       (.I0(\rgf_selc1_rn_wb[2]_i_9_n_0 ),
        .I1(\sr[11]_i_15_n_0 ),
        .I2(\rgf_selc1_rn_wb[2]_i_22_n_0 ),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_21_n_0 ),
        .I5(\rgf_selc1_rn_wb[2]_i_20_n_0 ),
        .O(\sr[11]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AAA8A8A8A8)) 
    \sr[11]_i_14 
       (.I0(\rgf_selc1_rn_wb[1]_i_4_n_0 ),
        .I1(\rgf_selc1_rn_wb[2]_i_15_n_0 ),
        .I2(\sr[11]_i_16_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_6_n_0 ),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [10]),
        .O(\sr[11]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[11]_i_15 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [5]),
        .O(\sr[11]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hABAAAAAAAAAAAAAA)) 
    \sr[11]_i_16 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\rgf_selc1_rn_wb[0]_i_32_n_0 ),
        .I2(\badr[31]_INST_0_i_146_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_17_n_0 ),
        .I4(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I5(\fch/ir1 [2]),
        .O(\sr[11]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[11]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/sreg/sr [11]),
        .O(\sr[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAEBAAAA)) 
    \sr[11]_i_3 
       (.I0(ctl_sr_upd1),
        .I1(\rgf/rctl/rgf_selc1_rn [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [2]),
        .I3(\rgf/rctl/rgf_selc1_rn [0]),
        .I4(\rgf/rctl/rgf_selc1 [1]),
        .I5(\rgf/rctl/rgf_selc1 [0]),
        .O(\sr[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[11]_i_4 
       (.I0(ctl_sr_ldie1),
        .I1(\rgf/c0bus_sel_cr [0]),
        .O(\sr[11]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_5 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[11]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [11]),
        .O(\rgf/rgf_c0bus_0 [11]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_6 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(\rgf_selc1_rn_wb[1]_i_1_n_0 ),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_rn_wb [1]),
        .O(\rgf/rctl/rgf_selc1_rn [1]));
  LUT6 #(
    .INIT(64'h444E000E000A000E)) 
    \sr[11]_i_7 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(\sr[11]_i_12_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[2] ),
        .I4(\rgf/rctl/rgf_selc1_stat ),
        .I5(\rgf/rctl/rgf_selc1_rn_wb [2]),
        .O(\rgf/rctl/rgf_selc1_rn [2]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_8 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(ctl_selc1_rn),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_rn_wb [0]),
        .O(\rgf/rctl/rgf_selc1_rn [0]));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[11]_i_9 
       (.I0(fch_wrbufn1),
        .I1(fch_term),
        .I2(ctl_selc1[1]),
        .I3(\rgf/rctl/rgf_selc1_stat ),
        .I4(\rgf/rctl/rgf_selc1_wb [1]),
        .O(\rgf/rctl/rgf_selc1 [1]));
  LUT4 #(
    .INIT(16'hCF44)) 
    \sr[12]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [12]),
        .I2(\sr[13]_i_2_n_0 ),
        .I3(cpuid[0]),
        .O(\rgf/sreg/p_0_in__0 [12]));
  LUT4 #(
    .INIT(16'hCF44)) 
    \sr[13]_i_1 
       (.I0(\sr[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [13]),
        .I2(\sr[13]_i_2_n_0 ),
        .I3(cpuid[1]),
        .O(\rgf/sreg/p_0_in__0 [13]));
  LUT5 #(
    .INIT(32'h00000200)) 
    \sr[13]_i_2 
       (.I0(\sr[5]_i_3_n_0 ),
        .I1(ctl_sr_upd0),
        .I2(ctl_sr_ldie0),
        .I3(rst_n),
        .I4(\sr[11]_i_3_n_0 ),
        .O(\sr[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \sr[13]_i_3 
       (.I0(\fch/ir0 [11]),
        .I1(stat[2]),
        .I2(\bbus_o[0]_INST_0_i_8_n_0 ),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [1]),
        .I5(\sr[13]_i_4_n_0 ),
        .O(ctl_sr_ldie0));
  LUT6 #(
    .INIT(64'hFFFFDFFFFFFFFFFF)) 
    \sr[13]_i_4 
       (.I0(brdy),
        .I1(\stat[1]_i_15__0_n_0 ),
        .I2(ctl_fetch0_fl_i_35_n_0),
        .I3(\fch/ir0 [0]),
        .I4(\ccmd[1]_INST_0_i_13_n_0 ),
        .I5(\rgf_selc0_wb[1]_i_12_n_0 ),
        .O(\sr[13]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[14]_i_1 
       (.I0(\rgf/sreg/sr [14]),
        .I1(\sr[15]_i_2_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [14]));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[15]_i_1 
       (.I0(\rgf/sreg/sr [15]),
        .I1(\sr[15]_i_2_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [15]));
  LUT6 #(
    .INIT(64'h7780778004048004)) 
    \sr[15]_i_10 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [4]),
        .I3(\fch/ir1 [6]),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [7]),
        .O(\sr[15]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hDDDDDDDF)) 
    \sr[15]_i_2 
       (.I0(rst_n),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/c1bus_sel_cr [5]),
        .I3(ctl_sr_upd1),
        .I4(\sr[11]_i_4_n_0 ),
        .O(\sr[15]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00000100)) 
    \sr[15]_i_3 
       (.I0(\rgf/rctl/rgf_selc1_rn [2]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .I2(\rgf/rctl/rgf_selc1_rn [1]),
        .I3(\rgf/rctl/rgf_selc1 [1]),
        .I4(\rgf/rctl/rgf_selc1 [0]),
        .O(\rgf/c1bus_sel_cr [0]));
  LUT5 #(
    .INIT(32'h00000800)) 
    \sr[15]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [2]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1 [1]),
        .I4(\rgf/rctl/rgf_selc1 [0]),
        .O(\rgf/c1bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'hF400F000F5000000)) 
    \sr[15]_i_5 
       (.I0(\fch/ir1 [13]),
        .I1(\sr[15]_i_6_n_0 ),
        .I2(\sr[15]_i_7_n_0 ),
        .I3(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [14]),
        .O(ctl_sr_upd1));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[15]_i_6 
       (.I0(\fch/ir1 [12]),
        .I1(\fch/ir1 [11]),
        .O(\sr[15]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00B0F0B0)) 
    \sr[15]_i_7 
       (.I0(\sr[15]_i_8_n_0 ),
        .I1(\sr[15]_i_9_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [12]),
        .O(\sr[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0040004000C040C0)) 
    \sr[15]_i_8 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [12]),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [9]),
        .O(\sr[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h15FFFFFFFFFFFFFF)) 
    \sr[15]_i_9 
       (.I0(\niss_dsp_a1[32]_INST_0_i_30_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [12]),
        .I4(\rgf_selc1_wb[1]_i_23_n_0 ),
        .I5(\sr[15]_i_10_n_0 ),
        .O(\sr[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h8C8C808C8C808080)) 
    \sr[1]_i_1 
       (.I0(\sr[1]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\sr[11]_i_3_n_0 ),
        .I3(\sr[11]_i_4_n_0 ),
        .I4(\rgf/sreg/sr [1]),
        .I5(\rgf/rgf_c0bus_0 [1]),
        .O(\rgf/sreg/p_0_in__0 [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[1]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/sreg/sr [1]),
        .O(\sr[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[1]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[1]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [1]),
        .O(\rgf/rgf_c0bus_0 [1]));
  LUT5 #(
    .INIT(32'hAA080008)) 
    \sr[2]_i_1 
       (.I0(rst_n),
        .I1(\sr[2]_i_2_n_0 ),
        .I2(\sr[2]_i_3_n_0 ),
        .I3(\sr[11]_i_3_n_0 ),
        .I4(\sr[2]_i_4_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [2]));
  LUT6 #(
    .INIT(64'hCCAFCCA0CCAFCCAF)) 
    \sr[2]_i_2 
       (.I0(\rgf/rgf_c0bus_0 [2]),
        .I1(fch_irq_lev[0]),
        .I2(\rgf/c0bus_sel_cr [0]),
        .I3(ctl_sr_ldie1),
        .I4(\rgf/sreg/sr [2]),
        .I5(\rgf/c0bus_sel_cr [5]),
        .O(\sr[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00D020F0)) 
    \sr[2]_i_3 
       (.I0(ctl_sr_ldie0),
        .I1(ctl_sr_upd0),
        .I2(\sr[5]_i_3_n_0 ),
        .I3(\rgf/sreg/sr [2]),
        .I4(fch_irq_lev[0]),
        .O(\sr[2]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[2]_i_4 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/sreg/sr [2]),
        .O(\sr[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000AAA8AAAAAAAA)) 
    \sr[3]_i_1 
       (.I0(rst_n),
        .I1(\sr[3]_i_2_n_0 ),
        .I2(\sr[5]_i_3_n_0 ),
        .I3(\sr[3]_i_3_n_0 ),
        .I4(\sr[3]_i_4_n_0 ),
        .I5(\sr[3]_i_5_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [3]));
  LUT4 #(
    .INIT(16'hB1A0)) 
    \sr[3]_i_2 
       (.I0(ctl_sr_ldie1),
        .I1(\rgf/c0bus_sel_cr [0]),
        .I2(fch_irq_lev[1]),
        .I3(\rgf/sreg/sr [3]),
        .O(\sr[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0F0B800)) 
    \sr[3]_i_3 
       (.I0(\rgf/rctl/rgf_c0bus_wb [3]),
        .I1(\rgf/rctl/rgf_selc0_stat ),
        .I2(c0bus[3]),
        .I3(fch_term),
        .I4(fch_wrbufn0),
        .I5(\sr[11]_i_4_n_0 ),
        .O(\sr[3]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hF0F2FDFFF0F0F0F0)) 
    \sr[3]_i_4 
       (.I0(ctl_sr_ldie0),
        .I1(ctl_sr_upd0),
        .I2(\sr[11]_i_3_n_0 ),
        .I3(fch_irq_lev[1]),
        .I4(\rgf/sreg/sr [3]),
        .I5(\sr[5]_i_3_n_0 ),
        .O(\sr[3]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h57F7)) 
    \sr[3]_i_5 
       (.I0(\sr[11]_i_3_n_0 ),
        .I1(\rgf/sreg/sr [3]),
        .I2(\rgf/c1bus_sel_cr [0]),
        .I3(\rgf/rgf_c1bus_0 [3]),
        .O(\sr[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEAAAEA)) 
    \sr[4]_i_1 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr[5]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [4]),
        .I3(ctl_sr_upd0),
        .I4(alu_sr_flag0[0]),
        .I5(\sr[4]_i_4_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [4]));
  LUT6 #(
    .INIT(64'hAAABAAAAABABABAB)) 
    \sr[4]_i_10 
       (.I0(\sr[4]_i_18_n_0 ),
        .I1(\sr[4]_i_19_n_0 ),
        .I2(\sr[4]_i_20_n_0 ),
        .I3(\sr[4]_i_21_n_0 ),
        .I4(\sr[4]_i_22_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010000)) 
    \sr[4]_i_11 
       (.I0(\sr[4]_i_23_n_0 ),
        .I1(\sr[4]_i_24_n_0 ),
        .I2(\sr[4]_i_25_n_0 ),
        .I3(\sr[4]_i_26_n_0 ),
        .I4(\sr[4]_i_27_n_0 ),
        .I5(\sr[4]_i_28_n_0 ),
        .O(alu_sr_flag1[0]));
  LUT3 #(
    .INIT(8'h1F)) 
    \sr[4]_i_12 
       (.I0(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h8088AAAA80888088)) 
    \sr[4]_i_13 
       (.I0(\rgf_c0bus_wb[2]_i_4_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_8_n_0 ),
        .I2(\sr[4]_i_29_n_0 ),
        .I3(\sr[4]_i_30_n_0 ),
        .I4(\sr[4]_i_31_n_0 ),
        .I5(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\sr[4]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_14 
       (.I0(\rgf_c0bus_wb[22]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[28]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb[17]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_2_n_0 ),
        .O(\sr[4]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_15 
       (.I0(\rgf_c0bus_wb[24]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[25]_i_2_n_0 ),
        .O(\sr[4]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_16 
       (.I0(\rgf_c0bus_wb[20]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[26]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[23]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .O(\sr[4]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_17 
       (.I0(\rgf_c0bus_wb[19]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb[29]_i_3_n_0 ),
        .O(\sr[4]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[4]_i_18 
       (.I0(\sr[4]_i_32_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I2(\sr[4]_i_33_n_0 ),
        .I3(\sr[4]_i_34_n_0 ),
        .O(\sr[4]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_19 
       (.I0(\rgf_c0bus_wb[4]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[3]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_7_n_0 ),
        .I3(\sr[4]_i_35_n_0 ),
        .O(\sr[4]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \sr[4]_i_2 
       (.I0(\sr[11]_i_3_n_0 ),
        .I1(\sr[7]_i_2_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(ctl_sr_ldie1),
        .I4(\rgf/sreg/sr [4]),
        .O(\sr[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_20 
       (.I0(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[12]_i_9_n_0 ),
        .I3(\sr[4]_i_36_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[11]_i_9_n_0 ),
        .O(\sr[4]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_21 
       (.I0(\rgf_c0bus_wb[17]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[22]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[28]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_8_n_0 ),
        .I4(\sr[4]_i_37_n_0 ),
        .O(\sr[4]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \sr[4]_i_22 
       (.I0(\rgf_c0bus_wb[29]_i_5_n_0 ),
        .I1(\rgf_c0bus_wb[19]_i_5_n_0 ),
        .I2(\rgf_c0bus_wb[26]_i_5_n_0 ),
        .I3(\rgf_c0bus_wb[24]_i_5_n_0 ),
        .I4(\sr[4]_i_38_n_0 ),
        .O(\sr[4]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_23 
       (.I0(\sr[4]_i_39_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[14]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[12]_i_3_n_0 ),
        .I4(\rgf_c1bus_wb[8]_i_3_n_0 ),
        .O(\sr[4]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_24 
       (.I0(\rgf_c1bus_wb[1]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[4]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[10]_i_3_n_0 ),
        .O(\sr[4]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_25 
       (.I0(\rgf_c1bus_wb[3]_i_3_n_0 ),
        .I1(\rgf_c1bus_wb[13]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[2]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_3_n_0 ),
        .O(\sr[4]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_26 
       (.I0(\rgf_c1bus_wb[7]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_3_n_0 ),
        .I3(\rgf_c1bus_wb[11]_i_3_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_27 
       (.I0(\rgf_c1bus_wb[16]_i_4_n_0 ),
        .I1(\sr[4]_i_40_n_0 ),
        .I2(\sr[4]_i_41_n_0 ),
        .I3(\sr[4]_i_42_n_0 ),
        .I4(\sr[4]_i_43_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAAABAAAAAAABAAAB)) 
    \sr[4]_i_28 
       (.I0(\sr[4]_i_44_n_0 ),
        .I1(\sr[4]_i_45_n_0 ),
        .I2(\sr[4]_i_46_n_0 ),
        .I3(\sr[4]_i_47_n_0 ),
        .I4(\sr[4]_i_48_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h4540FFFF45404540)) 
    \sr[4]_i_29 
       (.I0(\niss_dsp_b0[4]_INST_0_i_1_n_0 ),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\sr[4]_i_49_n_0 ),
        .I4(\rgf_c0bus_wb[18]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_8_n_0 ),
        .O(\sr[4]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010000)) 
    \sr[4]_i_3 
       (.I0(\sr[4]_i_5_n_0 ),
        .I1(\sr[4]_i_6_n_0 ),
        .I2(\sr[4]_i_7_n_0 ),
        .I3(\sr[4]_i_8_n_0 ),
        .I4(\sr[4]_i_9_n_0 ),
        .I5(\sr[4]_i_10_n_0 ),
        .O(alu_sr_flag0[0]));
  LUT6 #(
    .INIT(64'hAAAAABFBFFFFABFB)) 
    \sr[4]_i_30 
       (.I0(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I1(\sr[4]_i_49_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[18]_i_18_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_14_n_0 ),
        .I5(a0bus_0[31]),
        .O(\sr[4]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAE00AEAEAEAE)) 
    \sr[4]_i_31 
       (.I0(\rgf_c0bus_wb[2]_i_10_n_0 ),
        .I1(\sr[4]_i_50_n_0 ),
        .I2(\sr[4]_i_51_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\sr[4]_i_52_n_0 ),
        .I5(\sr[4]_i_53_n_0 ),
        .O(\sr[4]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_32 
       (.I0(\sr[4]_i_54_n_0 ),
        .I1(\rgf_c0bus_wb_reg[19]_i_11_n_4 ),
        .I2(\rgf_c0bus_wb_reg[29]_i_11_n_7 ),
        .I3(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .I4(\sr[4]_i_55_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_33 
       (.I0(\sr[4]_i_56_n_0 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_12_n_6 ),
        .I2(\rgf_c0bus_wb_reg[15]_i_19_n_4 ),
        .I3(\rgf_c0bus_wb_reg[3]_i_11_n_7 ),
        .I4(\rgf_c0bus_wb_reg[15]_i_19_n_7 ),
        .I5(\sr[4]_i_57_n_0 ),
        .O(\sr[4]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'h0000D1C0)) 
    \sr[4]_i_34 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_62_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .I4(\rgf/sreg/sr [4]),
        .O(\sr[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_35 
       (.I0(\rgf_c0bus_wb[7]_i_7_n_0 ),
        .I1(\rgf_c0bus_wb[5]_i_7_n_0 ),
        .I2(\rgf_c0bus_wb[0]_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[2]_i_9_n_0 ),
        .I4(\sr[4]_i_58_n_0 ),
        .I5(\rgf_c0bus_wb[14]_i_9_n_0 ),
        .O(\sr[4]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_36 
       (.I0(\rgf_c0bus_wb[9]_i_9_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_9_n_0 ),
        .O(\sr[4]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_37 
       (.I0(\rgf_c0bus_wb[27]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[21]_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[25]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[30]_i_8_n_0 ),
        .O(\sr[4]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_38 
       (.I0(\rgf_c0bus_wb[23]_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[20]_i_8_n_0 ),
        .O(\sr[4]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \sr[4]_i_39 
       (.I0(\rgf_c1bus_wb[4]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_8_n_0 ),
        .O(\sr[4]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[4]_i_4 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\sr[7]_i_9_n_0 ),
        .I2(alu_sr_flag1[0]),
        .I3(\sr[11]_i_3_n_0 ),
        .I4(rst_n),
        .O(\sr[4]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_40 
       (.I0(\rgf_c1bus_wb[22]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[28]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[30]_i_4_n_0 ),
        .O(\sr[4]_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_41 
       (.I0(\rgf_c1bus_wb[24]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[27]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[18]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[25]_i_4_n_0 ),
        .O(\sr[4]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_42 
       (.I0(\rgf_c1bus_wb[20]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[26]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_4_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .O(\sr[4]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_43 
       (.I0(\rgf_c1bus_wb[19]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[29]_i_4_n_0 ),
        .O(\sr[4]_i_43_n_0 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[4]_i_44 
       (.I0(\sr[4]_i_59_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I2(\sr[4]_i_60_n_0 ),
        .I3(\sr[4]_i_61_n_0 ),
        .O(\sr[4]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_45 
       (.I0(\rgf_c1bus_wb[4]_i_10_n_0 ),
        .I1(\rgf_c1bus_wb[3]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[6]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[14]_i_5_n_0 ),
        .I4(\sr[4]_i_62_n_0 ),
        .I5(\sr[4]_i_63_n_0 ),
        .O(\sr[4]_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_46 
       (.I0(\rgf_c1bus_wb[11]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[8]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[13]_i_5_n_0 ),
        .I3(\rgf_c1bus_wb[9]_i_5_n_0 ),
        .O(\sr[4]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_47 
       (.I0(\rgf_c1bus_wb[12]_i_5_n_0 ),
        .I1(\rgf_c1bus_wb[10]_i_5_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .O(\sr[4]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \sr[4]_i_48 
       (.I0(\sr[4]_i_64_n_0 ),
        .I1(\rgf_c1bus_wb[18]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[20]_i_2_n_0 ),
        .I3(\sr[4]_i_65_n_0 ),
        .I4(\sr[4]_i_66_n_0 ),
        .I5(\sr[4]_i_67_n_0 ),
        .O(\sr[4]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \sr[4]_i_49 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[10]_i_28_n_0 ),
        .O(\sr[4]_i_49_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_5 
       (.I0(\sr[4]_i_12_n_0 ),
        .I1(\rgf_c0bus_wb[0]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[14]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[12]_i_2_n_0 ),
        .I4(\rgf_c0bus_wb[8]_i_2_n_0 ),
        .O(\sr[4]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hABAA)) 
    \sr[4]_i_50 
       (.I0(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\sr[4]_i_68_n_0 ),
        .I3(\sr[4]_i_69_n_0 ),
        .O(\sr[4]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF04C404C404C4)) 
    \sr[4]_i_51 
       (.I0(\rgf_c0bus_wb[18]_i_13_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[19]_i_19_n_0 ),
        .I4(\rgf_c0bus_wb[2]_i_20_n_0 ),
        .I5(\bbus_o[5]_INST_0_i_1_n_0 ),
        .O(\sr[4]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFD50000)) 
    \sr[4]_i_52 
       (.I0(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I1(\rgf_c0bus_wb[10]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_28_n_0 ),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I5(\rgf_c0bus_wb[2]_i_20_n_0 ),
        .O(\sr[4]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'hAAEFAAEFAAEFAAAA)) 
    \sr[4]_i_53 
       (.I0(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I1(\sr[4]_i_70_n_0 ),
        .I2(\sr[4]_i_71_n_0 ),
        .I3(\sr[4]_i_72_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(\sr[4]_i_68_n_0 ),
        .O(\sr[4]_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF0E0)) 
    \sr[4]_i_54 
       (.I0(\rgf_c0bus_wb_reg[19]_i_11_n_7 ),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_7 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb_reg[29]_i_11_n_5 ),
        .I4(\sr[4]_i_73_n_0 ),
        .O(\sr[4]_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hEEEA)) 
    \sr[4]_i_55 
       (.I0(\sr[4]_i_74_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb_reg[27]_i_23_n_5 ),
        .I3(\alu0/art/add/tout [18]),
        .O(\sr[4]_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_56 
       (.I0(\rgf_c0bus_wb_reg[3]_i_11_n_6 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_12_n_5 ),
        .I2(\rgf_c0bus_wb_reg[11]_i_20_n_5 ),
        .I3(\rgf_c0bus_wb_reg[15]_i_19_n_6 ),
        .O(\sr[4]_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_57 
       (.I0(\rgf_c0bus_wb_reg[11]_i_20_n_4 ),
        .I1(\rgf_c0bus_wb_reg[7]_i_12_n_4 ),
        .I2(\rgf_c0bus_wb_reg[15]_i_19_n_5 ),
        .I3(\rgf_c0bus_wb_reg[3]_i_11_n_4 ),
        .I4(\sr[4]_i_75_n_0 ),
        .O(\sr[4]_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFE0037)) 
    \sr[4]_i_58 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I5(\rgf_c0bus_wb[1]_i_7_n_0 ),
        .O(\sr[4]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_59 
       (.I0(\sr[4]_i_76_n_0 ),
        .I1(\rgf_c1bus_wb_reg[19]_i_10_n_4 ),
        .I2(\rgf_c1bus_wb_reg[31]_i_11_n_7 ),
        .I3(\rgf_c1bus_wb_reg[31]_i_11_n_4 ),
        .I4(\sr[4]_i_77_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_59_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_6 
       (.I0(\rgf_c0bus_wb[1]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[4]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .I3(\rgf_c0bus_wb[10]_i_2_n_0 ),
        .O(\sr[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_60 
       (.I0(\sr[4]_i_78_n_0 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_6 ),
        .I2(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I3(\rgf_c1bus_wb_reg[3]_i_20_n_7 ),
        .I4(\rgf_c1bus_wb_reg[19]_i_18_n_7 ),
        .I5(\sr[4]_i_79_n_0 ),
        .O(\sr[4]_i_60_n_0 ));
  LUT5 #(
    .INIT(32'h0000F888)) 
    \sr[4]_i_61 
       (.I0(\rgf_c1bus_wb[31]_i_24_n_0 ),
        .I1(dctl_sign_f_i_2_n_0),
        .I2(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .I3(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I4(\rgf/sreg/sr [4]),
        .O(\sr[4]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFE0037)) 
    \sr[4]_i_62 
       (.I0(acmd1[0]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(acmd1[3]),
        .I4(acmd1[4]),
        .I5(\rgf_c1bus_wb[1]_i_9_n_0 ),
        .O(\sr[4]_i_62_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_63 
       (.I0(\rgf_c1bus_wb[2]_i_9_n_0 ),
        .I1(\rgf_c1bus_wb[0]_i_9_n_0 ),
        .I2(\rgf_c1bus_wb[5]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_11_n_0 ),
        .O(\sr[4]_i_63_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \sr[4]_i_64 
       (.I0(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_9_n_0 ),
        .I2(\sr[4]_i_80_n_0 ),
        .I3(\rgf_c1bus_wb[23]_i_5_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[4]_i_65 
       (.I0(\rgf_c1bus_wb_reg[24]_i_2_n_0 ),
        .I1(\rgf_c1bus_wb_reg[26]_i_2_n_0 ),
        .I2(\sr[4]_i_81_n_0 ),
        .I3(\sr[4]_i_82_n_0 ),
        .I4(\rgf_c1bus_wb[19]_i_8_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_2_n_0 ),
        .O(\sr[4]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_66 
       (.I0(\rgf_c1bus_wb[27]_i_2_n_0 ),
        .I1(\sr[4]_i_83_n_0 ),
        .I2(\sr[4]_i_84_n_0 ),
        .I3(\rgf_c1bus_wb[21]_i_8_n_0 ),
        .I4(\rgf_c1bus_wb[25]_i_2_n_0 ),
        .I5(\rgf_c1bus_wb_reg[30]_i_2_n_0 ),
        .O(\sr[4]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_67 
       (.I0(\sr[4]_i_85_n_0 ),
        .I1(\sr[4]_i_86_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_2_n_0 ),
        .I3(\rgf_c1bus_wb[22]_i_2_n_0 ),
        .I4(\sr[4]_i_87_n_0 ),
        .I5(\sr[4]_i_88_n_0 ),
        .O(\sr[4]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h0000021333330213)) 
    \sr[4]_i_68 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[27]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I5(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .O(\sr[4]_i_68_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \sr[4]_i_69 
       (.I0(\rgf_c0bus_wb[18]_i_15_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[18]_i_16_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\sr[4]_i_69_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_7 
       (.I0(\rgf_c0bus_wb[3]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[13]_i_2_n_0 ),
        .I2(\sr[4]_i_13_n_0 ),
        .I3(\rgf_c0bus_wb[9]_i_2_n_0 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_70 
       (.I0(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[27]_i_27_n_0 ),
        .O(\sr[4]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h3030303030201000)) 
    \sr[4]_i_71 
       (.I0(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I3(\rgf_c0bus_wb[27]_i_24_n_0 ),
        .I4(\rgf_c0bus_wb[14]_i_27_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\sr[4]_i_71_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_72 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(a0bus_0[1]),
        .O(\sr[4]_i_72_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0F0E0)) 
    \sr[4]_i_73 
       (.I0(\rgf_c0bus_wb_reg[23]_i_24_n_5 ),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_6 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c0bus_wb_reg[19]_i_11_n_5 ),
        .I4(\rgf_c0bus_wb_reg[23]_i_24_n_7 ),
        .O(\sr[4]_i_73_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_74 
       (.I0(\rgf_c0bus_wb_reg[29]_i_11_n_6 ),
        .I1(\rgf_c0bus_wb_reg[27]_i_23_n_4 ),
        .I2(\rgf_c0bus_wb_reg[23]_i_24_n_4 ),
        .I3(\rgf_c0bus_wb_reg[23]_i_24_n_6 ),
        .O(\sr[4]_i_74_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_75 
       (.I0(\rgf_c0bus_wb_reg[3]_i_11_n_5 ),
        .I1(\rgf_c0bus_wb_reg[11]_i_20_n_7 ),
        .I2(\rgf_c0bus_wb_reg[7]_i_12_n_7 ),
        .I3(\rgf_c0bus_wb_reg[11]_i_20_n_6 ),
        .O(\sr[4]_i_75_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF0E0)) 
    \sr[4]_i_76 
       (.I0(\rgf_c1bus_wb_reg[19]_i_10_n_7 ),
        .I1(\rgf_c1bus_wb_reg[27]_i_10_n_7 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c1bus_wb_reg[31]_i_11_n_5 ),
        .I4(\sr[4]_i_89_n_0 ),
        .O(\sr[4]_i_76_n_0 ));
  LUT4 #(
    .INIT(16'hEEEA)) 
    \sr[4]_i_77 
       (.I0(\sr[4]_i_90_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb_reg[27]_i_10_n_5 ),
        .I3(\alu1/art/add/tout [18]),
        .O(\sr[4]_i_77_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_78 
       (.I0(\rgf_c1bus_wb_reg[3]_i_20_n_6 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_5 ),
        .I2(\rgf_c1bus_wb_reg[11]_i_10_n_5 ),
        .I3(\rgf_c1bus_wb_reg[19]_i_18_n_6 ),
        .O(\sr[4]_i_78_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_79 
       (.I0(\rgf_c1bus_wb_reg[11]_i_10_n_4 ),
        .I1(\rgf_c1bus_wb_reg[7]_i_23_n_4 ),
        .I2(\rgf_c1bus_wb_reg[19]_i_18_n_5 ),
        .I3(\rgf_c1bus_wb_reg[3]_i_20_n_4 ),
        .I4(\sr[4]_i_91_n_0 ),
        .O(\sr[4]_i_79_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_8 
       (.I0(\rgf_c0bus_wb[7]_i_3_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I2(\rgf_c0bus_wb[5]_i_3_n_0 ),
        .I3(\rgf_c0bus_wb[11]_i_2_n_0 ),
        .O(\sr[4]_i_8_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \sr[4]_i_80 
       (.I0(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_7_n_0 ),
        .I2(\rgf_c1bus_wb[23]_i_8_n_0 ),
        .O(\sr[4]_i_80_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_81 
       (.I0(\sr[4]_i_92_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(\rgf_c1bus_wb[19]_i_16_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_81_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_82 
       (.I0(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[19]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[19]_i_7_n_0 ),
        .O(\sr[4]_i_82_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_83 
       (.I0(\sr[4]_i_93_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(\rgf_c1bus_wb[21]_i_14_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_83_n_0 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \sr[4]_i_84 
       (.I0(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .I1(\rgf_c1bus_wb[21]_i_6_n_0 ),
        .I2(\rgf_c1bus_wb[21]_i_7_n_0 ),
        .O(\sr[4]_i_84_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_85 
       (.I0(\sr[4]_i_94_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(\rgf_c1bus_wb[16]_i_14_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_85_n_0 ));
  LUT5 #(
    .INIT(32'hFFF44444)) 
    \sr[4]_i_86 
       (.I0(\sr[4]_i_95_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr[4]_i_86_n_0 ));
  LUT5 #(
    .INIT(32'hFE0E0000)) 
    \sr[4]_i_87 
       (.I0(\sr[4]_i_96_n_0 ),
        .I1(\rgf_c1bus_wb[23]_i_17_n_0 ),
        .I2(dctl_sign_f_i_2_n_0),
        .I3(\rgf_c1bus_wb[17]_i_14_n_0 ),
        .I4(acmd1[0]),
        .O(\sr[4]_i_87_n_0 ));
  LUT5 #(
    .INIT(32'hFF4F4444)) 
    \sr[4]_i_88 
       (.I0(\sr[4]_i_97_n_0 ),
        .I1(\niss_dsp_a1[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c1bus_wb[17]_i_7_n_0 ),
        .I3(\rgf_c1bus_wb[17]_i_6_n_0 ),
        .I4(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr[4]_i_88_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0F0E0)) 
    \sr[4]_i_89 
       (.I0(\rgf_c1bus_wb_reg[23]_i_11_n_5 ),
        .I1(\rgf_c1bus_wb_reg[27]_i_10_n_6 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\rgf_c1bus_wb_reg[19]_i_10_n_5 ),
        .I4(\rgf_c1bus_wb_reg[23]_i_11_n_7 ),
        .O(\sr[4]_i_89_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_9 
       (.I0(\rgf_c0bus_wb[16]_i_2_n_0 ),
        .I1(\sr[4]_i_14_n_0 ),
        .I2(\sr[4]_i_15_n_0 ),
        .I3(\sr[4]_i_16_n_0 ),
        .I4(\sr[4]_i_17_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[4]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_90 
       (.I0(\rgf_c1bus_wb_reg[31]_i_11_n_6 ),
        .I1(\rgf_c1bus_wb_reg[27]_i_10_n_4 ),
        .I2(\rgf_c1bus_wb_reg[23]_i_11_n_4 ),
        .I3(\rgf_c1bus_wb_reg[23]_i_11_n_6 ),
        .O(\sr[4]_i_90_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_91 
       (.I0(\rgf_c1bus_wb_reg[3]_i_20_n_5 ),
        .I1(\rgf_c1bus_wb_reg[11]_i_10_n_7 ),
        .I2(\rgf_c1bus_wb_reg[7]_i_23_n_7 ),
        .I3(\rgf_c1bus_wb_reg[11]_i_10_n_6 ),
        .O(\sr[4]_i_91_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_92 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[19]),
        .I2(b1bus_0[19]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_92_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_93 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[21]),
        .I2(b1bus_0[21]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_93_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_94 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[16]),
        .I2(b1bus_0[16]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_94_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \sr[4]_i_95 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[16]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\sr[4]_i_95_n_0 ));
  LUT4 #(
    .INIT(16'hC444)) 
    \sr[4]_i_96 
       (.I0(\rgf_c1bus_wb[29]_i_15_n_0 ),
        .I1(a1bus_0[17]),
        .I2(b1bus_0[17]),
        .I3(\rgf_c1bus_wb[29]_i_16_n_0 ),
        .O(\sr[4]_i_96_n_0 ));
  LUT5 #(
    .INIT(32'hFF74CFFF)) 
    \sr[4]_i_97 
       (.I0(b1bus_0[7]),
        .I1(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I2(a1bus_0[17]),
        .I3(acmd1[4]),
        .I4(acmd1[3]),
        .O(\sr[4]_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h00000000EEEAAAEA)) 
    \sr[5]_i_1 
       (.I0(\sr[5]_i_2_n_0 ),
        .I1(\sr[5]_i_3_n_0 ),
        .I2(\rgf/sreg/sr [5]),
        .I3(ctl_sr_upd0),
        .I4(alu_sr_flag0[1]),
        .I5(\sr[5]_i_6_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [5]));
  LUT5 #(
    .INIT(32'hB0F0F0F0)) 
    \sr[5]_i_10 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .O(\sr[5]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h00000060)) 
    \sr[5]_i_11 
       (.I0(\rgf_c0bus_wb[16]_i_2_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I2(\bbus_o[4]_INST_0_i_1_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\sr[5]_i_18_n_0 ),
        .O(\sr[5]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF2A40)) 
    \sr[5]_i_12 
       (.I0(\alu1/mul_a_i [31]),
        .I1(\rgf_c1bus_wb_reg[31]_i_11_n_4 ),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu1/art/p_0_in__0 ),
        .I4(\sr[5]_i_20_n_0 ),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(\sr[5]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hAABABAAAAAAAAAAA)) 
    \sr[5]_i_13 
       (.I0(\sr[5]_i_21_n_0 ),
        .I1(\sr[5]_i_22_n_0 ),
        .I2(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I3(\sr[6]_i_19_n_0 ),
        .I4(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[5]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h000000C000C040C0)) 
    \sr[5]_i_14 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [9]),
        .I5(\fch/ir0 [8]),
        .O(\sr[5]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFF00F1F1FFFFF1F1)) 
    \sr[5]_i_15 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\ccmd[1]_INST_0_i_10_n_0 ),
        .I3(\sr[5]_i_23_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [9]),
        .O(\sr[5]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h82)) 
    \sr[5]_i_16 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\sr[6]_i_16_n_0 ),
        .I2(b0bus_0[31]),
        .O(\alu0/art/p_0_in__0 ));
  LUT5 #(
    .INIT(32'h1D1D0010)) 
    \sr[5]_i_17 
       (.I0(\alu0/asr0 ),
        .I1(\alu0/art/add/p_0_in ),
        .I2(\rgf_c0bus_wb_reg[15]_i_19_n_4 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\niss_dsp_a0[32]_INST_0_i_2_n_0 ),
        .O(\sr[5]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \sr[5]_i_18 
       (.I0(\niss_dsp_a0[32]_INST_0_i_6_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I2(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_7_n_0 ),
        .O(\sr[5]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'h82)) 
    \sr[5]_i_19 
       (.I0(\rgf/sreg/sr [8]),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(b1bus_0[31]),
        .O(\alu1/art/p_0_in__0 ));
  LUT5 #(
    .INIT(32'hFFEAAAEA)) 
    \sr[5]_i_2 
       (.I0(\sr[11]_i_3_n_0 ),
        .I1(\sr[7]_i_2_n_0 ),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(ctl_sr_ldie1),
        .I4(\rgf/sreg/sr [5]),
        .O(\sr[5]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h0C0C0010)) 
    \sr[5]_i_20 
       (.I0(\mul_a[16]_i_1__0_n_0 ),
        .I1(\alu1/art/add/p_0_in ),
        .I2(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\niss_dsp_a1[32]_INST_0_i_2_n_0 ),
        .O(\sr[5]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h00000060)) 
    \sr[5]_i_21 
       (.I0(\rgf_c1bus_wb[16]_i_4_n_0 ),
        .I1(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I2(\bdatw[12]_INST_0_i_4_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\sr[5]_i_22_n_0 ),
        .O(\sr[5]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \sr[5]_i_22 
       (.I0(\niss_dsp_a1[32]_INST_0_i_5_n_0 ),
        .I1(acmd1[3]),
        .I2(acmd1[4]),
        .I3(\rgf_c1bus_wb[23]_i_6_n_0 ),
        .O(\sr[5]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hD9FF7726)) 
    \sr[5]_i_23 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [5]),
        .O(\sr[5]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'hD8)) 
    \sr[5]_i_24 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[16]),
        .I2(a0bus_0[15]),
        .O(\alu0/asr0 ));
  LUT4 #(
    .INIT(16'hE12D)) 
    \sr[5]_i_25 
       (.I0(b0bus_0[15]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\sr[6]_i_16_n_0 ),
        .I3(b0bus_0[16]),
        .O(\alu0/art/add/p_0_in ));
  LUT3 #(
    .INIT(8'h01)) 
    \sr[5]_i_3 
       (.I0(ctl_sr_ldie1),
        .I1(\rgf/c0bus_sel_cr [0]),
        .I2(\rgf/c0bus_sel_cr [5]),
        .O(\sr[5]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h88CC8000880C8000)) 
    \sr[5]_i_4 
       (.I0(\sr[5]_i_7_n_0 ),
        .I1(\bbus_o[5]_INST_0_i_8_n_0 ),
        .I2(\fch/ir0 [14]),
        .I3(\fch/ir0 [13]),
        .I4(\fch/ir0 [15]),
        .I5(\sr[5]_i_8_n_0 ),
        .O(ctl_sr_upd0));
  LUT6 #(
    .INIT(64'hFFFFFFFFAEEAAAAA)) 
    \sr[5]_i_5 
       (.I0(\sr[5]_i_9_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .I3(\sr[6]_i_13_n_0 ),
        .I4(\sr[5]_i_10_n_0 ),
        .I5(\sr[5]_i_11_n_0 ),
        .O(alu_sr_flag0[1]));
  LUT6 #(
    .INIT(64'h44470000FFFFFFFF)) 
    \sr[5]_i_6 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\sr[7]_i_9_n_0 ),
        .I2(\sr[5]_i_12_n_0 ),
        .I3(\sr[5]_i_13_n_0 ),
        .I4(\sr[11]_i_3_n_0 ),
        .I5(rst_n),
        .O(\sr[5]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4444EEEE5444EEEE)) 
    \sr[5]_i_7 
       (.I0(\fch/ir0 [15]),
        .I1(\sr[5]_i_14_n_0 ),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [12]),
        .I5(\sr[5]_i_15_n_0 ),
        .O(\sr[5]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[5]_i_8 
       (.I0(\fch/ir0 [12]),
        .I1(\fch/ir0 [11]),
        .O(\sr[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0820)) 
    \sr[5]_i_9 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .I3(\alu0/art/p_0_in__0 ),
        .I4(\sr[5]_i_17_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .O(\sr[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF40)) 
    \sr[6]_i_1 
       (.I0(ctl_sr_ldie1),
        .I1(\rgf/rgf_c0bus_0 [6]),
        .I2(\sr[7]_i_2_n_0 ),
        .I3(\sr[6]_i_4_n_0 ),
        .I4(\sr[6]_i_5_n_0 ),
        .I5(\sr[6]_i_6_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [6]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF44F4)) 
    \sr[6]_i_10 
       (.I0(\rgf_c0bus_wb[31]_i_2_n_0 ),
        .I1(bdatr[6]),
        .I2(\rgf_c1bus_wb[6]_i_2_n_0 ),
        .I3(\rgf_c0bus_wb[6]_i_5_n_0 ),
        .I4(\rgf_c0bus_wb[6]_i_4_n_0 ),
        .I5(\rgf_c0bus_wb[6]_i_3_n_0 ),
        .O(\sr[6]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_11 
       (.I0(cbus_i[6]),
        .I1(ccmd[4]),
        .O(\sr[6]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h45401015)) 
    \sr[6]_i_12 
       (.I0(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I1(\alu0/art/add/tout [34]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\alu0/art/add/tout [18]),
        .I4(\sr[6]_i_16_n_0 ),
        .O(\sr[6]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FDFFF8F0)) 
    \sr[6]_i_13 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(\rgf_c0bus_wb[31]_i_30_n_0 ),
        .I3(\rgf_c0bus_wb[7]_i_25_n_0 ),
        .I4(\sr[6]_i_17_n_0 ),
        .I5(\sr[6]_i_18_n_0 ),
        .O(\sr[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEEEBBBEB)) 
    \sr[6]_i_14 
       (.I0(\sr[6]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_23_n_0 ),
        .I2(\alu1/art/add/tout [18]),
        .I3(\rgf/sreg/sr [8]),
        .I4(\alu1/art/add/tout [34]),
        .I5(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .O(alu_sr_flag1[2]));
  LUT6 #(
    .INIT(64'hEEEEEEAEFFFFFFAF)) 
    \sr[6]_i_16 
       (.I0(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .I1(\niss_dsp_a0[32]_INST_0_i_4_n_0 ),
        .I2(\rgf_c0bus_wb[7]_i_34_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_7_n_0 ),
        .I4(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_58_n_0 ),
        .O(\sr[6]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \sr[6]_i_17 
       (.I0(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_29_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(\sr[6]_i_23_n_0 ),
        .O(\sr[6]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hCCFCCCDD)) 
    \sr[6]_i_18 
       (.I0(\sr[6]_i_24_n_0 ),
        .I1(\sr[6]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_16_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\bbus_o[4]_INST_0_i_1_n_0 ),
        .O(\sr[6]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FBEAFFEA)) 
    \sr[6]_i_19 
       (.I0(\rgf_c1bus_wb[16]_i_19_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_33_n_0 ),
        .I2(\alu1/mul_a_i [31]),
        .I3(\sr[6]_i_26_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\sr[6]_i_27_n_0 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \sr[6]_i_2 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\sr[6]_i_7_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\bcmd[1]_INST_0_i_14_n_0 ),
        .I4(\sr[6]_i_8_n_0 ),
        .I5(\sr[6]_i_9_n_0 ),
        .O(ctl_sr_ldie1));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_21 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .O(\sr[6]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'h78)) 
    \sr[6]_i_22 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a0bus_0[31]),
        .I2(\alu0/art/p_0_in__0 ),
        .O(\sr[6]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAFAEFFFE0F0CFFFC)) 
    \sr[6]_i_23 
       (.I0(\sr[6]_i_30_n_0 ),
        .I1(\sr[6]_i_31_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I3(\sr[6]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[15]_i_26_n_0 ),
        .I5(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .O(\sr[6]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FEE0F0E)) 
    \sr[6]_i_24 
       (.I0(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I1(\sr[6]_i_23_n_0 ),
        .I2(\rgf_c0bus_wb[16]_i_14_n_0 ),
        .I3(\niss_dsp_a0[32]_INST_0_i_8_n_0 ),
        .I4(a0bus_0[31]),
        .I5(\rgf_c0bus_wb[16]_i_13_n_0 ),
        .O(\sr[6]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABAAA)) 
    \sr[6]_i_25 
       (.I0(\sr[4]_i_12_n_0 ),
        .I1(\sr[6]_i_33_n_0 ),
        .I2(\bbus_o[5]_INST_0_i_1_n_0 ),
        .I3(\rgf/sreg/sr [8]),
        .I4(\sr[6]_i_34_n_0 ),
        .O(\sr[6]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \sr[6]_i_26 
       (.I0(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[16]_i_33_n_0 ),
        .I3(acmd1[3]),
        .I4(\sr[6]_i_35_n_0 ),
        .O(\sr[6]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF00F1)) 
    \sr[6]_i_27 
       (.I0(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .I1(\sr[6]_i_35_n_0 ),
        .I2(\sr[6]_i_36_n_0 ),
        .I3(\niss_dsp_b1[4]_INST_0_i_1_n_0 ),
        .I4(\sr[6]_i_37_n_0 ),
        .O(\sr[6]_i_27_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_28 
       (.I0(\rgf/sreg/sr [8]),
        .I1(a1bus_0[31]),
        .O(\sr[6]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hEEE4EEE0AAA0EEE0)) 
    \sr[6]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(\sr[6]_i_10_n_0 ),
        .I3(\sr[6]_i_11_n_0 ),
        .I4(\rgf/rctl/rgf_selc0_stat ),
        .I5(\rgf/rctl/rgf_c0bus_wb [6]),
        .O(\rgf/rgf_c0bus_0 [6]));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[6]_i_30 
       (.I0(\rgf_c0bus_wb[31]_i_42_n_0 ),
        .I1(\remden[31]_i_3_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .O(\sr[6]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h002EFF2E00000000)) 
    \sr[6]_i_31 
       (.I0(\rgf_c0bus_wb[30]_i_45_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_47_n_0 ),
        .I3(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I4(\sr[6]_i_38_n_0 ),
        .I5(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\sr[6]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_32 
       (.I0(\rgf_c0bus_wb[7]_i_37_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .O(\sr[6]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h47FF474700FF0000)) 
    \sr[6]_i_33 
       (.I0(\rgf_c0bus_wb[23]_i_29_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I2(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I3(\rgf_c0bus_wb[16]_i_32_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_16_n_0 ),
        .I5(\rgf_c0bus_wb[7]_i_23_n_0 ),
        .O(\sr[6]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h0101015151510151)) 
    \sr[6]_i_34 
       (.I0(\rgf_c0bus_wb[14]_i_21_n_0 ),
        .I1(\rgf_c0bus_wb[15]_i_25_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_29_n_0 ),
        .I3(\sr[6]_i_39_n_0 ),
        .I4(\rgf_c0bus_wb[31]_i_25_n_0 ),
        .I5(\rgf_c0bus_wb[28]_i_30_n_0 ),
        .O(\sr[6]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h44FF000F4F4F0F0F)) 
    \sr[6]_i_35 
       (.I0(\rgf_c1bus_wb[31]_i_41_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_57_n_0 ),
        .I2(\sr[6]_i_40_n_0 ),
        .I3(\rgf_c1bus_wb[15]_i_30_n_0 ),
        .I4(acmd1[0]),
        .I5(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .O(\sr[6]_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hFBAA)) 
    \sr[6]_i_36 
       (.I0(\rgf_c1bus_wb[16]_i_21_n_0 ),
        .I1(a1bus_0[31]),
        .I2(acmd1[3]),
        .I3(\rgf_c1bus_wb[16]_i_22_n_0 ),
        .O(\sr[6]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF2020FF20)) 
    \sr[6]_i_37 
       (.I0(\bdatw[12]_INST_0_i_4_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[16]_i_24_n_0 ),
        .I3(\sr[6]_i_41_n_0 ),
        .I4(\sr[6]_i_42_n_0 ),
        .I5(\sr[4]_i_39_n_0 ),
        .O(\sr[6]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_38 
       (.I0(\rgf_c0bus_wb[30]_i_49_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\rgf_c0bus_wb[30]_i_46_n_0 ),
        .O(\sr[6]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'h88BBB8BB)) 
    \sr[6]_i_39 
       (.I0(\rgf_c0bus_wb[30]_i_59_n_0 ),
        .I1(\rgf_c0bus_wb[30]_i_34_n_0 ),
        .I2(\bbus_o[0]_INST_0_i_1_n_0 ),
        .I3(a0bus_0[31]),
        .I4(\niss_dsp_a0[32]_INST_0_i_3_n_0 ),
        .O(\sr[6]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \sr[6]_i_4 
       (.I0(\sr[11]_i_3_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(ctl_sr_ldie1),
        .O(\sr[6]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h1013)) 
    \sr[6]_i_40 
       (.I0(\sr[6]_i_43_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c1bus_wb[7]_i_30_n_0 ),
        .O(\sr[6]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h8888888880888000)) 
    \sr[6]_i_41 
       (.I0(\niss_dsp_b1[5]_INST_0_i_1_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\sr[6]_i_44_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_36_n_0 ),
        .I4(\rgf_c1bus_wb[24]_i_27_n_0 ),
        .I5(\rgf_c1bus_wb[10]_i_20_n_0 ),
        .O(\sr[6]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h4F44)) 
    \sr[6]_i_42 
       (.I0(\rgf_c1bus_wb[16]_i_31_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_38_n_0 ),
        .I2(\rgf_c1bus_wb[15]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[16]_i_34_n_0 ),
        .O(\sr[6]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0F000FFF0F220F22)) 
    \sr[6]_i_43 
       (.I0(a1bus_0[0]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(\rgf_c1bus_wb[28]_i_29_n_0 ),
        .I3(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I4(\sr[6]_i_45_n_0 ),
        .I5(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .O(\sr[6]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888B8BBB888)) 
    \sr[6]_i_44 
       (.I0(\rgf_c1bus_wb[28]_i_30_n_0 ),
        .I1(\rgf_c1bus_wb[31]_i_51_n_0 ),
        .I2(\rgf_c1bus_wb[30]_i_48_n_0 ),
        .I3(\rgf_c1bus_wb[29]_i_38_n_0 ),
        .I4(\sr[6]_i_46_n_0 ),
        .I5(\rgf_c1bus_wb[27]_i_45_n_0 ),
        .O(\sr[6]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \sr[6]_i_45 
       (.I0(a1bus_0[1]),
        .I1(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I2(a1bus_0[2]),
        .O(\sr[6]_i_45_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[6]_i_46 
       (.I0(\niss_dsp_b1[0]_INST_0_i_1_n_0 ),
        .I1(a1bus_0[31]),
        .O(\sr[6]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hA8A8A808)) 
    \sr[6]_i_5 
       (.I0(\sr[5]_i_3_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(ctl_sr_upd0),
        .I3(\sr[6]_i_12_n_0 ),
        .I4(\sr[6]_i_13_n_0 ),
        .O(\sr[6]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[6]_i_6 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\sr[7]_i_9_n_0 ),
        .I2(alu_sr_flag1[2]),
        .I3(\sr[11]_i_3_n_0 ),
        .I4(rst_n),
        .O(\sr[6]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[6]_i_7 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [1]),
        .I2(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [6]),
        .I5(\fch/ir1 [9]),
        .O(\sr[6]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[6]_i_8 
       (.I0(\fch/ir1 [11]),
        .I1(\fch/ir1 [7]),
        .O(\sr[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \sr[6]_i_9 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [12]),
        .I3(\fch/ir1 [15]),
        .I4(\fch/ir1 [0]),
        .I5(\niss_dsp_b1[0]_INST_0_i_8_n_0 ),
        .O(\sr[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFAE)) 
    \sr[7]_i_1 
       (.I0(\sr[11]_i_3_n_0 ),
        .I1(\sr[7]_i_2_n_0 ),
        .I2(\sr[7]_i_3_n_0 ),
        .I3(\sr[7]_i_4_n_0 ),
        .I4(\sr[7]_i_5_n_0 ),
        .I5(\sr[7]_i_6_n_0 ),
        .O(\rgf/sreg/p_0_in__0 [7]));
  LUT4 #(
    .INIT(16'hFFE2)) 
    \sr[7]_i_10 
       (.I0(\rgf_c1bus_wb[15]_i_3_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c1bus_wb[31]_i_4_n_0 ),
        .I3(\sr[7]_i_12_n_0 ),
        .O(alu_sr_flag1[3]));
  LUT6 #(
    .INIT(64'hCFCFCCCCAFAAAFAA)) 
    \sr[7]_i_11 
       (.I0(\rgf_c0bus_wb[15]_i_10_n_0 ),
        .I1(\rgf_c0bus_wb[31]_i_9_n_0 ),
        .I2(\rgf_c0bus_wb[31]_i_36_n_0 ),
        .I3(\rgf_c0bus_wb_reg[15]_i_19_n_4 ),
        .I4(\rgf_c0bus_wb_reg[29]_i_11_n_4 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[7]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hCFCFCCCCAFAAAFAA)) 
    \sr[7]_i_12 
       (.I0(\rgf_c1bus_wb[15]_i_7_n_0 ),
        .I1(\rgf_c1bus_wb_reg[31]_i_2_n_0 ),
        .I2(\rgf_c1bus_wb[31]_i_10_n_0 ),
        .I3(\rgf_c1bus_wb_reg[19]_i_18_n_4 ),
        .I4(\rgf_c1bus_wb_reg[31]_i_11_n_4 ),
        .I5(\rgf/sreg/sr [8]),
        .O(\sr[7]_i_12_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[7]_i_2 
       (.I0(\rgf/c0bus_sel_cr [0]),
        .I1(\rgf/c0bus_sel_cr [5]),
        .O(\sr[7]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAFFAAFFBABFFFFF)) 
    \sr[7]_i_3 
       (.I0(ctl_sr_ldie1),
        .I1(\rgf/rctl/rgf_c0bus_wb [7]),
        .I2(\rgf/rctl/rgf_selc0_stat ),
        .I3(c0bus[7]),
        .I4(fch_term),
        .I5(fch_wrbufn0),
        .O(\sr[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[7]_i_4 
       (.I0(ctl_sr_ldie1),
        .I1(\rgf/sreg/sr [7]),
        .O(\sr[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[7]_i_5 
       (.I0(\sr[5]_i_3_n_0 ),
        .I1(\sr[7]_i_8_n_0 ),
        .O(\sr[7]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'h4700FFFF)) 
    \sr[7]_i_6 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\sr[7]_i_9_n_0 ),
        .I2(alu_sr_flag1[3]),
        .I3(\sr[11]_i_3_n_0 ),
        .I4(rst_n),
        .O(\sr[7]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h0008)) 
    \sr[7]_i_7 
       (.I0(\rgf/rctl/p_0_in [1]),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\rgf/rctl/p_0_in [0]),
        .I3(\pc[15]_i_11_n_0 ),
        .O(\rgf/c0bus_sel_cr [5]));
  LUT6 #(
    .INIT(64'hFFE2FFFFFFE20000)) 
    \sr[7]_i_8 
       (.I0(\rgf_c0bus_wb[15]_i_2_n_0 ),
        .I1(\rgf/sreg/sr [8]),
        .I2(\rgf_c0bus_wb[31]_i_3_n_0 ),
        .I3(\sr[7]_i_11_n_0 ),
        .I4(ctl_sr_upd0),
        .I5(\rgf/sreg/sr [7]),
        .O(\sr[7]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h04000004)) 
    \sr[7]_i_9 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .I2(\rgf/rctl/rgf_selc1_rn [0]),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .I4(\rgf/rctl/rgf_selc1_rn [1]),
        .O(\sr[7]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h8C8C808C8C808080)) 
    \sr[8]_i_1 
       (.I0(\sr[8]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\sr[11]_i_3_n_0 ),
        .I3(\sr[11]_i_4_n_0 ),
        .I4(\rgf/sreg/sr [8]),
        .I5(\rgf/rgf_c0bus_0 [8]),
        .O(\rgf/sreg/p_0_in__0 [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[8]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/sreg/sr [8]),
        .O(\sr[8]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[8]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[8]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [8]),
        .O(\rgf/rgf_c0bus_0 [8]));
  LUT6 #(
    .INIT(64'h8C8C808C8C808080)) 
    \sr[9]_i_1 
       (.I0(\sr[9]_i_2_n_0 ),
        .I1(rst_n),
        .I2(\sr[11]_i_3_n_0 ),
        .I3(\sr[11]_i_4_n_0 ),
        .I4(\rgf/sreg/sr [9]),
        .I5(\rgf/rgf_c0bus_0 [9]),
        .O(\rgf/sreg/p_0_in__0 [9]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[9]_i_2 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [0]),
        .I2(\rgf/sreg/sr [9]),
        .O(\sr[9]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hE4E0A0E0)) 
    \sr[9]_i_3 
       (.I0(fch_wrbufn0),
        .I1(fch_term),
        .I2(c0bus[9]),
        .I3(\rgf/rctl/rgf_selc0_stat ),
        .I4(\rgf/rctl/rgf_c0bus_wb [9]),
        .O(\rgf/rgf_c0bus_0 [9]));
  CARRY4 \sr_reg[6]_i_15 
       (.CI(\rgf_c0bus_wb_reg[29]_i_11_n_0 ),
        .CO(\alu0/art/add/tout [34]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_21_n_0 }),
        .S({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_22_n_0 }));
  CARRY4 \sr_reg[6]_i_20 
       (.CI(\rgf_c1bus_wb_reg[31]_i_11_n_0 ),
        .CO(\alu1/art/add/tout [34]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_28_n_0 }),
        .S({\<const0> ,\<const0> ,\<const0> ,\art/add/sr[6]_i_29_n_0 }));
  LUT6 #(
    .INIT(64'hBBB0BBB0BB000B00)) 
    \stat[0]_i_1 
       (.I0(\fch/stat [2]),
        .I1(\stat[0]_i_2_n_0 ),
        .I2(\fadr[15]_INST_0_i_5_n_0 ),
        .I3(\rgf/pcnt/pc [1]),
        .I4(\fadr[15]_INST_0_i_8_n_0 ),
        .I5(\stat[0]_i_3_n_0 ),
        .O(\fch/fctl/stat_nx [0]));
  LUT6 #(
    .INIT(64'h00000000BABBBABA)) 
    \stat[0]_i_10 
       (.I0(\stat[0]_i_17_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\stat[0]_i_18_n_0 ),
        .I3(\fch/ir1 [1]),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\stat[0]_i_19_n_0 ),
        .O(\stat[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF13030000)) 
    \stat[0]_i_10__0 
       (.I0(\fch/ir0 [8]),
        .I1(brdy),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [7]),
        .I4(\stat[0]_i_16__0_n_0 ),
        .I5(\stat[0]_i_17__0_n_0 ),
        .O(\stat[0]_i_10__0_n_0 ));
  LUT3 #(
    .INIT(8'h6F)) 
    \stat[0]_i_10__1 
       (.I0(\fch/ir0 [13]),
        .I1(\fch/ir0 [14]),
        .I2(brdy),
        .O(\stat[0]_i_10__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAEAEEEE)) 
    \stat[0]_i_11 
       (.I0(\stat[0]_i_18__0_n_0 ),
        .I1(brdy),
        .I2(\fch/ir0 [6]),
        .I3(\stat[0]_i_19__0_n_0 ),
        .I4(\fch/ir0 [10]),
        .I5(\stat[0]_i_20_n_0 ),
        .O(\stat[0]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h5525FBFF)) 
    \stat[0]_i_11__0 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .O(\stat[0]_i_11__0_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_11__1 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [14]),
        .O(\stat[0]_i_11__1_n_0 ));
  LUT6 #(
    .INIT(64'hFF0DFF0DFF0DFFFF)) 
    \stat[0]_i_12 
       (.I0(\stat[0]_i_21_n_0 ),
        .I1(\stat[0]_i_22_n_0 ),
        .I2(\stat[0]_i_20_n_0 ),
        .I3(\stat[0]_i_23_n_0 ),
        .I4(\rgf_selc0_rn_wb[1]_i_16_n_0 ),
        .I5(\stat[0]_i_24__0_n_0 ),
        .O(\stat[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFD)) 
    \stat[0]_i_12__0 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [10]),
        .I5(\fch/ir0 [11]),
        .O(\stat[0]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004140)) 
    \stat[0]_i_12__1 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [11]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir1 [13]),
        .I4(\fch/ir1 [14]),
        .I5(\ctl1/stat_reg_n_0_[2] ),
        .O(\stat[0]_i_12__1_n_0 ));
  LUT6 #(
    .INIT(64'h5DFD555FFFFFFFFF)) 
    \stat[0]_i_13 
       (.I0(\stat[0]_i_8__0_n_0 ),
        .I1(stat[2]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [1]),
        .I5(\stat[0]_i_25_n_0 ),
        .O(\stat[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF4FFF5F5F5F5)) 
    \stat[0]_i_13__0 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [3]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [7]),
        .I4(\rgf_selc1_rn_wb[0]_i_6_n_0 ),
        .I5(\fch/ir1 [10]),
        .O(\stat[0]_i_13__0_n_0 ));
  LUT4 #(
    .INIT(16'h0040)) 
    \stat[0]_i_13__1 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .O(\stat[0]_i_13__1_n_0 ));
  LUT6 #(
    .INIT(64'h0300A0A000000000)) 
    \stat[0]_i_14 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [3]),
        .I3(\rgf/sreg/sr [9]),
        .I4(\stat[0]_i_20__0_n_0 ),
        .I5(\stat[0]_i_21__0_n_0 ),
        .O(\stat[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_14__0 
       (.I0(stat[2]),
        .I1(stat[0]),
        .O(\stat[0]_i_14__0_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \stat[0]_i_14__1 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [11]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [10]),
        .O(\stat[0]_i_14__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000F800)) 
    \stat[0]_i_15 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\stat[0]_i_22__0_n_0 ),
        .I2(\stat[0]_i_23__0_n_0 ),
        .I3(\fch/ir1 [10]),
        .I4(\fch/ir1 [11]),
        .I5(\stat[0]_i_24_n_0 ),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000004140)) 
    \stat[0]_i_15__0 
       (.I0(stat[0]),
        .I1(\fch/ir0 [11]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir0 [13]),
        .I4(stat[2]),
        .I5(\fch/ir0 [14]),
        .O(\stat[0]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000B0FF)) 
    \stat[0]_i_16 
       (.I0(\rgf_selc1_rn_wb[0]_i_33_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [10]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\stat[0]_i_25__0_n_0 ),
        .I5(\stat[0]_i_26__0_n_0 ),
        .O(\stat[0]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \stat[0]_i_16__0 
       (.I0(\fch/ir0 [9]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [11]),
        .O(\stat[0]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000ABABABA0)) 
    \stat[0]_i_17 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [3]),
        .I4(fch_irq_req),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\stat[0]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h15FF)) 
    \stat[0]_i_17__0 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(crdy),
        .I2(div_crdy0),
        .I3(stat[0]),
        .O(\stat[0]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'h82888088AA88AA88)) 
    \stat[0]_i_18 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [1]),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [0]),
        .I4(\rgf/ivec/iv [0]),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\stat[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h5A5AFAFADAF2FAFA)) 
    \stat[0]_i_18__0 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [6]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [5]),
        .O(\stat[0]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'hEEFEFEFFEEFEEEEF)) 
    \stat[0]_i_19 
       (.I0(\niss_dsp_a1[32]_INST_0_i_26_n_0 ),
        .I1(\fch/ir1 [2]),
        .I2(\fch/ir1 [1]),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [3]),
        .I5(\ctl1/stat_reg_n_0_[2] ),
        .O(\stat[0]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \stat[0]_i_19__0 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [5]),
        .O(\stat[0]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[0]_i_1__0 
       (.I0(\stat[0]_i_2__0_n_0 ),
        .I1(stat[1]),
        .I2(\fch/ir0 [15]),
        .I3(\fch/ir0 [12]),
        .I4(stat[2]),
        .I5(\stat[0]_i_3__2_n_0 ),
        .O(\ctl0/stat_nx [0]));
  LUT6 #(
    .INIT(64'h0005030500050005)) 
    \stat[0]_i_1__1 
       (.I0(\stat[0]_i_2__1_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [15]),
        .I3(\fch/ir1 [12]),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\stat[0]_i_3__1_n_0 ),
        .O(\ctl1/stat_nx [0]));
  LUT6 #(
    .INIT(64'h01010100FFFFFFFF)) 
    \stat[0]_i_1__2 
       (.I0(\stat[0]_i_2__2_n_0 ),
        .I1(\stat[0]_i_3__0_n_0 ),
        .I2(\stat[0]_i_4__1_n_0 ),
        .I3(\stat[0]_i_5_n_0 ),
        .I4(\stat[0]_i_6_n_0 ),
        .I5(\bcmd[0]_INST_0_i_3_n_0 ),
        .O(\stat[0]_i_1__2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_2 
       (.I0(\fch/stat [0]),
        .I1(\fch/stat [1]),
        .O(\stat[0]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \stat[0]_i_20 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [11]),
        .O(\stat[0]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h45)) 
    \stat[0]_i_20__0 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [4]),
        .O(\stat[0]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'hECFCFFFFECFCEFFF)) 
    \stat[0]_i_21 
       (.I0(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [7]),
        .I4(brdy),
        .I5(\fch/ir0 [3]),
        .O(\stat[0]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_21__0 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [10]),
        .O(\stat[0]_i_21__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0020002)) 
    \stat[0]_i_22 
       (.I0(\rgf/sreg/sr [9]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [3]),
        .I3(\stat[0]_i_26_n_0 ),
        .I4(brdy),
        .I5(ctl_fetch0_fl_i_21_n_0),
        .O(\stat[0]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[0]_i_22__0 
       (.I0(\fch/ir1 [9]),
        .I1(\fch/ir1 [6]),
        .O(\stat[0]_i_22__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF3700)) 
    \stat[0]_i_23 
       (.I0(\bbus_o[5]_INST_0_i_25_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [8]),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\stat[0]_i_27_n_0 ),
        .I5(stat[0]),
        .O(\stat[0]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'h0F0A000C)) 
    \stat[0]_i_23__0 
       (.I0(div_crdy1),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [7]),
        .O(\stat[0]_i_23__0_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4FFF4F4F4)) 
    \stat[0]_i_24 
       (.I0(dctl_sign_f_i_9_n_0),
        .I1(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I2(\stat[0]_i_27__0_n_0 ),
        .I3(\rgf_selc1_rn_wb[2]_i_16_n_0 ),
        .I4(\bcmd[1]_INST_0_i_26_n_0 ),
        .I5(\fch/ir1 [9]),
        .O(\stat[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h3333031033330313)) 
    \stat[0]_i_24__0 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\rgf_selc0_rn_wb[0]_i_32_n_0 ),
        .I2(\fch/ir0 [7]),
        .I3(\fch/ir0 [9]),
        .I4(\fch/ir0 [8]),
        .I5(\rgf/sreg/sr [8]),
        .O(\stat[0]_i_24__0_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF00F2)) 
    \stat[0]_i_25 
       (.I0(stat[2]),
        .I1(\fch/ir0 [1]),
        .I2(\stat[0]_i_28_n_0 ),
        .I3(\fch/ir0 [11]),
        .I4(\stat[0]_i_29_n_0 ),
        .O(\stat[0]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h5FDF5FF7F0F0F0F0)) 
    \stat[0]_i_25__0 
       (.I0(\fch/ir1 [3]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [6]),
        .I3(\fch/ir1 [5]),
        .I4(\fch/ir1 [4]),
        .I5(\fch/ir1 [10]),
        .O(\stat[0]_i_25__0_n_0 ));
  LUT3 #(
    .INIT(8'hCE)) 
    \stat[0]_i_26 
       (.I0(\fch/ir0 [4]),
        .I1(\fch/ir0 [5]),
        .I2(\fch/ir0 [7]),
        .O(\stat[0]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \stat[0]_i_26__0 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [9]),
        .I2(\fch/ir1 [11]),
        .O(\stat[0]_i_26__0_n_0 ));
  LUT6 #(
    .INIT(64'h2030300020300000)) 
    \stat[0]_i_27 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\ccmd[2]_INST_0_i_12_n_0 ),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\rgf/sreg/sr [8]),
        .O(\stat[0]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h4440000000400000)) 
    \stat[0]_i_27__0 
       (.I0(dctl_sign_f_i_4_n_0),
        .I1(\fch/ir1 [11]),
        .I2(\rgf/sreg/sr [8]),
        .I3(\fch/ir1 [7]),
        .I4(\fch/ir1 [8]),
        .I5(div_crdy1),
        .O(\stat[0]_i_27__0_n_0 ));
  LUT6 #(
    .INIT(64'h82888088AA88AA88)) 
    \stat[0]_i_28 
       (.I0(stat[0]),
        .I1(\fch/ir0 [1]),
        .I2(\fch/ir0 [3]),
        .I3(\fch/ir0 [0]),
        .I4(\rgf/ivec/iv [0]),
        .I5(brdy),
        .O(\stat[0]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0F0E0EE)) 
    \stat[0]_i_29 
       (.I0(\fch/ir0 [3]),
        .I1(fch_irq_req),
        .I2(brdy),
        .I3(\fch/ir0 [0]),
        .I4(\fch/ir0 [1]),
        .I5(stat[0]),
        .O(\stat[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF2F2F200F2F2F2F2)) 
    \stat[0]_i_2__0 
       (.I0(\stat[0]_i_4_n_0 ),
        .I1(\stat[0]_i_5__0_n_0 ),
        .I2(stat[1]),
        .I3(\stat[0]_i_6__1_n_0 ),
        .I4(\stat[0]_i_7__1_n_0 ),
        .I5(\stat[0]_i_8__0_n_0 ),
        .O(\stat[0]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hF200F2F2F200F200)) 
    \stat[0]_i_2__1 
       (.I0(\stat[0]_i_4__0_n_0 ),
        .I1(\stat[0]_i_5__1_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[1] ),
        .I3(\stat[0]_i_6__0_n_0 ),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(\fch/ir1 [1]),
        .O(\stat[0]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'h8888008088000888)) 
    \stat[0]_i_2__2 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(\stat[0]_i_8__1_n_0 ),
        .I2(\fch/ir0 [1]),
        .I3(\stat[0]_i_9__0_n_0 ),
        .I4(\fch/ir0 [0]),
        .I5(stat[1]),
        .O(\stat[0]_i_2__2_n_0 ));
  LUT6 #(
    .INIT(64'hCC000000CC007600)) 
    \stat[0]_i_3 
       (.I0(\fch/fch_issu1_ir ),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [1]),
        .I3(\fadr[15]_INST_0_i_6_n_0 ),
        .I4(fch_heir_nir_i_3_n_0),
        .I5(\fch/stat [2]),
        .O(\stat[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFEFFFFFFFFFF)) 
    \stat[0]_i_3__0 
       (.I0(\stat[0]_i_10__1_n_0 ),
        .I1(stat[2]),
        .I2(\fch/ir0 [15]),
        .I3(\mem/bctl/fch_term_fl ),
        .I4(\mem/bctl/ctl/p_0_in [5]),
        .I5(\bcmd[0]_INST_0_i_7_n_0 ),
        .O(\stat[0]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'hC4C4C404FFFFFFFF)) 
    \stat[0]_i_3__1 
       (.I0(\stat[0]_i_7_n_0 ),
        .I1(ctl_fetch1_fl_i_16_n_0),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\stat[0]_i_8_n_0 ),
        .I4(\stat[0]_i_9_n_0 ),
        .I5(\stat[1]_i_6_n_0 ),
        .O(\stat[0]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'hFEFFAAAAAAAAAAAA)) 
    \stat[0]_i_3__2 
       (.I0(\stat[1]_i_3__0_n_0 ),
        .I1(\stat[0]_i_9__1_n_0 ),
        .I2(\stat[0]_i_10__0_n_0 ),
        .I3(\stat[0]_i_11_n_0 ),
        .I4(\bcmd[2]_INST_0_i_8_n_0 ),
        .I5(\stat[0]_i_12_n_0 ),
        .O(\stat[0]_i_3__2_n_0 ));
  LUT6 #(
    .INIT(64'hFF8FFF8FFFCFCFCF)) 
    \stat[0]_i_4 
       (.I0(stat[0]),
        .I1(\stat[0]_i_13_n_0 ),
        .I2(\stat[2]_i_13__0_n_0 ),
        .I3(stat[2]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [11]),
        .O(\stat[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFF4FFF4FFF5F5F5F)) 
    \stat[0]_i_4__0 
       (.I0(\stat[0]_i_10_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\stat[0]_i_11__1_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[2] ),
        .I4(\fch/ir1 [3]),
        .I5(\fch/ir1 [11]),
        .O(\stat[0]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'hBFFFBFBFBFFCBFFC)) 
    \stat[0]_i_4__1 
       (.I0(stat[1]),
        .I1(\fch/ir0 [13]),
        .I2(\fch/ir0 [12]),
        .I3(\fch/ir0 [10]),
        .I4(stat[0]),
        .I5(\fch/ir0 [11]),
        .O(\stat[0]_i_4__1_n_0 ));
  LUT6 #(
    .INIT(64'h0020282800202222)) 
    \stat[0]_i_5 
       (.I0(\ccmd[0]_INST_0_i_14_n_0 ),
        .I1(stat[0]),
        .I2(\fch/ir0 [8]),
        .I3(\stat[0]_i_11__0_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [7]),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF04010400)) 
    \stat[0]_i_5__0 
       (.I0(\stat[0]_i_14__0_n_0 ),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [11]),
        .I4(\fch/ir0 [14]),
        .I5(\stat[0]_i_15__0_n_0 ),
        .O(\stat[0]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0C020000)) 
    \stat[0]_i_5__1 
       (.I0(\fch/ir1 [14]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [13]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\niss_dsp_a1[32]_INST_0_i_13_n_0 ),
        .I5(\stat[0]_i_12__1_n_0 ),
        .O(\stat[0]_i_5__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF014545)) 
    \stat[0]_i_6 
       (.I0(\stat[0]_i_12__0_n_0 ),
        .I1(\fch/ir0 [3]),
        .I2(stat[1]),
        .I3(\stat[0]_i_13__1_n_0 ),
        .I4(stat[0]),
        .I5(\stat[0]_i_14__1_n_0 ),
        .O(\stat[0]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFBFF)) 
    \stat[0]_i_6__0 
       (.I0(\stat[1]_i_11__0_n_0 ),
        .I1(\fch/ir1 [0]),
        .I2(\fch/ir1 [3]),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\ctl1/stat_reg_n_0_[2] ),
        .O(\stat[0]_i_6__0_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \stat[0]_i_6__1 
       (.I0(\fch/ir0 [14]),
        .I1(brdy),
        .I2(\fch/ir0 [1]),
        .O(\stat[0]_i_6__1_n_0 ));
  LUT6 #(
    .INIT(64'h000000002FFFFFFF)) 
    \stat[0]_i_7 
       (.I0(\stat[0]_i_13__0_n_0 ),
        .I1(\stat[0]_i_14_n_0 ),
        .I2(\fch/ir1 [8]),
        .I3(\fch/ir1 [9]),
        .I4(\fch/ir1 [11]),
        .I5(\stat[0]_i_15_n_0 ),
        .O(\stat[0]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \stat[0]_i_7__0 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [4]),
        .I2(\fch/ir0 [2]),
        .I3(\fch/ir0 [6]),
        .O(\stat[0]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \stat[0]_i_7__1 
       (.I0(stat[1]),
        .I1(\fch/ir0 [0]),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(\fch/ir0 [13]),
        .I4(stat[0]),
        .I5(\fch/ir0 [3]),
        .O(\stat[0]_i_7__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFAAAAEAEE)) 
    \stat[0]_i_8 
       (.I0(\stat[0]_i_16_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_12_n_0 ),
        .I2(\bcmd[1]_INST_0_i_26_n_0 ),
        .I3(\fch/ir1 [6]),
        .I4(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I5(ctl_fetch1_fl_i_13_n_0),
        .O(\stat[0]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h00000002)) 
    \stat[0]_i_8__0 
       (.I0(\stat[0]_i_7__0_n_0 ),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [8]),
        .I3(\fch/ir0 [10]),
        .I4(\fch/ir0 [9]),
        .O(\stat[0]_i_8__0_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \stat[0]_i_8__1 
       (.I0(\fch/ir0 [8]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [7]),
        .O(\stat[0]_i_8__1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000041710000)) 
    \stat[0]_i_9 
       (.I0(div_crdy1),
        .I1(\fch/ir1 [8]),
        .I2(\fch/ir1 [11]),
        .I3(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I4(\fch/ir1 [7]),
        .I5(dctl_sign_f_i_4_n_0),
        .O(\stat[0]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_9__0 
       (.I0(stat[0]),
        .I1(\fch/ir0 [3]),
        .O(\stat[0]_i_9__0_n_0 ));
  LUT6 #(
    .INIT(64'h4171000000000000)) 
    \stat[0]_i_9__1 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [11]),
        .I3(brdy),
        .I4(\ccmd[3]_INST_0_i_15_n_0 ),
        .I5(\fch/ir0 [10]),
        .O(\stat[0]_i_9__1_n_0 ));
  LUT6 #(
    .INIT(64'h020202020202A202)) 
    \stat[1]_i_1 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\stat[1]_i_2_n_0 ),
        .I2(\stat[1]_i_3__1_n_0 ),
        .I3(\fch/stat [1]),
        .I4(\fch/stat [0]),
        .I5(\fadr[15]_INST_0_i_8_n_0 ),
        .O(\fch/fctl/stat_nx [1]));
  LUT6 #(
    .INIT(64'h00000000202203E0)) 
    \stat[1]_i_10 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .I5(\bcmd[1]_INST_0_i_14_n_0 ),
        .O(\stat[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000015101510101)) 
    \stat[1]_i_10__0 
       (.I0(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I1(\ccmd[2]_INST_0_i_10_n_0 ),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(\stat[1]_i_16__0_n_0 ),
        .I4(\fch/ir0 [11]),
        .I5(\fch/ir0 [9]),
        .O(\stat[1]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \stat[1]_i_11 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\fch/ir0 [9]),
        .I2(\ccmd[2]_INST_0_i_10_n_0 ),
        .I3(stat[1]),
        .I4(\fch/ir0 [7]),
        .I5(\bcmd[3]_INST_0_i_9_n_0 ),
        .O(\stat[1]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \stat[1]_i_11__0 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [11]),
        .I2(\niss_dsp_a1[32]_INST_0_i_26_n_0 ),
        .I3(\fch/ir1 [2]),
        .I4(\fch/ir1 [14]),
        .O(\stat[1]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hDDFCFCCCDDFCFCFC)) 
    \stat[1]_i_12 
       (.I0(\stat[1]_i_17__0_n_0 ),
        .I1(\stat[1]_i_18__0_n_0 ),
        .I2(\ccmd[1]_INST_0_i_16_n_0 ),
        .I3(\fch/ir0 [7]),
        .I4(stat[0]),
        .I5(\rgf/sreg/sr [9]),
        .O(\stat[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000B0)) 
    \stat[1]_i_12__0 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\fch/ir1 [13]),
        .I2(\fch/ir1 [11]),
        .I3(\ctl1/stat_reg_n_0_[1] ),
        .I4(\ctl1/stat_reg_n_0_[2] ),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\stat[1]_i_12__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFAFAFAFFBFFFB)) 
    \stat[1]_i_13 
       (.I0(\stat[1]_i_19__0_n_0 ),
        .I1(brdy),
        .I2(\fch/ir0 [11]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [7]),
        .I5(\fch/ir0 [6]),
        .O(\stat[1]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB0)) 
    \stat[1]_i_13__0 
       (.I0(\fch/ir1 [13]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir1 [14]),
        .O(\stat[1]_i_13__0_n_0 ));
  LUT6 #(
    .INIT(64'h1555FFFFFFFFFFFF)) 
    \stat[1]_i_14 
       (.I0(\stat[1]_i_20__0_n_0 ),
        .I1(stat[0]),
        .I2(\fch/ir0 [7]),
        .I3(\stat[1]_i_21_n_0 ),
        .I4(\stat[1]_i_22__0_n_0 ),
        .I5(\fch/ir0 [10]),
        .O(\stat[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h00000020000A0020)) 
    \stat[1]_i_14__0 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [14]),
        .I5(\rgf/sreg/sr [5]),
        .O(\stat[1]_i_14__0_n_0 ));
  LUT5 #(
    .INIT(32'hA65656A6)) 
    \stat[1]_i_15 
       (.I0(\fch/ir1 [11]),
        .I1(\rgf/sreg/sr [4]),
        .I2(\fch/ir1 [14]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\rgf/sreg/sr [7]),
        .O(\stat[1]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[1]_i_15__0 
       (.I0(stat[1]),
        .I1(stat[0]),
        .O(\stat[1]_i_15__0_n_0 ));
  LUT6 #(
    .INIT(64'h5F00FFF75FFFFFF7)) 
    \stat[1]_i_16 
       (.I0(div_crdy1),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\rgf/sreg/sr [10]),
        .I3(\fch/ir1 [8]),
        .I4(\fch/ir1 [11]),
        .I5(\stat[1]_i_24_n_0 ),
        .O(\stat[1]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \stat[1]_i_16__0 
       (.I0(\fch/ir0 [10]),
        .I1(\fch/ir0 [8]),
        .I2(brdy),
        .I3(\fch/ir0 [6]),
        .I4(\fch/ir0 [7]),
        .O(\stat[1]_i_16__0_n_0 ));
  LUT6 #(
    .INIT(64'hAEFFFFFFAEAEAEAE)) 
    \stat[1]_i_17 
       (.I0(\fch/ir1 [7]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [8]),
        .I5(\rgf/sreg/sr [11]),
        .O(\stat[1]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[1]_i_17__0 
       (.I0(\fch/ir0 [8]),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\stat[1]_i_17__0_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAEFEE)) 
    \stat[1]_i_18 
       (.I0(\rgf/sreg/sr [11]),
        .I1(\bcmd[2]_INST_0_i_6_n_0 ),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(div_crdy1),
        .I4(\fch/ir1 [11]),
        .I5(\fch/ir1 [8]),
        .O(\stat[1]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h2400000000000000)) 
    \stat[1]_i_18__0 
       (.I0(\fch/ir0 [5]),
        .I1(\fch/ir0 [7]),
        .I2(\fch/ir0 [4]),
        .I3(stat[0]),
        .I4(\fch/ir0 [3]),
        .I5(\fch/ir0 [8]),
        .O(\stat[1]_i_18__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFBF00FFFFFFFF)) 
    \stat[1]_i_19 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_31_n_0 ),
        .I2(\stat[1]_i_25_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\ctl1/stat_reg_n_0_[0] ),
        .I5(\ctl1/stat_reg_n_0_[1] ),
        .O(\stat[1]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \stat[1]_i_19__0 
       (.I0(stat[1]),
        .I1(\fch/ir0 [9]),
        .I2(\fch/ir0 [10]),
        .O(\stat[1]_i_19__0_n_0 ));
  LUT6 #(
    .INIT(64'h00001010000000FF)) 
    \stat[1]_i_1__0 
       (.I0(\ctl1/stat_reg_n_0_[2] ),
        .I1(\stat[1]_i_2__1_n_0 ),
        .I2(\stat[1]_i_3_n_0 ),
        .I3(\stat[1]_i_4_n_0 ),
        .I4(\fch/ir1 [15]),
        .I5(\fch/ir1 [12]),
        .O(\ctl1/stat_nx [1]));
  LUT6 #(
    .INIT(64'hEAEAEAEAAAEAAAAA)) 
    \stat[1]_i_1__1 
       (.I0(\stat[1]_i_2__0_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(stat[1]),
        .I4(\stat[1]_i_3__0_n_0 ),
        .I5(\stat[1]_i_4__0_n_0 ),
        .O(\ctl0/stat_nx [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \stat[1]_i_1__2 
       (.I0(\bcmd[0]_INST_0_i_7_n_0 ),
        .I1(\mem/bctl/fch_term_fl ),
        .I2(\mem/bctl/ctl/p_0_in [5]),
        .O(\mem/bctl/ctl/stat_nx ));
  LUT5 #(
    .INIT(32'h2F3A2F30)) 
    \stat[1]_i_2 
       (.I0(\fadr[15]_INST_0_i_16_n_0 ),
        .I1(\fadr[15]_INST_0_i_10_n_0 ),
        .I2(\fch/stat [1]),
        .I3(\fch/stat [0]),
        .I4(fch_leir_nir_i_2_n_0),
        .O(\stat[1]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAABBAABBAFBBAABB)) 
    \stat[1]_i_20 
       (.I0(\fch/ir1 [11]),
        .I1(div_crdy1),
        .I2(\rgf_selc1_rn_wb[2]_i_14_n_0 ),
        .I3(\bcmd[2]_INST_0_i_6_n_0 ),
        .I4(\rgf_selc1_wb[1]_i_31_n_0 ),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\stat[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F000000E)) 
    \stat[1]_i_20__0 
       (.I0(\stat[1]_i_23__0_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\rgf/sreg/sr [11]),
        .I3(\fch/ir0 [8]),
        .I4(\fch/ir0 [11]),
        .I5(\stat[1]_i_24__0_n_0 ),
        .O(\stat[1]_i_20__0_n_0 ));
  LUT6 #(
    .INIT(64'hD0101310D0101010)) 
    \stat[1]_i_21 
       (.I0(\rgf_selc0_rn_wb[1]_i_17_n_0 ),
        .I1(\fch/ir0 [8]),
        .I2(\fch/ir0 [11]),
        .I3(\ccmd[2]_INST_0_i_10_n_0 ),
        .I4(\rgf/sreg/sr [10]),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\stat[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \stat[1]_i_21__0 
       (.I0(\rgf_selc1_rn_wb[2]_i_19_n_0 ),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [8]),
        .I3(\bcmd[2]_INST_0_i_5_n_0 ),
        .I4(\fch/ir1 [9]),
        .I5(\fch/ir1 [7]),
        .O(\stat[1]_i_21__0_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[1]_i_22 
       (.I0(\fch/ir1 [10]),
        .I1(\fch/ir1 [9]),
        .O(\stat[1]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_22__0 
       (.I0(stat[1]),
        .I1(\fch/ir0 [9]),
        .O(\stat[1]_i_22__0_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFF77F)) 
    \stat[1]_i_23 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [11]),
        .I2(\fch/ir1 [7]),
        .I3(\fch/ir1 [6]),
        .I4(\stat[1]_i_26_n_0 ),
        .I5(\stat[1]_i_27_n_0 ),
        .O(\stat[1]_i_23_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \stat[1]_i_23__0 
       (.I0(div_crdy0),
        .I1(crdy),
        .I2(stat[0]),
        .O(\stat[1]_i_23__0_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \stat[1]_i_24 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\fch/ir1 [6]),
        .O(\stat[1]_i_24_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \stat[1]_i_24__0 
       (.I0(stat[0]),
        .I1(\rgf/sreg/sr [8]),
        .I2(\fch/ir0 [7]),
        .O(\stat[1]_i_24__0_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \stat[1]_i_25 
       (.I0(\fch/ir1 [6]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .O(\stat[1]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF3C3FFFFFF2)) 
    \stat[1]_i_26 
       (.I0(\rgf/sreg/sr [9]),
        .I1(\ctl1/stat_reg_n_0_[0] ),
        .I2(\fch/ir1 [3]),
        .I3(\fch/ir1 [4]),
        .I4(\fch/ir1 [5]),
        .I5(\fch/ir1 [7]),
        .O(\stat[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \stat[1]_i_27 
       (.I0(\rgf_selc1_wb[1]_i_29_n_0 ),
        .I1(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I2(\bcmd[2]_INST_0_i_6_n_0 ),
        .I3(\fch/ir1 [11]),
        .I4(\fch/ir1 [8]),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\stat[1]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h1010101011101111)) 
    \stat[1]_i_2__0 
       (.I0(\fch/ir0 [15]),
        .I1(\fch/ir0 [12]),
        .I2(\stat[1]_i_5_n_0 ),
        .I3(\stat[1]_i_6__0_n_0 ),
        .I4(\stat[1]_i_7__0_n_0 ),
        .I5(\stat[1]_i_8__0_n_0 ),
        .O(\stat[1]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'h1114441455555555)) 
    \stat[1]_i_2__1 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [11]),
        .I2(\rgf/sreg/sr [4]),
        .I3(\fch/ir1 [14]),
        .I4(\stat[1]_i_5__0_n_0 ),
        .I5(\bcmd[2]_INST_0_i_5_n_0 ),
        .O(\stat[1]_i_2__1_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF111311111111)) 
    \stat[1]_i_3 
       (.I0(\stat[1]_i_6_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(dctl_sign_f_i_4_n_0),
        .I3(\stat[1]_i_7_n_0 ),
        .I4(\stat[1]_i_8_n_0 ),
        .I5(\fch/ir1 [14]),
        .O(\stat[1]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h004F00400010001F)) 
    \stat[1]_i_3__0 
       (.I0(\fch/ir0 [14]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir0 [13]),
        .I3(stat[0]),
        .I4(\stat[1]_i_9__0_n_0 ),
        .I5(\fch/ir0 [11]),
        .O(\stat[1]_i_3__0_n_0 ));
  LUT5 #(
    .INIT(32'h55554540)) 
    \stat[1]_i_3__1 
       (.I0(\fch/stat [2]),
        .I1(\fch/fch_issu1 ),
        .I2(\fch/fch_term_fl ),
        .I3(\fch/fch_issu1_fl ),
        .I4(\fch/stat [0]),
        .O(\stat[1]_i_3__1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F2F200F2)) 
    \stat[1]_i_4 
       (.I0(\stat[1]_i_9_n_0 ),
        .I1(\stat[1]_i_10_n_0 ),
        .I2(\stat[1]_i_11__0_n_0 ),
        .I3(\stat[1]_i_12__0_n_0 ),
        .I4(\stat[1]_i_13__0_n_0 ),
        .I5(\stat[1]_i_14__0_n_0 ),
        .O(\stat[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8AAA8AAAAAAAA)) 
    \stat[1]_i_4__0 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\stat[1]_i_10__0_n_0 ),
        .I2(\stat[1]_i_11_n_0 ),
        .I3(\stat[1]_i_12_n_0 ),
        .I4(\stat[1]_i_13_n_0 ),
        .I5(\stat[1]_i_14_n_0 ),
        .O(\stat[1]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h0A0A0F00BA8ABA8A)) 
    \stat[1]_i_5 
       (.I0(fch_heir_nir_i_7_n_0),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [14]),
        .I3(\stat[2]_i_4_n_0 ),
        .I4(\rgf/sreg/sr [6]),
        .I5(\fch/ir0 [13]),
        .O(\stat[1]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \stat[1]_i_5__0 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .O(\stat[1]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFF3CAAAA)) 
    \stat[1]_i_6 
       (.I0(\stat[1]_i_15_n_0 ),
        .I1(\fch/ir1 [11]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [13]),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\stat[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0005000000050010)) 
    \stat[1]_i_6__0 
       (.I0(\rgf_selc0_rn_wb[1]_i_5_n_0 ),
        .I1(brdy),
        .I2(\fch/ir0 [3]),
        .I3(stat[2]),
        .I4(\fch/ir0 [0]),
        .I5(\fch/ir0 [1]),
        .O(\stat[1]_i_6__0_n_0 ));
  LUT5 #(
    .INIT(32'hBF00BFBF)) 
    \stat[1]_i_7 
       (.I0(\stat[1]_i_16_n_0 ),
        .I1(\fch/ir1 [7]),
        .I2(\ctl1/stat_reg_n_0_[0] ),
        .I3(\stat[1]_i_17_n_0 ),
        .I4(\stat[1]_i_18_n_0 ),
        .O(\stat[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFBAFBEBFFFFFBEF)) 
    \stat[1]_i_7__0 
       (.I0(\stat[1]_i_15__0_n_0 ),
        .I1(\fch/ir0 [0]),
        .I2(\fch/ir0 [3]),
        .I3(stat[2]),
        .I4(\fch/ir0 [1]),
        .I5(brdy),
        .O(\stat[1]_i_7__0_n_0 ));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4F4F4FF)) 
    \stat[1]_i_8 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(\stat[1]_i_20_n_0 ),
        .I2(\stat[1]_i_21__0_n_0 ),
        .I3(\stat[1]_i_22_n_0 ),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\stat[1]_i_23_n_0 ),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \stat[1]_i_8__0 
       (.I0(\fch/ir0 [11]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(ctl_fetch0_fl_i_29_n_0),
        .I4(\stat[0]_i_7__0_n_0 ),
        .I5(\stat[2]_i_13__0_n_0 ),
        .O(\stat[1]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFBF3F3FFFFF)) 
    \stat[1]_i_9 
       (.I0(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\niss_dsp_a1[32]_INST_0_i_13_n_0 ),
        .I3(\fch/ir1 [1]),
        .I4(\fch/ir1 [0]),
        .I5(\fch/ir1 [3]),
        .O(\stat[1]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h6F60)) 
    \stat[1]_i_9__0 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [14]),
        .I3(\rgf/sreg/sr [4]),
        .O(\stat[1]_i_9__0_n_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    \stat[2]_i_1 
       (.I0(\fch/rst_n_fl ),
        .O(\stat[2]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h8F00800000000000)) 
    \stat[2]_i_10 
       (.I0(\stat[2]_i_13_n_0 ),
        .I1(\rgf_selc1_wb[1]_i_33_n_0 ),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [12]),
        .I4(\stat[1]_i_5__0_n_0 ),
        .I5(\fch/ir1 [14]),
        .O(\stat[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00000ACF)) 
    \stat[2]_i_10__0 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [12]),
        .I5(\stat[2]_i_14__0_n_0 ),
        .O(\stat[2]_i_10__0_n_0 ));
  LUT6 #(
    .INIT(64'h37FFF7FFF7FFF7FF)) 
    \stat[2]_i_11 
       (.I0(\stat[1]_i_5__0_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [14]),
        .I4(\stat[2]_i_15_n_0 ),
        .I5(\fch_irq_lev[1]_i_3_n_0 ),
        .O(\stat[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF7FFFDFFFFFFF)) 
    \stat[2]_i_11__0 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [6]),
        .I2(\fch/ir1 [3]),
        .I3(\stat[2]_i_14_n_0 ),
        .I4(\fch/ir1 [7]),
        .I5(\fch/ir1 [4]),
        .O(\stat[2]_i_11__0_n_0 ));
  LUT6 #(
    .INIT(64'hAA2AA2AAAAAAAAAA)) 
    \stat[2]_i_12 
       (.I0(stat[0]),
        .I1(\fch/ir0 [3]),
        .I2(\fch/ir0 [4]),
        .I3(\fch/ir0 [7]),
        .I4(\fch/ir0 [6]),
        .I5(\stat[2]_i_16_n_0 ),
        .O(\stat[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h9000000000000000)) 
    \stat[2]_i_12__0 
       (.I0(\fch/ir1 [5]),
        .I1(\fch/ir1 [4]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [14]),
        .I4(\fch/ir1 [12]),
        .I5(\fch/ir1 [10]),
        .O(\stat[2]_i_12__0_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \stat[2]_i_13 
       (.I0(\fch/ir1 [8]),
        .I1(\fch/ir1 [7]),
        .I2(\fch/ir1 [9]),
        .I3(\fch/ir1 [10]),
        .O(\stat[2]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[2]_i_13__0 
       (.I0(\fch/ir0 [14]),
        .I1(\fch/ir0 [13]),
        .O(\stat[2]_i_13__0_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[2]_i_14 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\fch/ir1 [9]),
        .O(\stat[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBBBAAABAAABAAABA)) 
    \stat[2]_i_14__0 
       (.I0(stat[0]),
        .I1(\fch/ir0 [14]),
        .I2(\rgf/sreg/sr [4]),
        .I3(\fch/ir0 [13]),
        .I4(\rgf/sreg/sr [7]),
        .I5(\fch/ir0 [12]),
        .O(\stat[2]_i_14__0_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \stat[2]_i_15 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [10]),
        .I2(\fch/ir0 [9]),
        .I3(\fch/ir0 [8]),
        .O(\stat[2]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000080)) 
    \stat[2]_i_16 
       (.I0(\bcmd[2]_INST_0_i_8_n_0 ),
        .I1(\fch/ir0 [12]),
        .I2(\fch/ir0 [10]),
        .I3(\fch/ir0 [4]),
        .I4(\fch/ir0 [5]),
        .I5(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\stat[2]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h0005003500050005)) 
    \stat[2]_i_1__0 
       (.I0(\stat[2]_i_2__0_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[2] ),
        .I2(\fch/ir1 [11]),
        .I3(\fch/ir1 [15]),
        .I4(\ctl1/stat_reg_n_0_[1] ),
        .I5(\stat[2]_i_3__0_n_0 ),
        .O(\ctl1/stat_nx [2]));
  LUT6 #(
    .INIT(64'h5555510055555555)) 
    \stat[2]_i_1__1 
       (.I0(\fch/ir0 [15]),
        .I1(\stat[2]_i_2__1_n_0 ),
        .I2(\stat[2]_i_3__1_n_0 ),
        .I3(\stat[2]_i_4_n_0 ),
        .I4(\stat[2]_i_5_n_0 ),
        .I5(\stat[2]_i_6_n_0 ),
        .O(\stat[2]_i_1__1_n_0 ));
  LUT6 #(
    .INIT(64'hA0A0A2AA0000222A)) 
    \stat[2]_i_2 
       (.I0(\fadr[15]_INST_0_i_5_n_0 ),
        .I1(\fch/stat [0]),
        .I2(\fch/stat [2]),
        .I3(\fch/fch_issu1_ir ),
        .I4(\stat[2]_i_3_n_0 ),
        .I5(\fadr[15]_INST_0_i_10_n_0 ),
        .O(\fch/fctl/stat_nx [2]));
  LUT6 #(
    .INIT(64'h005D5D5D5D5D5D5D)) 
    \stat[2]_i_2__0 
       (.I0(\rgf_selc1_wb[0]_i_6_n_0 ),
        .I1(\stat[2]_i_4__0_n_0 ),
        .I2(\stat[2]_i_5__0_n_0 ),
        .I3(ctl_fetch1_fl_i_11_n_0),
        .I4(\stat[2]_i_6__0_n_0 ),
        .I5(\stat[2]_i_7_n_0 ),
        .O(\stat[2]_i_2__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFAAFFFFFFCCF0FF)) 
    \stat[2]_i_2__1 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [6]),
        .I2(\rgf/sreg/sr [5]),
        .I3(\fch/ir0 [14]),
        .I4(\fch/ir0 [13]),
        .I5(\fch/ir0 [12]),
        .O(\stat[2]_i_2__1_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF444)) 
    \stat[2]_i_3 
       (.I0(\fadr[15]_INST_0_i_7_n_0 ),
        .I1(\nir_id[24]_i_6_n_0 ),
        .I2(\fch/stat [0]),
        .I3(\fch/stat [1]),
        .I4(fch_term),
        .O(\stat[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00FBFFFF00FB00FB)) 
    \stat[2]_i_3__0 
       (.I0(\stat[2]_i_8_n_0 ),
        .I1(\stat[2]_i_9_n_0 ),
        .I2(\stat[2]_i_10_n_0 ),
        .I3(\ctl1/stat_reg_n_0_[0] ),
        .I4(\stat[2]_i_11__0_n_0 ),
        .I5(\stat[2]_i_12__0_n_0 ),
        .O(\stat[2]_i_3__0_n_0 ));
  LUT6 #(
    .INIT(64'h0900090000000F00)) 
    \stat[2]_i_3__1 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir0 [13]),
        .I3(\fch/ir0 [12]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\fch/ir0 [14]),
        .O(\stat[2]_i_3__1_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \stat[2]_i_4 
       (.I0(stat[0]),
        .I1(stat[1]),
        .I2(\fch/ir0 [11]),
        .I3(stat[2]),
        .O(\stat[2]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFCFCFFFF0AFAF)) 
    \stat[2]_i_4__0 
       (.I0(\rgf/sreg/sr [6]),
        .I1(\rgf/sreg/sr [7]),
        .I2(\fch/ir1 [13]),
        .I3(\rgf/sreg/sr [5]),
        .I4(\fch/ir1 [14]),
        .I5(\fch/ir1 [12]),
        .O(\stat[2]_i_4__0_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \stat[2]_i_5 
       (.I0(\stat[2]_i_7__0_n_0 ),
        .I1(\fch/ir0 [6]),
        .I2(\fch/ir0 [2]),
        .I3(\rgf_selc0_wb[1]_i_3_n_0 ),
        .I4(\stat[2]_i_8__0_n_0 ),
        .I5(\stat[2]_i_9__0_n_0 ),
        .O(\stat[2]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0900090000000F00)) 
    \stat[2]_i_5__0 
       (.I0(\rgf/sreg/sr [7]),
        .I1(\rgf/sreg/sr [5]),
        .I2(\fch/ir1 [13]),
        .I3(\fch/ir1 [12]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\fch/ir1 [14]),
        .O(\stat[2]_i_5__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFF4FFFFFFFF)) 
    \stat[2]_i_6 
       (.I0(\stat[2]_i_10__0_n_0 ),
        .I1(\stat[2]_i_11_n_0 ),
        .I2(\stat[2]_i_12_n_0 ),
        .I3(stat[2]),
        .I4(stat[1]),
        .I5(\fch/ir0 [11]),
        .O(\stat[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4544544544445444)) 
    \stat[2]_i_6__0 
       (.I0(\niss_dsp_a1[32]_INST_0_i_26_n_0 ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\ctl1/stat_reg_n_0_[2] ),
        .I3(\fch/ir1 [0]),
        .I4(\fch/ir1 [3]),
        .I5(\ctl1/stat_reg_n_0_[0] ),
        .O(\stat[2]_i_6__0_n_0 ));
  LUT6 #(
    .INIT(64'hFF4F44F4000000F0)) 
    \stat[2]_i_7 
       (.I0(\ctl1/stat_reg_n_0_[0] ),
        .I1(\ctl1/stat_reg_n_0_[1] ),
        .I2(\fch/ir1 [0]),
        .I3(\fch/ir1 [3]),
        .I4(\fch/ir1 [1]),
        .I5(\rgf_selc1_rn_wb[1]_i_15_n_0 ),
        .O(\stat[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF2F22F2000000F0)) 
    \stat[2]_i_7__0 
       (.I0(stat[1]),
        .I1(stat[0]),
        .I2(\fch/ir0 [0]),
        .I3(\fch/ir0 [3]),
        .I4(\fch/ir0 [1]),
        .I5(brdy),
        .O(\stat[2]_i_7__0_n_0 ));
  LUT4 #(
    .INIT(16'h0080)) 
    \stat[2]_i_8 
       (.I0(\fch/ir1 [13]),
        .I1(\fch/ir1 [12]),
        .I2(\rgf/sreg/sr [7]),
        .I3(\fch/ir1 [14]),
        .O(\stat[2]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \stat[2]_i_8__0 
       (.I0(\fch/ir0 [7]),
        .I1(\fch/ir0 [8]),
        .I2(\rgf_selc0_rn_wb[2]_i_25_n_0 ),
        .I3(\stat[2]_i_13__0_n_0 ),
        .I4(\fch/ir0 [12]),
        .I5(\fch/ir0 [11]),
        .O(\stat[2]_i_8__0_n_0 ));
  LUT6 #(
    .INIT(64'hFFDDFFDDCF00CFCC)) 
    \stat[2]_i_9 
       (.I0(\rgf/sreg/sr [5]),
        .I1(\fch/ir1 [12]),
        .I2(\rgf/sreg/sr [6]),
        .I3(\fch/ir1 [13]),
        .I4(\rgf/sreg/sr [4]),
        .I5(\fch/ir1 [14]),
        .O(\stat[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFBFBB6BF)) 
    \stat[2]_i_9__0 
       (.I0(\fch/ir0 [3]),
        .I1(\fch/ir0 [0]),
        .I2(stat[2]),
        .I3(stat[0]),
        .I4(stat[1]),
        .O(\stat[2]_i_9__0_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[0]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [0]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [0]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [0]),
        .O(\rgf/treg/p_1_in [0]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[10]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [10]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [10]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [10]),
        .O(\rgf/treg/p_1_in [10]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[11]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [11]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [11]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [11]),
        .O(\rgf/treg/p_1_in [11]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[12]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [12]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [12]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [12]),
        .O(\rgf/treg/p_1_in [12]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[13]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [13]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [13]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [13]),
        .O(\rgf/treg/p_1_in [13]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[14]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [14]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [14]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [14]),
        .O(\rgf/treg/p_1_in [14]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[15]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [15]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [15]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [15]),
        .O(\rgf/treg/p_1_in [15]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[16]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [16]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [16]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [16]),
        .O(\rgf/treg/p_1_in [16]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[17]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [17]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [17]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [17]),
        .O(\rgf/treg/p_1_in [17]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[18]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [18]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [18]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [18]),
        .O(\rgf/treg/p_1_in [18]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[19]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [19]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [19]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [19]),
        .O(\rgf/treg/p_1_in [19]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[1]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [1]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [1]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [1]),
        .O(\rgf/treg/p_1_in [1]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[20]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [20]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [20]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [20]),
        .O(\rgf/treg/p_1_in [20]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[21]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [21]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [21]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [21]),
        .O(\rgf/treg/p_1_in [21]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[22]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [22]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [22]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [22]),
        .O(\rgf/treg/p_1_in [22]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[23]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [23]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [23]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [23]),
        .O(\rgf/treg/p_1_in [23]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[24]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [24]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [24]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [24]),
        .O(\rgf/treg/p_1_in [24]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[25]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [25]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [25]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [25]),
        .O(\rgf/treg/p_1_in [25]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[26]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [26]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [26]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [26]),
        .O(\rgf/treg/p_1_in [26]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[27]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [27]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [27]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [27]),
        .O(\rgf/treg/p_1_in [27]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[28]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [28]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [28]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [28]),
        .O(\rgf/treg/p_1_in [28]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[29]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [29]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [29]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [29]),
        .O(\rgf/treg/p_1_in [29]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[2]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [2]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [2]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [2]),
        .O(\rgf/treg/p_1_in [2]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[30]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [30]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [30]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [30]),
        .O(\rgf/treg/p_1_in [30]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[31]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [31]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [31]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [31]),
        .O(\rgf/treg/p_1_in [31]));
  LUT4 #(
    .INIT(16'h0400)) 
    \tr[31]_i_2 
       (.I0(\rgf/rctl/rgf_selc1 [0]),
        .I1(\rgf/rctl/rgf_selc1 [1]),
        .I2(\tr[31]_i_4_n_0 ),
        .I3(\rgf/rctl/rgf_selc1_rn [2]),
        .O(\rgf/c1bus_sel_cr [4]));
  LUT3 #(
    .INIT(8'h04)) 
    \tr[31]_i_3 
       (.I0(\grn[15]_i_4__2_n_0 ),
        .I1(\rgf/rctl/p_0_in [2]),
        .I2(\pc[15]_i_11_n_0 ),
        .O(\rgf/c0bus_sel_cr [4]));
  LUT2 #(
    .INIT(4'hE)) 
    \tr[31]_i_4 
       (.I0(\rgf/rctl/rgf_selc1_rn [1]),
        .I1(\rgf/rctl/rgf_selc1_rn [0]),
        .O(\tr[31]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[3]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [3]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [3]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [3]),
        .O(\rgf/treg/p_1_in [3]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[4]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [4]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [4]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [4]),
        .O(\rgf/treg/p_1_in [4]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[5]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [5]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [5]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [5]),
        .O(\rgf/treg/p_1_in [5]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[6]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [6]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [6]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [6]),
        .O(\rgf/treg/p_1_in [6]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[7]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [7]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [7]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [7]),
        .O(\rgf/treg/p_1_in [7]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[8]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [8]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [8]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [8]),
        .O(\rgf/treg/p_1_in [8]));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[9]_i_1 
       (.I0(\rgf/rgf_c1bus_0 [9]),
        .I1(\rgf/c1bus_sel_cr [4]),
        .I2(\rgf/rgf_c0bus_0 [9]),
        .I3(\rgf/c0bus_sel_cr [4]),
        .I4(\rgf/treg/tr [9]),
        .O(\rgf/treg/p_1_in [9]));
endmodule
