
module niho_alu
   (mul_rslt,
    dctl_sign_f,
    div_crdy,
    niho_dsp_b,
    div_crdy_reg,
    \niho_dsp_c[31] ,
    mul_rslt_reg,
    Q,
    \rem_reg[30] ,
    \remden_reg[13] ,
    \remden_reg[15] ,
    \remden_reg[22] ,
    \remden_reg[23] ,
    \remden_reg[24] ,
    \remden_reg[26] ,
    \remden_reg[25] ,
    \remden_reg[21] ,
    \remden_reg[20] ,
    \remden_reg[19] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] ,
    \remden_reg[12] ,
    \remden_reg[14] ,
    div_crdy_reg_0,
    crdy_0,
    div_crdy_reg_1,
    mulh,
    mul_a,
    \mul_b_reg[32] ,
    \mul_b_reg[30] ,
    \mul_b_reg[29] ,
    \mul_b_reg[28] ,
    \mul_b_reg[27] ,
    \mul_b_reg[26] ,
    \mul_b_reg[25] ,
    \mul_b_reg[24] ,
    \mul_b_reg[23] ,
    \mul_b_reg[22] ,
    \mul_b_reg[21] ,
    \mul_b_reg[20] ,
    \mul_b_reg[19] ,
    \mul_b_reg[18] ,
    \mul_b_reg[17] ,
    \mul_b_reg[16] ,
    \mul_b_reg[15] ,
    \mul_b_reg[14] ,
    \mul_b_reg[13] ,
    \mul_b_reg[12] ,
    \mul_b_reg[11] ,
    \mul_b_reg[10] ,
    \mul_b_reg[9] ,
    \mul_b_reg[8] ,
    \mul_b_reg[7] ,
    \mul_b_reg[6] ,
    \mul_b_reg[5] ,
    \mul_b_reg[3] ,
    \mul_b_reg[2] ,
    \mul_b_reg[1] ,
    \mul_b_reg[0] ,
    p_0_in,
    mul_rslt0,
    clk,
    dctl_sign,
    rgf_sr_nh,
    \niho_dsp_b[4] ,
    \niho_dsp_b[4]_0 ,
    abus_0,
    niho_dsp_c,
    \tr[31]_i_5 ,
    \tr[31]_i_5_0 ,
    \dctl_stat_reg[2] ,
    crdy,
    \bcmd[2]_INST_0_i_1 ,
    rst_n,
    out,
    \niho_dsp_a[32]_INST_0_i_12 ,
    \dso_reg[19] ,
    \dso_reg[19]_0 ,
    \dso_reg[19]_1 ,
    \dso_reg[19]_2 ,
    \dso_reg[23] ,
    \dso_reg[23]_0 ,
    \dso_reg[23]_1 ,
    \dso_reg[23]_2 ,
    \dso_reg[27] ,
    \dso_reg[27]_0 ,
    \dso_reg[27]_1 ,
    \dso_reg[27]_2 ,
    \dso_reg[31] ,
    \dso_reg[31]_0 ,
    \dso_reg[31]_1 ,
    \dso_reg[31]_2 ,
    \remden_reg[31] ,
    \remden_reg[29] ,
    \remden_reg[25]_0 ,
    \remden_reg[24]_0 ,
    \remden_reg[23]_0 ,
    \remden_reg[22]_0 ,
    \remden_reg[21]_0 ,
    \remden_reg[20]_0 ,
    \remden_reg[18]_0 ,
    \remden_reg[17]_0 ,
    \remden_reg[16]_0 ,
    \remden_reg[30] ,
    \remden_reg[19]_0 ,
    \mulh_reg[0] ,
    mul_b,
    D,
    mul_a_i,
    \mul_a_reg[16] ,
    \mul_b_reg[0]_0 ,
    \mul_b_reg[32]_0 ,
    bbus_0,
    \remden_reg[28] ,
    \remden_reg[27] ,
    \remden_reg[26]_0 );
  output mul_rslt;
  output dctl_sign_f;
  output div_crdy;
  output [0:0]niho_dsp_b;
  output div_crdy_reg;
  output \niho_dsp_c[31] ;
  output mul_rslt_reg;
  output [30:0]Q;
  output [30:0]\rem_reg[30] ;
  output \remden_reg[13] ;
  output \remden_reg[15] ;
  output \remden_reg[22] ;
  output \remden_reg[23] ;
  output \remden_reg[24] ;
  output \remden_reg[26] ;
  output \remden_reg[25] ;
  output \remden_reg[21] ;
  output \remden_reg[20] ;
  output \remden_reg[19] ;
  output \remden_reg[18] ;
  output \remden_reg[17] ;
  output \remden_reg[16] ;
  output \remden_reg[12] ;
  output \remden_reg[14] ;
  output div_crdy_reg_0;
  output crdy_0;
  output div_crdy_reg_1;
  output [15:0]mulh;
  output [32:0]mul_a;
  output [1:0]\mul_b_reg[32] ;
  output \mul_b_reg[30] ;
  output \mul_b_reg[29] ;
  output \mul_b_reg[28] ;
  output \mul_b_reg[27] ;
  output \mul_b_reg[26] ;
  output \mul_b_reg[25] ;
  output \mul_b_reg[24] ;
  output \mul_b_reg[23] ;
  output \mul_b_reg[22] ;
  output \mul_b_reg[21] ;
  output \mul_b_reg[20] ;
  output \mul_b_reg[19] ;
  output \mul_b_reg[18] ;
  output \mul_b_reg[17] ;
  output \mul_b_reg[16] ;
  output \mul_b_reg[15] ;
  output \mul_b_reg[14] ;
  output \mul_b_reg[13] ;
  output \mul_b_reg[12] ;
  output \mul_b_reg[11] ;
  output \mul_b_reg[10] ;
  output \mul_b_reg[9] ;
  output \mul_b_reg[8] ;
  output \mul_b_reg[7] ;
  output \mul_b_reg[6] ;
  output \mul_b_reg[5] ;
  output \mul_b_reg[3] ;
  output \mul_b_reg[2] ;
  output \mul_b_reg[1] ;
  output \mul_b_reg[0] ;
  input p_0_in;
  input mul_rslt0;
  input clk;
  input dctl_sign;
  input rgf_sr_nh;
  input \niho_dsp_b[4] ;
  input \niho_dsp_b[4]_0 ;
  input [15:0]abus_0;
  input [15:0]niho_dsp_c;
  input \tr[31]_i_5 ;
  input \tr[31]_i_5_0 ;
  input \dctl_stat_reg[2] ;
  input crdy;
  input \bcmd[2]_INST_0_i_1 ;
  input rst_n;
  input [0:0]out;
  input [0:0]\niho_dsp_a[32]_INST_0_i_12 ;
  input \dso_reg[19] ;
  input \dso_reg[19]_0 ;
  input \dso_reg[19]_1 ;
  input \dso_reg[19]_2 ;
  input \dso_reg[23] ;
  input \dso_reg[23]_0 ;
  input \dso_reg[23]_1 ;
  input \dso_reg[23]_2 ;
  input \dso_reg[27] ;
  input \dso_reg[27]_0 ;
  input \dso_reg[27]_1 ;
  input \dso_reg[27]_2 ;
  input \dso_reg[31] ;
  input \dso_reg[31]_0 ;
  input \dso_reg[31]_1 ;
  input \dso_reg[31]_2 ;
  input \remden_reg[31] ;
  input \remden_reg[29] ;
  input \remden_reg[25]_0 ;
  input \remden_reg[24]_0 ;
  input \remden_reg[23]_0 ;
  input \remden_reg[22]_0 ;
  input \remden_reg[21]_0 ;
  input \remden_reg[20]_0 ;
  input \remden_reg[18]_0 ;
  input \remden_reg[17]_0 ;
  input \remden_reg[16]_0 ;
  input \remden_reg[30] ;
  input \remden_reg[19]_0 ;
  input \mulh_reg[0] ;
  input mul_b;
  input [1:0]D;
  input [13:0]mul_a_i;
  input \mul_a_reg[16] ;
  input \mul_b_reg[0]_0 ;
  input [1:0]\mul_b_reg[32]_0 ;
  input [30:0]bbus_0;
  input \remden_reg[28] ;
  input \remden_reg[27] ;
  input \remden_reg[26]_0 ;

  wire [1:0]D;
  wire [30:0]Q;
  wire [15:0]abus_0;
  wire [30:0]bbus_0;
  wire \bcmd[2]_INST_0_i_1 ;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[2] ;
  wire div_crdy;
  wire div_crdy_reg;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire \dso_reg[19] ;
  wire \dso_reg[19]_0 ;
  wire \dso_reg[19]_1 ;
  wire \dso_reg[19]_2 ;
  wire \dso_reg[23] ;
  wire \dso_reg[23]_0 ;
  wire \dso_reg[23]_1 ;
  wire \dso_reg[23]_2 ;
  wire \dso_reg[27] ;
  wire \dso_reg[27]_0 ;
  wire \dso_reg[27]_1 ;
  wire \dso_reg[27]_2 ;
  wire \dso_reg[31] ;
  wire \dso_reg[31]_0 ;
  wire \dso_reg[31]_1 ;
  wire \dso_reg[31]_2 ;
  wire [32:0]mul_a;
  wire [13:0]mul_a_i;
  wire \mul_a_reg[16] ;
  wire mul_b;
  wire \mul_b_reg[0] ;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[10] ;
  wire \mul_b_reg[11] ;
  wire \mul_b_reg[12] ;
  wire \mul_b_reg[13] ;
  wire \mul_b_reg[14] ;
  wire \mul_b_reg[15] ;
  wire \mul_b_reg[16] ;
  wire \mul_b_reg[17] ;
  wire \mul_b_reg[18] ;
  wire \mul_b_reg[19] ;
  wire \mul_b_reg[1] ;
  wire \mul_b_reg[20] ;
  wire \mul_b_reg[21] ;
  wire \mul_b_reg[22] ;
  wire \mul_b_reg[23] ;
  wire \mul_b_reg[24] ;
  wire \mul_b_reg[25] ;
  wire \mul_b_reg[26] ;
  wire \mul_b_reg[27] ;
  wire \mul_b_reg[28] ;
  wire \mul_b_reg[29] ;
  wire \mul_b_reg[2] ;
  wire \mul_b_reg[30] ;
  wire [1:0]\mul_b_reg[32] ;
  wire [1:0]\mul_b_reg[32]_0 ;
  wire \mul_b_reg[3] ;
  wire \mul_b_reg[5] ;
  wire \mul_b_reg[6] ;
  wire \mul_b_reg[7] ;
  wire \mul_b_reg[8] ;
  wire \mul_b_reg[9] ;
  wire mul_rslt;
  wire mul_rslt0;
  wire mul_rslt_reg;
  wire [15:0]mulh;
  wire \mulh_reg[0] ;
  wire [0:0]\niho_dsp_a[32]_INST_0_i_12 ;
  wire [0:0]niho_dsp_b;
  wire \niho_dsp_b[4] ;
  wire \niho_dsp_b[4]_0 ;
  wire [15:0]niho_dsp_c;
  wire \niho_dsp_c[31] ;
  wire [0:0]out;
  wire p_0_in;
  wire [30:0]\rem_reg[30] ;
  wire \remden_reg[12] ;
  wire \remden_reg[13] ;
  wire \remden_reg[14] ;
  wire \remden_reg[15] ;
  wire \remden_reg[16] ;
  wire \remden_reg[16]_0 ;
  wire \remden_reg[17] ;
  wire \remden_reg[17]_0 ;
  wire \remden_reg[18] ;
  wire \remden_reg[18]_0 ;
  wire \remden_reg[19] ;
  wire \remden_reg[19]_0 ;
  wire \remden_reg[20] ;
  wire \remden_reg[20]_0 ;
  wire \remden_reg[21] ;
  wire \remden_reg[21]_0 ;
  wire \remden_reg[22] ;
  wire \remden_reg[22]_0 ;
  wire \remden_reg[23] ;
  wire \remden_reg[23]_0 ;
  wire \remden_reg[24] ;
  wire \remden_reg[24]_0 ;
  wire \remden_reg[25] ;
  wire \remden_reg[25]_0 ;
  wire \remden_reg[26] ;
  wire \remden_reg[26]_0 ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire \tr[31]_i_5 ;
  wire \tr[31]_i_5_0 ;

  niho_alu_div div
       (.Q(Q),
        .abus_0(abus_0),
        .bbus_0(bbus_0[15:0]),
        .\bcmd[2]_INST_0_i_1 (\bcmd[2]_INST_0_i_1 ),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(crdy_0),
        .dctl_sign(dctl_sign),
        .dctl_sign_f(dctl_sign_f),
        .\dctl_stat_reg[2] (\dctl_stat_reg[2] ),
        .div_crdy_reg(div_crdy),
        .div_crdy_reg_0(div_crdy_reg),
        .div_crdy_reg_1(div_crdy_reg_0),
        .div_crdy_reg_2(div_crdy_reg_1),
        .\dso_reg[19] (\dso_reg[19] ),
        .\dso_reg[19]_0 (\dso_reg[19]_0 ),
        .\dso_reg[19]_1 (\dso_reg[19]_1 ),
        .\dso_reg[19]_2 (\dso_reg[19]_2 ),
        .\dso_reg[23] (\dso_reg[23] ),
        .\dso_reg[23]_0 (\dso_reg[23]_0 ),
        .\dso_reg[23]_1 (\dso_reg[23]_1 ),
        .\dso_reg[23]_2 (\dso_reg[23]_2 ),
        .\dso_reg[27] (\dso_reg[27] ),
        .\dso_reg[27]_0 (\dso_reg[27]_0 ),
        .\dso_reg[27]_1 (\dso_reg[27]_1 ),
        .\dso_reg[27]_2 (\dso_reg[27]_2 ),
        .\dso_reg[31] (\dso_reg[31] ),
        .\dso_reg[31]_0 (\dso_reg[31]_0 ),
        .\dso_reg[31]_1 (\dso_reg[31]_1 ),
        .\dso_reg[31]_2 (\dso_reg[31]_2 ),
        .\niho_dsp_a[32]_INST_0_i_12 (\niho_dsp_a[32]_INST_0_i_12 ),
        .niho_dsp_c(niho_dsp_c[15]),
        .\niho_dsp_c[31] (\niho_dsp_c[31] ),
        .out(out),
        .p_0_in(p_0_in),
        .\rem_reg[30] (\rem_reg[30] ),
        .\remden_reg[12] (\remden_reg[12] ),
        .\remden_reg[13] (\remden_reg[13] ),
        .\remden_reg[14] (\remden_reg[14] ),
        .\remden_reg[15] (\remden_reg[15] ),
        .\remden_reg[16] (\remden_reg[16] ),
        .\remden_reg[16]_0 (\remden_reg[16]_0 ),
        .\remden_reg[17] (\remden_reg[17] ),
        .\remden_reg[17]_0 (\remden_reg[17]_0 ),
        .\remden_reg[18] (\remden_reg[18] ),
        .\remden_reg[18]_0 (\remden_reg[18]_0 ),
        .\remden_reg[19] (\remden_reg[19] ),
        .\remden_reg[19]_0 (\remden_reg[19]_0 ),
        .\remden_reg[20] (\remden_reg[20] ),
        .\remden_reg[20]_0 (\remden_reg[20]_0 ),
        .\remden_reg[21] (\remden_reg[21] ),
        .\remden_reg[21]_0 (\remden_reg[21]_0 ),
        .\remden_reg[22] (\remden_reg[22] ),
        .\remden_reg[22]_0 (\remden_reg[22]_0 ),
        .\remden_reg[23] (\remden_reg[23] ),
        .\remden_reg[23]_0 (\remden_reg[23]_0 ),
        .\remden_reg[24] (\remden_reg[24] ),
        .\remden_reg[24]_0 (\remden_reg[24]_0 ),
        .\remden_reg[25] (\remden_reg[25] ),
        .\remden_reg[25]_0 (\remden_reg[25]_0 ),
        .\remden_reg[26] (\remden_reg[26] ),
        .\remden_reg[26]_0 (\remden_reg[26]_0 ),
        .\remden_reg[27] (\remden_reg[27] ),
        .\remden_reg[28] (\remden_reg[28] ),
        .\remden_reg[29] (\remden_reg[29] ),
        .\remden_reg[30] (\remden_reg[30] ),
        .\remden_reg[31] (\remden_reg[31] ),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .\tr[31]_i_5 (mul_rslt_reg),
        .\tr[31]_i_5_0 (\tr[31]_i_5 ),
        .\tr[31]_i_5_1 (\tr[31]_i_5_0 ));
  niho_alu_mul mul
       (.D(D),
        .abus_0(abus_0),
        .bbus_0(bbus_0),
        .clk(clk),
        .mul_a(mul_a),
        .mul_a_i(mul_a_i),
        .\mul_a_reg[16]_0 (\mul_a_reg[16] ),
        .mul_b(mul_b),
        .\mul_b_reg[0]_0 (\mul_b_reg[0] ),
        .\mul_b_reg[0]_1 (\mul_b_reg[0]_0 ),
        .\mul_b_reg[10]_0 (\mul_b_reg[10] ),
        .\mul_b_reg[11]_0 (\mul_b_reg[11] ),
        .\mul_b_reg[12]_0 (\mul_b_reg[12] ),
        .\mul_b_reg[13]_0 (\mul_b_reg[13] ),
        .\mul_b_reg[14]_0 (\mul_b_reg[14] ),
        .\mul_b_reg[15]_0 (\mul_b_reg[15] ),
        .\mul_b_reg[16]_0 (\mul_b_reg[16] ),
        .\mul_b_reg[17]_0 (\mul_b_reg[17] ),
        .\mul_b_reg[18]_0 (\mul_b_reg[18] ),
        .\mul_b_reg[19]_0 (\mul_b_reg[19] ),
        .\mul_b_reg[1]_0 (\mul_b_reg[1] ),
        .\mul_b_reg[20]_0 (\mul_b_reg[20] ),
        .\mul_b_reg[21]_0 (\mul_b_reg[21] ),
        .\mul_b_reg[22]_0 (\mul_b_reg[22] ),
        .\mul_b_reg[23]_0 (\mul_b_reg[23] ),
        .\mul_b_reg[24]_0 (\mul_b_reg[24] ),
        .\mul_b_reg[25]_0 (\mul_b_reg[25] ),
        .\mul_b_reg[26]_0 (\mul_b_reg[26] ),
        .\mul_b_reg[27]_0 (\mul_b_reg[27] ),
        .\mul_b_reg[28]_0 (\mul_b_reg[28] ),
        .\mul_b_reg[29]_0 (\mul_b_reg[29] ),
        .\mul_b_reg[2]_0 (\mul_b_reg[2] ),
        .\mul_b_reg[30]_0 (\mul_b_reg[30] ),
        .\mul_b_reg[32]_0 (\mul_b_reg[32] ),
        .\mul_b_reg[32]_1 (\mul_b_reg[32]_0 ),
        .\mul_b_reg[3]_0 (\mul_b_reg[3] ),
        .\mul_b_reg[5]_0 (\mul_b_reg[5] ),
        .\mul_b_reg[6]_0 (\mul_b_reg[6] ),
        .\mul_b_reg[7]_0 (\mul_b_reg[7] ),
        .\mul_b_reg[8]_0 (\mul_b_reg[8] ),
        .\mul_b_reg[9]_0 (\mul_b_reg[9] ),
        .mul_rslt(mul_rslt),
        .mul_rslt0(mul_rslt0),
        .mul_rslt_reg_0(mul_rslt_reg),
        .mulh(mulh),
        .\mulh_reg[0]_0 (\mulh_reg[0] ),
        .niho_dsp_b(niho_dsp_b),
        .\niho_dsp_b[4] (\niho_dsp_b[4] ),
        .\niho_dsp_b[4]_0 (\niho_dsp_b[4]_0 ),
        .niho_dsp_c(niho_dsp_c),
        .p_0_in(p_0_in),
        .rgf_sr_nh(rgf_sr_nh));
endmodule

module niho_alu_div
   (dctl_sign_f,
    div_crdy_reg,
    div_crdy_reg_0,
    \niho_dsp_c[31] ,
    Q,
    \remden_reg[13] ,
    \remden_reg[15] ,
    \remden_reg[22] ,
    \remden_reg[23] ,
    \remden_reg[24] ,
    \remden_reg[26] ,
    \remden_reg[25] ,
    \remden_reg[21] ,
    \remden_reg[20] ,
    \remden_reg[19] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] ,
    \remden_reg[12] ,
    \rem_reg[30] ,
    \remden_reg[14] ,
    div_crdy_reg_1,
    crdy_0,
    div_crdy_reg_2,
    p_0_in,
    clk,
    dctl_sign,
    abus_0,
    rgf_sr_nh,
    \tr[31]_i_5 ,
    niho_dsp_c,
    \tr[31]_i_5_0 ,
    \tr[31]_i_5_1 ,
    \dctl_stat_reg[2] ,
    crdy,
    \bcmd[2]_INST_0_i_1 ,
    rst_n,
    out,
    \niho_dsp_a[32]_INST_0_i_12 ,
    \dso_reg[19] ,
    \dso_reg[19]_0 ,
    \dso_reg[19]_1 ,
    \dso_reg[19]_2 ,
    \dso_reg[23] ,
    \dso_reg[23]_0 ,
    \dso_reg[23]_1 ,
    \dso_reg[23]_2 ,
    \dso_reg[27] ,
    \dso_reg[27]_0 ,
    \dso_reg[27]_1 ,
    \dso_reg[27]_2 ,
    \dso_reg[31] ,
    \dso_reg[31]_0 ,
    \dso_reg[31]_1 ,
    \dso_reg[31]_2 ,
    \remden_reg[31] ,
    \remden_reg[29] ,
    \remden_reg[25]_0 ,
    \remden_reg[24]_0 ,
    \remden_reg[23]_0 ,
    \remden_reg[22]_0 ,
    \remden_reg[21]_0 ,
    \remden_reg[20]_0 ,
    \remden_reg[18]_0 ,
    \remden_reg[17]_0 ,
    \remden_reg[16]_0 ,
    \remden_reg[30] ,
    \remden_reg[19]_0 ,
    \remden_reg[28] ,
    \remden_reg[27] ,
    \remden_reg[26]_0 ,
    bbus_0);
  output dctl_sign_f;
  output div_crdy_reg;
  output div_crdy_reg_0;
  output \niho_dsp_c[31] ;
  output [30:0]Q;
  output \remden_reg[13] ;
  output \remden_reg[15] ;
  output \remden_reg[22] ;
  output \remden_reg[23] ;
  output \remden_reg[24] ;
  output \remden_reg[26] ;
  output \remden_reg[25] ;
  output \remden_reg[21] ;
  output \remden_reg[20] ;
  output \remden_reg[19] ;
  output \remden_reg[18] ;
  output \remden_reg[17] ;
  output \remden_reg[16] ;
  output \remden_reg[12] ;
  output [30:0]\rem_reg[30] ;
  output \remden_reg[14] ;
  output div_crdy_reg_1;
  output crdy_0;
  output div_crdy_reg_2;
  input p_0_in;
  input clk;
  input dctl_sign;
  input [15:0]abus_0;
  input rgf_sr_nh;
  input \tr[31]_i_5 ;
  input [0:0]niho_dsp_c;
  input \tr[31]_i_5_0 ;
  input \tr[31]_i_5_1 ;
  input \dctl_stat_reg[2] ;
  input crdy;
  input \bcmd[2]_INST_0_i_1 ;
  input rst_n;
  input [0:0]out;
  input [0:0]\niho_dsp_a[32]_INST_0_i_12 ;
  input \dso_reg[19] ;
  input \dso_reg[19]_0 ;
  input \dso_reg[19]_1 ;
  input \dso_reg[19]_2 ;
  input \dso_reg[23] ;
  input \dso_reg[23]_0 ;
  input \dso_reg[23]_1 ;
  input \dso_reg[23]_2 ;
  input \dso_reg[27] ;
  input \dso_reg[27]_0 ;
  input \dso_reg[27]_1 ;
  input \dso_reg[27]_2 ;
  input \dso_reg[31] ;
  input \dso_reg[31]_0 ;
  input \dso_reg[31]_1 ;
  input \dso_reg[31]_2 ;
  input \remden_reg[31] ;
  input \remden_reg[29] ;
  input \remden_reg[25]_0 ;
  input \remden_reg[24]_0 ;
  input \remden_reg[23]_0 ;
  input \remden_reg[22]_0 ;
  input \remden_reg[21]_0 ;
  input \remden_reg[20]_0 ;
  input \remden_reg[18]_0 ;
  input \remden_reg[17]_0 ;
  input \remden_reg[16]_0 ;
  input \remden_reg[30] ;
  input \remden_reg[19]_0 ;
  input \remden_reg[28] ;
  input \remden_reg[27] ;
  input \remden_reg[26]_0 ;
  input [15:0]bbus_0;

  wire [30:0]Q;
  wire [15:0]abus_0;
  wire [31:0]add_out;
  wire [15:0]bbus_0;
  wire \bcmd[2]_INST_0_i_1 ;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire dadd_n_51;
  wire dadd_n_52;
  wire dadd_n_53;
  wire dadd_n_54;
  wire dadd_n_55;
  wire dadd_n_56;
  wire dadd_n_57;
  wire dadd_n_58;
  wire dadd_n_59;
  wire dctl_long_f;
  wire dctl_n_10;
  wire dctl_n_100;
  wire dctl_n_101;
  wire dctl_n_102;
  wire dctl_n_103;
  wire dctl_n_104;
  wire dctl_n_105;
  wire dctl_n_106;
  wire dctl_n_107;
  wire dctl_n_108;
  wire dctl_n_109;
  wire dctl_n_11;
  wire dctl_n_110;
  wire dctl_n_111;
  wire dctl_n_112;
  wire dctl_n_113;
  wire dctl_n_114;
  wire dctl_n_115;
  wire dctl_n_116;
  wire dctl_n_117;
  wire dctl_n_118;
  wire dctl_n_119;
  wire dctl_n_12;
  wire dctl_n_120;
  wire dctl_n_121;
  wire dctl_n_122;
  wire dctl_n_123;
  wire dctl_n_124;
  wire dctl_n_125;
  wire dctl_n_126;
  wire dctl_n_127;
  wire dctl_n_128;
  wire dctl_n_129;
  wire dctl_n_13;
  wire dctl_n_130;
  wire dctl_n_131;
  wire dctl_n_132;
  wire dctl_n_133;
  wire dctl_n_134;
  wire dctl_n_135;
  wire dctl_n_136;
  wire dctl_n_137;
  wire dctl_n_138;
  wire dctl_n_139;
  wire dctl_n_14;
  wire dctl_n_140;
  wire dctl_n_141;
  wire dctl_n_142;
  wire dctl_n_143;
  wire dctl_n_144;
  wire dctl_n_145;
  wire dctl_n_146;
  wire dctl_n_147;
  wire dctl_n_148;
  wire dctl_n_149;
  wire dctl_n_15;
  wire dctl_n_150;
  wire dctl_n_151;
  wire dctl_n_152;
  wire dctl_n_153;
  wire dctl_n_154;
  wire dctl_n_155;
  wire dctl_n_156;
  wire dctl_n_157;
  wire dctl_n_158;
  wire dctl_n_159;
  wire dctl_n_16;
  wire dctl_n_160;
  wire dctl_n_161;
  wire dctl_n_162;
  wire dctl_n_163;
  wire dctl_n_164;
  wire dctl_n_165;
  wire dctl_n_166;
  wire dctl_n_167;
  wire dctl_n_168;
  wire dctl_n_169;
  wire dctl_n_17;
  wire dctl_n_170;
  wire dctl_n_171;
  wire dctl_n_172;
  wire dctl_n_173;
  wire dctl_n_174;
  wire dctl_n_175;
  wire dctl_n_176;
  wire dctl_n_177;
  wire dctl_n_178;
  wire dctl_n_179;
  wire dctl_n_18;
  wire dctl_n_180;
  wire dctl_n_181;
  wire dctl_n_182;
  wire dctl_n_183;
  wire dctl_n_184;
  wire dctl_n_185;
  wire dctl_n_186;
  wire dctl_n_187;
  wire dctl_n_188;
  wire dctl_n_189;
  wire dctl_n_19;
  wire dctl_n_190;
  wire dctl_n_191;
  wire dctl_n_192;
  wire dctl_n_193;
  wire dctl_n_194;
  wire dctl_n_195;
  wire dctl_n_196;
  wire dctl_n_197;
  wire dctl_n_24;
  wire dctl_n_25;
  wire dctl_n_26;
  wire dctl_n_27;
  wire dctl_n_28;
  wire dctl_n_29;
  wire dctl_n_3;
  wire dctl_n_30;
  wire dctl_n_31;
  wire dctl_n_32;
  wire dctl_n_33;
  wire dctl_n_34;
  wire dctl_n_35;
  wire dctl_n_36;
  wire dctl_n_37;
  wire dctl_n_4;
  wire dctl_n_40;
  wire dctl_n_42;
  wire dctl_n_43;
  wire dctl_n_44;
  wire dctl_n_45;
  wire dctl_n_46;
  wire dctl_n_47;
  wire dctl_n_48;
  wire dctl_n_49;
  wire dctl_n_50;
  wire dctl_n_51;
  wire dctl_n_52;
  wire dctl_n_53;
  wire dctl_n_54;
  wire dctl_n_55;
  wire dctl_n_56;
  wire dctl_n_57;
  wire dctl_n_58;
  wire dctl_n_59;
  wire dctl_n_6;
  wire dctl_n_60;
  wire dctl_n_61;
  wire dctl_n_62;
  wire dctl_n_63;
  wire dctl_n_64;
  wire dctl_n_65;
  wire dctl_n_66;
  wire dctl_n_67;
  wire dctl_n_68;
  wire dctl_n_69;
  wire dctl_n_7;
  wire dctl_n_70;
  wire dctl_n_71;
  wire dctl_n_72;
  wire dctl_n_73;
  wire dctl_n_74;
  wire dctl_n_75;
  wire dctl_n_76;
  wire dctl_n_77;
  wire dctl_n_78;
  wire dctl_n_79;
  wire dctl_n_8;
  wire dctl_n_80;
  wire dctl_n_81;
  wire dctl_n_82;
  wire dctl_n_83;
  wire dctl_n_84;
  wire dctl_n_85;
  wire dctl_n_86;
  wire dctl_n_87;
  wire dctl_n_88;
  wire dctl_n_89;
  wire dctl_n_9;
  wire dctl_n_90;
  wire dctl_n_91;
  wire dctl_n_92;
  wire dctl_n_93;
  wire dctl_n_94;
  wire dctl_n_95;
  wire dctl_n_96;
  wire dctl_n_97;
  wire dctl_n_98;
  wire dctl_n_99;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[2] ;
  wire [3:3]den2;
  wire div_crdy_reg;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire div_crdy_reg_2;
  wire [31:0]dso_0;
  wire \dso_reg[19] ;
  wire \dso_reg[19]_0 ;
  wire \dso_reg[19]_1 ;
  wire \dso_reg[19]_2 ;
  wire \dso_reg[23] ;
  wire \dso_reg[23]_0 ;
  wire \dso_reg[23]_1 ;
  wire \dso_reg[23]_2 ;
  wire \dso_reg[27] ;
  wire \dso_reg[27]_0 ;
  wire \dso_reg[27]_1 ;
  wire \dso_reg[27]_2 ;
  wire \dso_reg[31] ;
  wire \dso_reg[31]_0 ;
  wire \dso_reg[31]_1 ;
  wire \dso_reg[31]_2 ;
  wire [31:0]fdiv_rem;
  wire \fsm/chg_rem_sgn0 ;
  wire [0:0]\niho_dsp_a[32]_INST_0_i_12 ;
  wire [0:0]niho_dsp_c;
  wire \niho_dsp_c[31] ;
  wire [0:0]out;
  wire p_0_in;
  wire p_0_in0;
  wire [0:0]p_1_in5_in;
  wire [31:0]p_2_in;
  wire [31:31]quo;
  wire rden_n_1;
  wire rden_n_10;
  wire rden_n_11;
  wire rden_n_12;
  wire rden_n_13;
  wire rden_n_14;
  wire rden_n_15;
  wire rden_n_16;
  wire rden_n_17;
  wire rden_n_18;
  wire rden_n_19;
  wire rden_n_2;
  wire rden_n_20;
  wire rden_n_21;
  wire rden_n_22;
  wire rden_n_23;
  wire rden_n_24;
  wire rden_n_25;
  wire rden_n_26;
  wire rden_n_27;
  wire rden_n_28;
  wire rden_n_29;
  wire rden_n_3;
  wire rden_n_30;
  wire rden_n_31;
  wire rden_n_32;
  wire rden_n_33;
  wire rden_n_34;
  wire rden_n_35;
  wire rden_n_36;
  wire rden_n_37;
  wire rden_n_38;
  wire rden_n_39;
  wire rden_n_40;
  wire rden_n_41;
  wire rden_n_42;
  wire rden_n_43;
  wire rden_n_44;
  wire rden_n_45;
  wire rden_n_46;
  wire rden_n_47;
  wire rden_n_48;
  wire rden_n_49;
  wire rden_n_50;
  wire rden_n_51;
  wire rden_n_52;
  wire rden_n_53;
  wire rden_n_54;
  wire rden_n_55;
  wire rden_n_56;
  wire rden_n_57;
  wire rden_n_58;
  wire rden_n_59;
  wire rden_n_6;
  wire rden_n_60;
  wire rden_n_61;
  wire rden_n_62;
  wire rden_n_63;
  wire rden_n_64;
  wire rden_n_65;
  wire rden_n_66;
  wire rden_n_67;
  wire rden_n_68;
  wire rden_n_69;
  wire rden_n_7;
  wire rden_n_70;
  wire rden_n_71;
  wire rden_n_72;
  wire rden_n_8;
  wire rden_n_86;
  wire rden_n_87;
  wire rden_n_88;
  wire rden_n_89;
  wire rden_n_9;
  wire rden_n_90;
  wire rden_n_91;
  wire rden_n_92;
  wire rden_n_93;
  wire rden_n_95;
  wire rden_n_96;
  wire rden_n_97;
  wire rden_n_98;
  wire rden_n_99;
  wire rdso_n_0;
  wire rdso_n_1;
  wire [31:31]rem;
  wire [33:33]rem1;
  wire [33:33]rem2;
  wire [33:33]rem3;
  wire [30:0]\rem_reg[30] ;
  wire \remden_reg[12] ;
  wire \remden_reg[13] ;
  wire \remden_reg[14] ;
  wire \remden_reg[15] ;
  wire \remden_reg[16] ;
  wire \remden_reg[16]_0 ;
  wire \remden_reg[17] ;
  wire \remden_reg[17]_0 ;
  wire \remden_reg[18] ;
  wire \remden_reg[18]_0 ;
  wire \remden_reg[19] ;
  wire \remden_reg[19]_0 ;
  wire \remden_reg[20] ;
  wire \remden_reg[20]_0 ;
  wire \remden_reg[21] ;
  wire \remden_reg[21]_0 ;
  wire \remden_reg[22] ;
  wire \remden_reg[22]_0 ;
  wire \remden_reg[23] ;
  wire \remden_reg[23]_0 ;
  wire \remden_reg[24] ;
  wire \remden_reg[24]_0 ;
  wire \remden_reg[25] ;
  wire \remden_reg[25]_0 ;
  wire \remden_reg[26] ;
  wire \remden_reg[26]_0 ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire \tr[31]_i_5 ;
  wire \tr[31]_i_5_0 ;
  wire \tr[31]_i_5_1 ;

  niho_div_add dadd
       (.D(p_2_in[27:0]),
        .DI({dctl_n_26,dctl_n_27,dctl_n_28,dctl_n_29}),
        .O(rem3),
        .Q(Q[23:0]),
        .S({dctl_n_34,dctl_n_35,dctl_n_36,dctl_n_37}),
        .\quo_reg[0] (p_0_in0),
        .\quo_reg[11] ({dctl_n_61,dctl_n_62,dctl_n_63,dctl_n_64}),
        .\quo_reg[11]_0 ({dctl_n_85,dctl_n_86,dctl_n_87,dctl_n_88}),
        .\quo_reg[15] ({dctl_n_57,dctl_n_58,dctl_n_59,dctl_n_60}),
        .\quo_reg[15]_0 ({dctl_n_81,dctl_n_82,dctl_n_83,dctl_n_84}),
        .\quo_reg[19] ({dctl_n_53,dctl_n_54,dctl_n_55,dctl_n_56}),
        .\quo_reg[19]_0 ({dctl_n_77,dctl_n_78,dctl_n_79,dctl_n_80}),
        .\quo_reg[1] (rem1),
        .\quo_reg[27] ({dctl_n_45,dctl_n_46,dctl_n_47,dctl_n_48}),
        .\quo_reg[27]_0 ({dctl_n_69,dctl_n_70,dctl_n_71,dctl_n_72}),
        .\quo_reg[27]_1 (dctl_n_17),
        .\quo_reg[2] (rem2),
        .\quo_reg[7] ({dctl_n_65,dctl_n_66,dctl_n_67,dctl_n_68}),
        .\quo_reg[7]_0 ({dctl_n_89,dctl_n_90,dctl_n_91,dctl_n_92}),
        .\rem_reg[30] ({add_out[31:26],add_out[19],add_out[15:0]}),
        .\remden_reg[16] (\remden_reg[16]_0 ),
        .\remden_reg[17] (\remden_reg[17]_0 ),
        .\remden_reg[18] (\remden_reg[18]_0 ),
        .\remden_reg[20] (\remden_reg[20]_0 ),
        .\remden_reg[21] (\remden_reg[21]_0 ),
        .\remden_reg[22] (\remden_reg[22]_0 ),
        .\remden_reg[23] ({dctl_n_49,dctl_n_50,dctl_n_51,dctl_n_52}),
        .\remden_reg[23]_0 ({dctl_n_73,dctl_n_74,dctl_n_75,dctl_n_76}),
        .\remden_reg[23]_1 (\remden_reg[23]_0 ),
        .\remden_reg[24] (\remden_reg[24]_0 ),
        .\remden_reg[25] (dctl_n_4),
        .\remden_reg[25]_0 (\remden_reg[25]_0 ),
        .\remden_reg[31] ({dctl_n_42,dctl_n_43,dctl_n_44}),
        .\remden_reg[31]_0 ({dctl_n_30,dctl_n_31,dctl_n_32,dctl_n_33}),
        .rst_n(rst_n),
        .rst_n_0(dadd_n_51),
        .rst_n_1(dadd_n_52),
        .rst_n_2(dadd_n_53),
        .rst_n_3(dadd_n_54),
        .rst_n_4(dadd_n_55),
        .rst_n_5(dadd_n_56),
        .rst_n_6(dadd_n_57),
        .rst_n_7(dadd_n_58),
        .rst_n_8(dadd_n_59));
  niho_div_ctl dctl
       (.D(p_2_in[31:28]),
        .DI(rden_n_67),
        .E(dctl_n_19),
        .Q({quo,Q}),
        .S({dctl_n_34,dctl_n_35,dctl_n_36,dctl_n_37}),
        .abus_0(abus_0),
        .add_out0_carry__2_i_10(\remden_reg[14] ),
        .add_out0_carry__2_i_11(\remden_reg[13] ),
        .add_out0_carry__2_i_12(\remden_reg[12] ),
        .add_out0_carry__2_i_9(\remden_reg[15] ),
        .add_out0_carry__3_i_10(\remden_reg[18] ),
        .add_out0_carry__3_i_11(\remden_reg[17] ),
        .add_out0_carry__3_i_12(\remden_reg[16] ),
        .add_out0_carry__3_i_9(\remden_reg[19] ),
        .add_out0_carry__4_i_10(\remden_reg[22] ),
        .add_out0_carry__4_i_11(\remden_reg[21] ),
        .add_out0_carry__4_i_12(\remden_reg[20] ),
        .add_out0_carry__4_i_9(\remden_reg[23] ),
        .add_out0_carry__5_i_10(\remden_reg[26] ),
        .add_out0_carry__5_i_11(\remden_reg[25] ),
        .add_out0_carry__5_i_12(\remden_reg[24] ),
        .add_out0_carry__6(dso_0),
        .add_out0_carry__6_i_10(rden_n_71),
        .add_out0_carry__6_i_9(rden_n_69),
        .bbus_0(bbus_0),
        .\bcmd[2]_INST_0_i_1 (\bcmd[2]_INST_0_i_1 ),
        .chg_quo_sgn_reg(rdso_n_1),
        .chg_rem_sgn0(\fsm/chg_rem_sgn0 ),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(crdy_0),
        .dctl_long_f(dctl_long_f),
        .dctl_sign(dctl_sign),
        .dctl_sign_f(dctl_sign_f),
        .\dctl_stat_reg[1] (dctl_n_18),
        .\dctl_stat_reg[2] (dctl_n_17),
        .\dctl_stat_reg[2]_0 (dctl_n_25),
        .\dctl_stat_reg[2]_1 (\dctl_stat_reg[2] ),
        .\dctl_stat_reg[3] (dctl_n_4),
        .\dctl_stat_reg[3]_0 (rdso_n_0),
        .den2(den2),
        .div_crdy_reg_0(div_crdy_reg),
        .div_crdy_reg_1(div_crdy_reg_0),
        .div_crdy_reg_2(dctl_n_24),
        .div_crdy_reg_3(div_crdy_reg_1),
        .div_crdy_reg_4(div_crdy_reg_2),
        .\dso_reg[19] (\dso_reg[19] ),
        .\dso_reg[19]_0 (\dso_reg[19]_0 ),
        .\dso_reg[19]_1 (\dso_reg[19]_1 ),
        .\dso_reg[19]_2 (\dso_reg[19]_2 ),
        .\dso_reg[23] (\dso_reg[23] ),
        .\dso_reg[23]_0 (\dso_reg[23]_0 ),
        .\dso_reg[23]_1 (\dso_reg[23]_1 ),
        .\dso_reg[23]_2 (\dso_reg[23]_2 ),
        .\dso_reg[27] (\dso_reg[27] ),
        .\dso_reg[27]_0 (\dso_reg[27]_0 ),
        .\dso_reg[27]_1 (\dso_reg[27]_1 ),
        .\dso_reg[27]_2 (\dso_reg[27]_2 ),
        .\dso_reg[31] ({dctl_n_30,dctl_n_31,dctl_n_32,dctl_n_33}),
        .\dso_reg[31]_0 (\dso_reg[31] ),
        .\dso_reg[31]_1 (\dso_reg[31]_0 ),
        .\dso_reg[31]_2 (\dso_reg[31]_1 ),
        .\dso_reg[31]_3 (\dso_reg[31]_2 ),
        .fdiv_rem(fdiv_rem),
        .fdiv_rem_msb_f_reg(p_0_in0),
        .\niho_dsp_a[32]_INST_0_i_12 (\niho_dsp_a[32]_INST_0_i_12 ),
        .out(out),
        .p_0_in(p_0_in),
        .\rem_reg[11] ({dctl_n_61,dctl_n_62,dctl_n_63,dctl_n_64}),
        .\rem_reg[11]_0 ({dctl_n_85,dctl_n_86,dctl_n_87,dctl_n_88}),
        .\rem_reg[15] ({dctl_n_57,dctl_n_58,dctl_n_59,dctl_n_60}),
        .\rem_reg[15]_0 ({dctl_n_81,dctl_n_82,dctl_n_83,dctl_n_84}),
        .\rem_reg[19] ({dctl_n_53,dctl_n_54,dctl_n_55,dctl_n_56}),
        .\rem_reg[19]_0 ({dctl_n_77,dctl_n_78,dctl_n_79,dctl_n_80}),
        .\rem_reg[23] ({dctl_n_49,dctl_n_50,dctl_n_51,dctl_n_52}),
        .\rem_reg[23]_0 ({dctl_n_73,dctl_n_74,dctl_n_75,dctl_n_76}),
        .\rem_reg[27] ({dctl_n_45,dctl_n_46,dctl_n_47,dctl_n_48}),
        .\rem_reg[27]_0 ({dctl_n_69,dctl_n_70,dctl_n_71,dctl_n_72}),
        .\rem_reg[30] ({dctl_n_42,dctl_n_43,dctl_n_44}),
        .\rem_reg[31] ({dctl_n_134,dctl_n_135,dctl_n_136,dctl_n_137,dctl_n_138,dctl_n_139,dctl_n_140,dctl_n_141,dctl_n_142,dctl_n_143,dctl_n_144,dctl_n_145,dctl_n_146,dctl_n_147,dctl_n_148,dctl_n_149,dctl_n_150,dctl_n_151,dctl_n_152,dctl_n_153,dctl_n_154,dctl_n_155,dctl_n_156,dctl_n_157,dctl_n_158,dctl_n_159,dctl_n_160,dctl_n_161,dctl_n_162,dctl_n_163,dctl_n_164,dctl_n_165}),
        .\rem_reg[31]_0 ({rem,\rem_reg[30] }),
        .\rem_reg[3] ({dctl_n_26,dctl_n_27,dctl_n_28,dctl_n_29}),
        .\rem_reg[7] ({dctl_n_65,dctl_n_66,dctl_n_67,dctl_n_68}),
        .\rem_reg[7]_0 ({dctl_n_89,dctl_n_90,dctl_n_91,dctl_n_92}),
        .\remden_reg[10] (rden_n_91),
        .\remden_reg[11] (rden_n_90),
        .\remden_reg[12] (rden_n_89),
        .\remden_reg[13] (rden_n_88),
        .\remden_reg[14] (rden_n_87),
        .\remden_reg[15] (rden_n_86),
        .\remden_reg[19] (\remden_reg[19]_0 ),
        .\remden_reg[28] (dctl_n_122),
        .\remden_reg[28]_0 (dctl_n_123),
        .\remden_reg[28]_1 (dctl_n_124),
        .\remden_reg[28]_2 (dctl_n_125),
        .\remden_reg[29] (\remden_reg[29] ),
        .\remden_reg[30] (\remden_reg[30] ),
        .\remden_reg[31] ({add_out[31:28],add_out[19],add_out[15:0]}),
        .\remden_reg[31]_0 (rden_n_99),
        .\remden_reg[31]_1 (\remden_reg[31] ),
        .\remden_reg[4] (rden_n_98),
        .\remden_reg[5] (rden_n_97),
        .\remden_reg[6] (rden_n_96),
        .\remden_reg[7] (rden_n_95),
        .\remden_reg[8] (rden_n_93),
        .\remden_reg[9] (rden_n_92),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .rst_n_0(dctl_n_40),
        .rst_n_1(dctl_n_93),
        .rst_n_10(dctl_n_102),
        .rst_n_11(dctl_n_103),
        .rst_n_12(dctl_n_104),
        .rst_n_13(dctl_n_105),
        .rst_n_14(dctl_n_106),
        .rst_n_15(dctl_n_107),
        .rst_n_16(dctl_n_108),
        .rst_n_17(dctl_n_109),
        .rst_n_18(dctl_n_110),
        .rst_n_19(dctl_n_111),
        .rst_n_2(dctl_n_94),
        .rst_n_20(dctl_n_112),
        .rst_n_21(dctl_n_113),
        .rst_n_22(dctl_n_114),
        .rst_n_23(dctl_n_115),
        .rst_n_24(dctl_n_116),
        .rst_n_25(dctl_n_117),
        .rst_n_26(dctl_n_118),
        .rst_n_27(dctl_n_119),
        .rst_n_28(dctl_n_120),
        .rst_n_29(dctl_n_121),
        .rst_n_3(dctl_n_95),
        .rst_n_30(dctl_n_126),
        .rst_n_31(dctl_n_127),
        .rst_n_32(dctl_n_128),
        .rst_n_33(dctl_n_129),
        .rst_n_34(dctl_n_130),
        .rst_n_35(dctl_n_131),
        .rst_n_36(dctl_n_132),
        .rst_n_37(dctl_n_133),
        .rst_n_4(dctl_n_96),
        .rst_n_5(dctl_n_97),
        .rst_n_6(dctl_n_98),
        .rst_n_7(dctl_n_99),
        .rst_n_8(dctl_n_100),
        .rst_n_9(dctl_n_101),
        .\sr_reg[8] (dctl_n_3),
        .\sr_reg[8]_0 (dctl_n_6),
        .\sr_reg[8]_1 (dctl_n_7),
        .\sr_reg[8]_10 (dctl_n_16),
        .\sr_reg[8]_11 ({dctl_n_166,dctl_n_167,dctl_n_168,dctl_n_169,dctl_n_170,dctl_n_171,dctl_n_172,dctl_n_173,dctl_n_174,dctl_n_175,dctl_n_176,dctl_n_177,dctl_n_178,dctl_n_179,dctl_n_180,dctl_n_181,dctl_n_182,dctl_n_183,dctl_n_184,dctl_n_185,dctl_n_186,dctl_n_187,dctl_n_188,dctl_n_189,dctl_n_190,dctl_n_191,dctl_n_192,dctl_n_193,dctl_n_194,dctl_n_195,dctl_n_196,dctl_n_197}),
        .\sr_reg[8]_2 (dctl_n_8),
        .\sr_reg[8]_3 (dctl_n_9),
        .\sr_reg[8]_4 (dctl_n_10),
        .\sr_reg[8]_5 (dctl_n_11),
        .\sr_reg[8]_6 (dctl_n_12),
        .\sr_reg[8]_7 (dctl_n_13),
        .\sr_reg[8]_8 (dctl_n_14),
        .\sr_reg[8]_9 (dctl_n_15));
  niho_div_fdiv fdiv
       (.DI({rden_n_1,rden_n_2,rden_n_3,den2}),
        .O(rem3),
        .Q(dso_0[31:1]),
        .S({rden_n_6,rden_n_7,rden_n_8,rden_n_9}),
        .fdiv_rem(fdiv_rem),
        .p_1_in5_in(p_1_in5_in),
        .\quo_reg[3] (rden_n_72),
        .rem0_carry_0(rden_n_69),
        .rem0_carry_1(rden_n_68),
        .rem0_carry__7_i_1_0(p_0_in0),
        .rem1_carry_0(rden_n_67),
        .rem1_carry_1(rden_n_66),
        .rem1_carry__7_i_1_0(rem1),
        .rem2_carry__0_0({rden_n_14,rden_n_15,rden_n_16,rden_n_17}),
        .rem2_carry__0_1({rden_n_10,rden_n_11,rden_n_12,rden_n_13}),
        .rem2_carry__1_0({rden_n_22,rden_n_23,rden_n_24,rden_n_25}),
        .rem2_carry__1_1({rden_n_18,rden_n_19,rden_n_20,rden_n_21}),
        .rem2_carry__2_0({rden_n_30,rden_n_31,rden_n_32,rden_n_33}),
        .rem2_carry__2_1({rden_n_26,rden_n_27,rden_n_28,rden_n_29}),
        .rem2_carry__3_0({rden_n_38,rden_n_39,rden_n_40,rden_n_41}),
        .rem2_carry__3_1({rden_n_34,rden_n_35,rden_n_36,rden_n_37}),
        .rem2_carry__4_0({rden_n_46,rden_n_47,rden_n_48,rden_n_49}),
        .rem2_carry__4_1({rden_n_42,rden_n_43,rden_n_44,rden_n_45}),
        .rem2_carry__5_0({rden_n_54,rden_n_55,rden_n_56,rden_n_57}),
        .rem2_carry__5_1({rden_n_50,rden_n_51,rden_n_52,rden_n_53}),
        .rem2_carry__6_0({rden_n_62,rden_n_63,rden_n_64,rden_n_65}),
        .rem2_carry__6_1({rden_n_58,rden_n_59,rden_n_60,rden_n_61}),
        .rem2_carry__7_i_1_0(rem2),
        .\remden_reg[35] (rden_n_71),
        .\remden_reg[35]_0 (rden_n_70));
  niho_div_reg_den rden
       (.DI({rden_n_1,rden_n_2,rden_n_3,den2}),
        .O(rem3),
        .Q(dso_0),
        .S({rden_n_6,rden_n_7,rden_n_8,rden_n_9}),
        .chg_rem_sgn0(\fsm/chg_rem_sgn0 ),
        .clk(clk),
        .dctl_sign(dctl_sign),
        .p_1_in5_in(p_1_in5_in),
        .rem0_carry(rem1),
        .rem1_carry(rem2),
        .\remden_reg[0]_0 (rden_n_98),
        .\remden_reg[0]_1 (dctl_n_133),
        .\remden_reg[10]_0 (rden_n_87),
        .\remden_reg[10]_1 (dctl_n_10),
        .\remden_reg[11]_0 (rden_n_86),
        .\remden_reg[11]_1 (dctl_n_9),
        .\remden_reg[12]_0 (\remden_reg[12] ),
        .\remden_reg[12]_1 (dctl_n_8),
        .\remden_reg[13]_0 (\remden_reg[13] ),
        .\remden_reg[13]_1 (dctl_n_7),
        .\remden_reg[14]_0 (\remden_reg[14] ),
        .\remden_reg[14]_1 (dctl_n_6),
        .\remden_reg[15]_0 (\remden_reg[15] ),
        .\remden_reg[15]_1 (dctl_n_3),
        .\remden_reg[16]_0 (\remden_reg[16] ),
        .\remden_reg[16]_1 (dadd_n_59),
        .\remden_reg[17]_0 (\remden_reg[17] ),
        .\remden_reg[17]_1 (dadd_n_58),
        .\remden_reg[18]_0 (\remden_reg[18] ),
        .\remden_reg[18]_1 (dadd_n_57),
        .\remden_reg[19]_0 (\remden_reg[19] ),
        .\remden_reg[19]_1 (dctl_n_129),
        .\remden_reg[1]_0 (rden_n_97),
        .\remden_reg[1]_1 (dctl_n_132),
        .\remden_reg[20]_0 (\remden_reg[20] ),
        .\remden_reg[20]_1 (dadd_n_56),
        .\remden_reg[21]_0 (\remden_reg[21] ),
        .\remden_reg[21]_1 (dadd_n_55),
        .\remden_reg[22]_0 (\remden_reg[22] ),
        .\remden_reg[22]_1 (dadd_n_54),
        .\remden_reg[23]_0 (\remden_reg[23] ),
        .\remden_reg[23]_1 (dadd_n_53),
        .\remden_reg[24]_0 (\remden_reg[24] ),
        .\remden_reg[24]_1 (dadd_n_52),
        .\remden_reg[25]_0 (\remden_reg[25] ),
        .\remden_reg[25]_1 (dadd_n_51),
        .\remden_reg[26]_0 (\remden_reg[26] ),
        .\remden_reg[26]_1 (\remden_reg[26]_0 ),
        .\remden_reg[27]_0 (rden_n_99),
        .\remden_reg[27]_1 (\remden_reg[27] ),
        .\remden_reg[28]_0 (rden_n_70),
        .\remden_reg[28]_1 (rden_n_71),
        .\remden_reg[28]_2 (\remden_reg[28] ),
        .\remden_reg[28]_3 (dctl_n_4),
        .\remden_reg[28]_4 (add_out[28:26]),
        .\remden_reg[29]_0 (rden_n_68),
        .\remden_reg[29]_1 (rden_n_69),
        .\remden_reg[29]_2 (dctl_n_127),
        .\remden_reg[2]_0 (rden_n_96),
        .\remden_reg[2]_1 (dctl_n_131),
        .\remden_reg[30]_0 (rden_n_66),
        .\remden_reg[30]_1 (rden_n_67),
        .\remden_reg[30]_2 (dctl_n_128),
        .\remden_reg[31]_0 (dctl_n_126),
        .\remden_reg[32]_0 (dctl_n_125),
        .\remden_reg[33]_0 (dctl_n_124),
        .\remden_reg[34]_0 (dctl_n_123),
        .\remden_reg[35]_0 (dctl_n_122),
        .\remden_reg[36]_0 (dctl_n_121),
        .\remden_reg[37]_0 (dctl_n_120),
        .\remden_reg[38]_0 ({rden_n_10,rden_n_11,rden_n_12,rden_n_13}),
        .\remden_reg[38]_1 ({rden_n_14,rden_n_15,rden_n_16,rden_n_17}),
        .\remden_reg[38]_2 (dctl_n_119),
        .\remden_reg[39]_0 (dctl_n_118),
        .\remden_reg[3]_0 (rden_n_95),
        .\remden_reg[3]_1 (dctl_n_130),
        .\remden_reg[40]_0 (dctl_n_117),
        .\remden_reg[41]_0 (dctl_n_116),
        .\remden_reg[42]_0 ({rden_n_18,rden_n_19,rden_n_20,rden_n_21}),
        .\remden_reg[42]_1 ({rden_n_22,rden_n_23,rden_n_24,rden_n_25}),
        .\remden_reg[42]_2 (dctl_n_115),
        .\remden_reg[43]_0 (dctl_n_114),
        .\remden_reg[44]_0 (dctl_n_113),
        .\remden_reg[45]_0 (dctl_n_112),
        .\remden_reg[46]_0 ({rden_n_26,rden_n_27,rden_n_28,rden_n_29}),
        .\remden_reg[46]_1 ({rden_n_30,rden_n_31,rden_n_32,rden_n_33}),
        .\remden_reg[46]_2 (dctl_n_111),
        .\remden_reg[47]_0 (dctl_n_110),
        .\remden_reg[48]_0 (dctl_n_109),
        .\remden_reg[49]_0 (dctl_n_108),
        .\remden_reg[4]_0 (rden_n_93),
        .\remden_reg[4]_1 (dctl_n_40),
        .\remden_reg[4]_2 (dctl_n_16),
        .\remden_reg[50]_0 ({rden_n_34,rden_n_35,rden_n_36,rden_n_37}),
        .\remden_reg[50]_1 ({rden_n_38,rden_n_39,rden_n_40,rden_n_41}),
        .\remden_reg[50]_2 (dctl_n_107),
        .\remden_reg[51]_0 (dctl_n_106),
        .\remden_reg[52]_0 (dctl_n_105),
        .\remden_reg[53]_0 (dctl_n_104),
        .\remden_reg[54]_0 ({rden_n_42,rden_n_43,rden_n_44,rden_n_45}),
        .\remden_reg[54]_1 ({rden_n_46,rden_n_47,rden_n_48,rden_n_49}),
        .\remden_reg[54]_2 (dctl_n_103),
        .\remden_reg[55]_0 (dctl_n_102),
        .\remden_reg[56]_0 (dctl_n_101),
        .\remden_reg[57]_0 (dctl_n_100),
        .\remden_reg[58]_0 ({rden_n_50,rden_n_51,rden_n_52,rden_n_53}),
        .\remden_reg[58]_1 ({rden_n_54,rden_n_55,rden_n_56,rden_n_57}),
        .\remden_reg[58]_2 (dctl_n_99),
        .\remden_reg[59]_0 (dctl_n_98),
        .\remden_reg[5]_0 (rden_n_92),
        .\remden_reg[5]_1 (dctl_n_15),
        .\remden_reg[60]_0 (dctl_n_97),
        .\remden_reg[61]_0 (dctl_n_96),
        .\remden_reg[62]_0 ({rden_n_58,rden_n_59,rden_n_60,rden_n_61}),
        .\remden_reg[62]_1 ({rden_n_62,rden_n_63,rden_n_64,rden_n_65}),
        .\remden_reg[62]_2 (dctl_n_95),
        .\remden_reg[63]_0 (dctl_n_94),
        .\remden_reg[64]_0 (rden_n_72),
        .\remden_reg[64]_1 (dctl_n_18),
        .\remden_reg[64]_2 (dctl_n_93),
        .\remden_reg[6]_0 (rden_n_91),
        .\remden_reg[6]_1 (dctl_n_14),
        .\remden_reg[7]_0 (rden_n_90),
        .\remden_reg[7]_1 (dctl_n_13),
        .\remden_reg[8]_0 (rden_n_89),
        .\remden_reg[8]_1 (dctl_n_12),
        .\remden_reg[9]_0 (rden_n_88),
        .\remden_reg[9]_1 (dctl_n_11),
        .rst_n(rst_n));
  niho_div_reg_dso rdso
       (.D({dctl_n_166,dctl_n_167,dctl_n_168,dctl_n_169,dctl_n_170,dctl_n_171,dctl_n_172,dctl_n_173,dctl_n_174,dctl_n_175,dctl_n_176,dctl_n_177,dctl_n_178,dctl_n_179,dctl_n_180,dctl_n_181,dctl_n_182,dctl_n_183,dctl_n_184,dctl_n_185,dctl_n_186,dctl_n_187,dctl_n_188,dctl_n_189,dctl_n_190,dctl_n_191,dctl_n_192,dctl_n_193,dctl_n_194,dctl_n_195,dctl_n_196,dctl_n_197}),
        .DI(den2),
        .E(dctl_n_24),
        .Q(dso_0),
        .chg_quo_sgn_reg(div_crdy_reg),
        .clk(clk),
        .dctl_long_f(dctl_long_f),
        .dctl_sign(dctl_sign),
        .\dso_reg[31]_0 (rdso_n_1),
        .p_0_in(p_0_in),
        .\remden_reg[31] (rdso_n_0),
        .rgf_sr_nh(rgf_sr_nh));
  niho_div_reg_quo rquo
       (.D(p_2_in),
        .E(dctl_n_19),
        .Q({quo,Q}),
        .clk(clk),
        .niho_dsp_c(niho_dsp_c),
        .\niho_dsp_c[31] (\niho_dsp_c[31] ),
        .p_0_in(p_0_in),
        .\tr[31]_i_5 (\tr[31]_i_5 ),
        .\tr[31]_i_5_0 (\tr[31]_i_5_0 ),
        .\tr[31]_i_5_1 (rem),
        .\tr[31]_i_5_2 (\tr[31]_i_5_1 ));
  niho_div_reg_rem rrem
       (.D({dctl_n_134,dctl_n_135,dctl_n_136,dctl_n_137,dctl_n_138,dctl_n_139,dctl_n_140,dctl_n_141,dctl_n_142,dctl_n_143,dctl_n_144,dctl_n_145,dctl_n_146,dctl_n_147,dctl_n_148,dctl_n_149,dctl_n_150,dctl_n_151,dctl_n_152,dctl_n_153,dctl_n_154,dctl_n_155,dctl_n_156,dctl_n_157,dctl_n_158,dctl_n_159,dctl_n_160,dctl_n_161,dctl_n_162,dctl_n_163,dctl_n_164,dctl_n_165}),
        .E(dctl_n_25),
        .Q({rem,\rem_reg[30] }),
        .clk(clk),
        .p_0_in(p_0_in));
endmodule

module niho_alu_mul
   (mul_rslt,
    niho_dsp_b,
    mul_rslt_reg_0,
    mulh,
    mul_a,
    \mul_b_reg[32]_0 ,
    \mul_b_reg[30]_0 ,
    \mul_b_reg[29]_0 ,
    \mul_b_reg[28]_0 ,
    \mul_b_reg[27]_0 ,
    \mul_b_reg[26]_0 ,
    \mul_b_reg[25]_0 ,
    \mul_b_reg[24]_0 ,
    \mul_b_reg[23]_0 ,
    \mul_b_reg[22]_0 ,
    \mul_b_reg[21]_0 ,
    \mul_b_reg[20]_0 ,
    \mul_b_reg[19]_0 ,
    \mul_b_reg[18]_0 ,
    \mul_b_reg[17]_0 ,
    \mul_b_reg[16]_0 ,
    \mul_b_reg[15]_0 ,
    \mul_b_reg[14]_0 ,
    \mul_b_reg[13]_0 ,
    \mul_b_reg[12]_0 ,
    \mul_b_reg[11]_0 ,
    \mul_b_reg[10]_0 ,
    \mul_b_reg[9]_0 ,
    \mul_b_reg[8]_0 ,
    \mul_b_reg[7]_0 ,
    \mul_b_reg[6]_0 ,
    \mul_b_reg[5]_0 ,
    \mul_b_reg[3]_0 ,
    \mul_b_reg[2]_0 ,
    \mul_b_reg[1]_0 ,
    \mul_b_reg[0]_0 ,
    p_0_in,
    mul_rslt0,
    clk,
    rgf_sr_nh,
    \niho_dsp_b[4] ,
    \niho_dsp_b[4]_0 ,
    \mulh_reg[0]_0 ,
    mul_b,
    niho_dsp_c,
    D,
    mul_a_i,
    \mul_a_reg[16]_0 ,
    \mul_b_reg[0]_1 ,
    abus_0,
    \mul_b_reg[32]_1 ,
    bbus_0);
  output mul_rslt;
  output [0:0]niho_dsp_b;
  output mul_rslt_reg_0;
  output [15:0]mulh;
  output [32:0]mul_a;
  output [1:0]\mul_b_reg[32]_0 ;
  output \mul_b_reg[30]_0 ;
  output \mul_b_reg[29]_0 ;
  output \mul_b_reg[28]_0 ;
  output \mul_b_reg[27]_0 ;
  output \mul_b_reg[26]_0 ;
  output \mul_b_reg[25]_0 ;
  output \mul_b_reg[24]_0 ;
  output \mul_b_reg[23]_0 ;
  output \mul_b_reg[22]_0 ;
  output \mul_b_reg[21]_0 ;
  output \mul_b_reg[20]_0 ;
  output \mul_b_reg[19]_0 ;
  output \mul_b_reg[18]_0 ;
  output \mul_b_reg[17]_0 ;
  output \mul_b_reg[16]_0 ;
  output \mul_b_reg[15]_0 ;
  output \mul_b_reg[14]_0 ;
  output \mul_b_reg[13]_0 ;
  output \mul_b_reg[12]_0 ;
  output \mul_b_reg[11]_0 ;
  output \mul_b_reg[10]_0 ;
  output \mul_b_reg[9]_0 ;
  output \mul_b_reg[8]_0 ;
  output \mul_b_reg[7]_0 ;
  output \mul_b_reg[6]_0 ;
  output \mul_b_reg[5]_0 ;
  output \mul_b_reg[3]_0 ;
  output \mul_b_reg[2]_0 ;
  output \mul_b_reg[1]_0 ;
  output \mul_b_reg[0]_0 ;
  input p_0_in;
  input mul_rslt0;
  input clk;
  input rgf_sr_nh;
  input \niho_dsp_b[4] ;
  input \niho_dsp_b[4]_0 ;
  input \mulh_reg[0]_0 ;
  input mul_b;
  input [15:0]niho_dsp_c;
  input [1:0]D;
  input [13:0]mul_a_i;
  input \mul_a_reg[16]_0 ;
  input \mul_b_reg[0]_1 ;
  input [15:0]abus_0;
  input [1:0]\mul_b_reg[32]_1 ;
  input [30:0]bbus_0;

  wire \<const0> ;
  wire \<const1> ;
  wire [1:0]D;
  wire [15:0]abus_0;
  wire [30:0]bbus_0;
  wire clk;
  wire [32:0]mul_a;
  wire [13:0]mul_a_i;
  wire \mul_a_reg[16]_0 ;
  wire mul_b;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[0]_1 ;
  wire \mul_b_reg[10]_0 ;
  wire \mul_b_reg[11]_0 ;
  wire \mul_b_reg[12]_0 ;
  wire \mul_b_reg[13]_0 ;
  wire \mul_b_reg[14]_0 ;
  wire \mul_b_reg[15]_0 ;
  wire \mul_b_reg[16]_0 ;
  wire \mul_b_reg[17]_0 ;
  wire \mul_b_reg[18]_0 ;
  wire \mul_b_reg[19]_0 ;
  wire \mul_b_reg[1]_0 ;
  wire \mul_b_reg[20]_0 ;
  wire \mul_b_reg[21]_0 ;
  wire \mul_b_reg[22]_0 ;
  wire \mul_b_reg[23]_0 ;
  wire \mul_b_reg[24]_0 ;
  wire \mul_b_reg[25]_0 ;
  wire \mul_b_reg[26]_0 ;
  wire \mul_b_reg[27]_0 ;
  wire \mul_b_reg[28]_0 ;
  wire \mul_b_reg[29]_0 ;
  wire \mul_b_reg[2]_0 ;
  wire \mul_b_reg[30]_0 ;
  wire [1:0]\mul_b_reg[32]_0 ;
  wire [1:0]\mul_b_reg[32]_1 ;
  wire \mul_b_reg[3]_0 ;
  wire \mul_b_reg[5]_0 ;
  wire \mul_b_reg[6]_0 ;
  wire \mul_b_reg[7]_0 ;
  wire \mul_b_reg[8]_0 ;
  wire \mul_b_reg[9]_0 ;
  wire \mul_b_reg_n_0_[4] ;
  wire mul_rslt;
  wire mul_rslt0;
  wire mul_rslt_reg_0;
  wire [15:0]mulh;
  wire \mulh_reg[0]_0 ;
  wire [0:0]niho_dsp_b;
  wire \niho_dsp_b[4] ;
  wire \niho_dsp_b[4]_0 ;
  wire [15:0]niho_dsp_c;
  wire p_0_in;
  wire rgf_sr_nh;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  FDRE \mul_a_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[0]),
        .Q(mul_a[0]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[10]),
        .Q(mul_a[10]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[11]),
        .Q(mul_a[11]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[12]),
        .Q(mul_a[12]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[13]),
        .Q(mul_a[13]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[14]),
        .Q(mul_a[14]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[15]),
        .Q(mul_a[15]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[16] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_a_reg[16]_0 ),
        .Q(mul_a[16]),
        .R(p_0_in));
  FDRE \mul_a_reg[17] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[0]),
        .Q(mul_a[17]),
        .R(p_0_in));
  FDRE \mul_a_reg[18] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[1]),
        .Q(mul_a[18]),
        .R(p_0_in));
  FDRE \mul_a_reg[19] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[2]),
        .Q(mul_a[19]),
        .R(p_0_in));
  FDRE \mul_a_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[1]),
        .Q(mul_a[1]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[20] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[3]),
        .Q(mul_a[20]),
        .R(p_0_in));
  FDRE \mul_a_reg[21] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[4]),
        .Q(mul_a[21]),
        .R(p_0_in));
  FDRE \mul_a_reg[22] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[5]),
        .Q(mul_a[22]),
        .R(p_0_in));
  FDRE \mul_a_reg[23] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[6]),
        .Q(mul_a[23]),
        .R(p_0_in));
  FDRE \mul_a_reg[24] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[7]),
        .Q(mul_a[24]),
        .R(p_0_in));
  FDRE \mul_a_reg[25] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[8]),
        .Q(mul_a[25]),
        .R(p_0_in));
  FDRE \mul_a_reg[26] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[9]),
        .Q(mul_a[26]),
        .R(p_0_in));
  FDRE \mul_a_reg[27] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[10]),
        .Q(mul_a[27]),
        .R(p_0_in));
  FDRE \mul_a_reg[28] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[11]),
        .Q(mul_a[28]),
        .R(p_0_in));
  FDRE \mul_a_reg[29] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[12]),
        .Q(mul_a[29]),
        .R(p_0_in));
  FDRE \mul_a_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[2]),
        .Q(mul_a[2]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[30] 
       (.C(clk),
        .CE(mul_b),
        .D(mul_a_i[13]),
        .Q(mul_a[30]),
        .R(p_0_in));
  FDRE \mul_a_reg[31] 
       (.C(clk),
        .CE(mul_b),
        .D(D[0]),
        .Q(mul_a[31]),
        .R(\<const0> ));
  FDRE \mul_a_reg[32] 
       (.C(clk),
        .CE(mul_b),
        .D(D[1]),
        .Q(mul_a[32]),
        .R(\<const0> ));
  FDRE \mul_a_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[3]),
        .Q(mul_a[3]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[4]),
        .Q(mul_a[4]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[5]),
        .Q(mul_a[5]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[6]),
        .Q(mul_a[6]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[7]),
        .Q(mul_a[7]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[8]),
        .Q(mul_a[8]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_a_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(abus_0[9]),
        .Q(mul_a[9]),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[0]),
        .Q(\mul_b_reg[0]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[10]),
        .Q(\mul_b_reg[10]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[11]),
        .Q(\mul_b_reg[11]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[12]),
        .Q(\mul_b_reg[12]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[13]),
        .Q(\mul_b_reg[13]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[14]),
        .Q(\mul_b_reg[14]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[15]),
        .Q(\mul_b_reg[15]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[16] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[16]),
        .Q(\mul_b_reg[16]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[17] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[17]),
        .Q(\mul_b_reg[17]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[18] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[18]),
        .Q(\mul_b_reg[18]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[19] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[19]),
        .Q(\mul_b_reg[19]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[1]),
        .Q(\mul_b_reg[1]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[20] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[20]),
        .Q(\mul_b_reg[20]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[21] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[21]),
        .Q(\mul_b_reg[21]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[22] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[22]),
        .Q(\mul_b_reg[22]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[23] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[23]),
        .Q(\mul_b_reg[23]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[24] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[24]),
        .Q(\mul_b_reg[24]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[25] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[25]),
        .Q(\mul_b_reg[25]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[26] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[26]),
        .Q(\mul_b_reg[26]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[27] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[27]),
        .Q(\mul_b_reg[27]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[28] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[28]),
        .Q(\mul_b_reg[28]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[29] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[29]),
        .Q(\mul_b_reg[29]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[2]),
        .Q(\mul_b_reg[2]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[30] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[30]),
        .Q(\mul_b_reg[30]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[31] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_b_reg[32]_1 [0]),
        .Q(\mul_b_reg[32]_0 [0]),
        .R(\<const0> ));
  FDRE \mul_b_reg[32] 
       (.C(clk),
        .CE(mul_b),
        .D(\mul_b_reg[32]_1 [1]),
        .Q(\mul_b_reg[32]_0 [1]),
        .R(\<const0> ));
  FDRE \mul_b_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[3]),
        .Q(\mul_b_reg[3]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[4]),
        .Q(\mul_b_reg_n_0_[4] ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[5]),
        .Q(\mul_b_reg[5]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[6]),
        .Q(\mul_b_reg[6]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[7]),
        .Q(\mul_b_reg[7]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[8]),
        .Q(\mul_b_reg[8]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE \mul_b_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(bbus_0[9]),
        .Q(\mul_b_reg[9]_0 ),
        .R(\mul_b_reg[0]_1 ));
  FDRE mul_rslt_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(mul_rslt0),
        .Q(mul_rslt),
        .R(p_0_in));
  FDRE \mulh_reg[0] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[0]),
        .Q(mulh[0]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[10] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[10]),
        .Q(mulh[10]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[11] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[11]),
        .Q(mulh[11]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[12] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[12]),
        .Q(mulh[12]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[13] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[13]),
        .Q(mulh[13]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[14] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[14]),
        .Q(mulh[14]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[15] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[15]),
        .Q(mulh[15]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[1] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[1]),
        .Q(mulh[1]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[2] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[2]),
        .Q(mulh[2]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[3] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[3]),
        .Q(mulh[3]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[4] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[4]),
        .Q(mulh[4]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[5] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[5]),
        .Q(mulh[5]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[6] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[6]),
        .Q(mulh[6]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[7] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[7]),
        .Q(mulh[7]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[8] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[8]),
        .Q(mulh[8]),
        .R(\mulh_reg[0]_0 ));
  FDRE \mulh_reg[9] 
       (.C(clk),
        .CE(mul_b),
        .D(niho_dsp_c[9]),
        .Q(mulh[9]),
        .R(\mulh_reg[0]_0 ));
  LUT5 #(
    .INIT(32'h80FF8080)) 
    \niho_dsp_b[4]_INST_0 
       (.I0(rgf_sr_nh),
        .I1(mul_rslt),
        .I2(\mul_b_reg_n_0_[4] ),
        .I3(\niho_dsp_b[4] ),
        .I4(\niho_dsp_b[4]_0 ),
        .O(niho_dsp_b));
  LUT3 #(
    .INIT(8'h4F)) 
    \tr[30]_i_4 
       (.I0(mul_rslt),
        .I1(\niho_dsp_b[4] ),
        .I2(rgf_sr_nh),
        .O(mul_rslt_reg_0));
endmodule

module niho_div_add
   (\rem_reg[30] ,
    D,
    rst_n_0,
    rst_n_1,
    rst_n_2,
    rst_n_3,
    rst_n_4,
    rst_n_5,
    rst_n_6,
    rst_n_7,
    rst_n_8,
    DI,
    S,
    \quo_reg[7] ,
    \quo_reg[7]_0 ,
    \quo_reg[11] ,
    \quo_reg[11]_0 ,
    \quo_reg[15] ,
    \quo_reg[15]_0 ,
    \quo_reg[19] ,
    \quo_reg[19]_0 ,
    \remden_reg[23] ,
    \remden_reg[23]_0 ,
    \quo_reg[27] ,
    \quo_reg[27]_0 ,
    \remden_reg[31] ,
    \remden_reg[31]_0 ,
    \quo_reg[27]_1 ,
    Q,
    O,
    \quo_reg[2] ,
    \quo_reg[1] ,
    \quo_reg[0] ,
    rst_n,
    \remden_reg[25] ,
    \remden_reg[25]_0 ,
    \remden_reg[24] ,
    \remden_reg[23]_1 ,
    \remden_reg[22] ,
    \remden_reg[21] ,
    \remden_reg[20] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] );
  output [22:0]\rem_reg[30] ;
  output [27:0]D;
  output rst_n_0;
  output rst_n_1;
  output rst_n_2;
  output rst_n_3;
  output rst_n_4;
  output rst_n_5;
  output rst_n_6;
  output rst_n_7;
  output rst_n_8;
  input [3:0]DI;
  input [3:0]S;
  input [3:0]\quo_reg[7] ;
  input [3:0]\quo_reg[7]_0 ;
  input [3:0]\quo_reg[11] ;
  input [3:0]\quo_reg[11]_0 ;
  input [3:0]\quo_reg[15] ;
  input [3:0]\quo_reg[15]_0 ;
  input [3:0]\quo_reg[19] ;
  input [3:0]\quo_reg[19]_0 ;
  input [3:0]\remden_reg[23] ;
  input [3:0]\remden_reg[23]_0 ;
  input [3:0]\quo_reg[27] ;
  input [3:0]\quo_reg[27]_0 ;
  input [2:0]\remden_reg[31] ;
  input [3:0]\remden_reg[31]_0 ;
  input \quo_reg[27]_1 ;
  input [23:0]Q;
  input [0:0]O;
  input [0:0]\quo_reg[2] ;
  input [0:0]\quo_reg[1] ;
  input [0:0]\quo_reg[0] ;
  input rst_n;
  input \remden_reg[25] ;
  input \remden_reg[25]_0 ;
  input \remden_reg[24] ;
  input \remden_reg[23]_1 ;
  input \remden_reg[22] ;
  input \remden_reg[21] ;
  input \remden_reg[20] ;
  input \remden_reg[18] ;
  input \remden_reg[17] ;
  input \remden_reg[16] ;

  wire \<const0> ;
  wire [27:0]D;
  wire [3:0]DI;
  wire [0:0]O;
  wire [23:0]Q;
  wire [3:0]S;
  wire [25:16]add_out;
  wire add_out0_carry__0_n_0;
  wire add_out0_carry__0_n_1;
  wire add_out0_carry__0_n_2;
  wire add_out0_carry__0_n_3;
  wire add_out0_carry__1_n_0;
  wire add_out0_carry__1_n_1;
  wire add_out0_carry__1_n_2;
  wire add_out0_carry__1_n_3;
  wire add_out0_carry__2_n_0;
  wire add_out0_carry__2_n_1;
  wire add_out0_carry__2_n_2;
  wire add_out0_carry__2_n_3;
  wire add_out0_carry__3_n_0;
  wire add_out0_carry__3_n_1;
  wire add_out0_carry__3_n_2;
  wire add_out0_carry__3_n_3;
  wire add_out0_carry__4_n_0;
  wire add_out0_carry__4_n_1;
  wire add_out0_carry__4_n_2;
  wire add_out0_carry__4_n_3;
  wire add_out0_carry__5_n_0;
  wire add_out0_carry__5_n_1;
  wire add_out0_carry__5_n_2;
  wire add_out0_carry__5_n_3;
  wire add_out0_carry__6_n_1;
  wire add_out0_carry__6_n_2;
  wire add_out0_carry__6_n_3;
  wire add_out0_carry_n_0;
  wire add_out0_carry_n_1;
  wire add_out0_carry_n_2;
  wire add_out0_carry_n_3;
  wire [0:0]\quo_reg[0] ;
  wire [3:0]\quo_reg[11] ;
  wire [3:0]\quo_reg[11]_0 ;
  wire [3:0]\quo_reg[15] ;
  wire [3:0]\quo_reg[15]_0 ;
  wire [3:0]\quo_reg[19] ;
  wire [3:0]\quo_reg[19]_0 ;
  wire [0:0]\quo_reg[1] ;
  wire [3:0]\quo_reg[27] ;
  wire [3:0]\quo_reg[27]_0 ;
  wire \quo_reg[27]_1 ;
  wire [0:0]\quo_reg[2] ;
  wire [3:0]\quo_reg[7] ;
  wire [3:0]\quo_reg[7]_0 ;
  wire [22:0]\rem_reg[30] ;
  wire \remden_reg[16] ;
  wire \remden_reg[17] ;
  wire \remden_reg[18] ;
  wire \remden_reg[20] ;
  wire \remden_reg[21] ;
  wire \remden_reg[22] ;
  wire [3:0]\remden_reg[23] ;
  wire [3:0]\remden_reg[23]_0 ;
  wire \remden_reg[23]_1 ;
  wire \remden_reg[24] ;
  wire \remden_reg[25] ;
  wire \remden_reg[25]_0 ;
  wire [2:0]\remden_reg[31] ;
  wire [3:0]\remden_reg[31]_0 ;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_1;
  wire rst_n_2;
  wire rst_n_3;
  wire rst_n_4;
  wire rst_n_5;
  wire rst_n_6;
  wire rst_n_7;
  wire rst_n_8;

  GND GND
       (.G(\<const0> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry
       (.CI(\<const0> ),
        .CO({add_out0_carry_n_0,add_out0_carry_n_1,add_out0_carry_n_2,add_out0_carry_n_3}),
        .CYINIT(\<const0> ),
        .DI(DI),
        .O(\rem_reg[30] [3:0]),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__0
       (.CI(add_out0_carry_n_0),
        .CO({add_out0_carry__0_n_0,add_out0_carry__0_n_1,add_out0_carry__0_n_2,add_out0_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[7] ),
        .O(\rem_reg[30] [7:4]),
        .S(\quo_reg[7]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__1
       (.CI(add_out0_carry__0_n_0),
        .CO({add_out0_carry__1_n_0,add_out0_carry__1_n_1,add_out0_carry__1_n_2,add_out0_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[11] ),
        .O(\rem_reg[30] [11:8]),
        .S(\quo_reg[11]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__2
       (.CI(add_out0_carry__1_n_0),
        .CO({add_out0_carry__2_n_0,add_out0_carry__2_n_1,add_out0_carry__2_n_2,add_out0_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[15] ),
        .O(\rem_reg[30] [15:12]),
        .S(\quo_reg[15]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__3
       (.CI(add_out0_carry__2_n_0),
        .CO({add_out0_carry__3_n_0,add_out0_carry__3_n_1,add_out0_carry__3_n_2,add_out0_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[19] ),
        .O({\rem_reg[30] [16],add_out[18:16]}),
        .S(\quo_reg[19]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__4
       (.CI(add_out0_carry__3_n_0),
        .CO({add_out0_carry__4_n_0,add_out0_carry__4_n_1,add_out0_carry__4_n_2,add_out0_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(\remden_reg[23] ),
        .O(add_out[23:20]),
        .S(\remden_reg[23]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__5
       (.CI(add_out0_carry__4_n_0),
        .CO({add_out0_carry__5_n_0,add_out0_carry__5_n_1,add_out0_carry__5_n_2,add_out0_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(\quo_reg[27] ),
        .O({\rem_reg[30] [18:17],add_out[25:24]}),
        .S(\quo_reg[27]_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 add_out0_carry__6
       (.CI(add_out0_carry__5_n_0),
        .CO({add_out0_carry__6_n_1,add_out0_carry__6_n_2,add_out0_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\remden_reg[31] }),
        .O(\rem_reg[30] [22:19]),
        .S(\remden_reg[31]_0 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[0]_i_1 
       (.I0(\rem_reg[30] [0]),
        .I1(\quo_reg[27]_1 ),
        .I2(\quo_reg[0] ),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[10]_i_1 
       (.I0(\rem_reg[30] [10]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[6]),
        .O(D[10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[11]_i_1 
       (.I0(\rem_reg[30] [11]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[7]),
        .O(D[11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[12]_i_1 
       (.I0(\rem_reg[30] [12]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[8]),
        .O(D[12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[13]_i_1 
       (.I0(\rem_reg[30] [13]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[9]),
        .O(D[13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[14]_i_1 
       (.I0(\rem_reg[30] [14]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[10]),
        .O(D[14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[15]_i_1 
       (.I0(\rem_reg[30] [15]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[11]),
        .O(D[15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[16]_i_1 
       (.I0(add_out[16]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[12]),
        .O(D[16]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[17]_i_1 
       (.I0(add_out[17]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[13]),
        .O(D[17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[18]_i_1 
       (.I0(add_out[18]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[14]),
        .O(D[18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[19]_i_1 
       (.I0(\rem_reg[30] [16]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[15]),
        .O(D[19]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[1]_i_1 
       (.I0(\rem_reg[30] [1]),
        .I1(\quo_reg[27]_1 ),
        .I2(\quo_reg[1] ),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[20]_i_1 
       (.I0(add_out[20]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[16]),
        .O(D[20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[21]_i_1 
       (.I0(add_out[21]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[17]),
        .O(D[21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[22]_i_1 
       (.I0(add_out[22]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[18]),
        .O(D[22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[23]_i_1 
       (.I0(add_out[23]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[19]),
        .O(D[23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[24]_i_1 
       (.I0(add_out[24]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[20]),
        .O(D[24]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[25]_i_1 
       (.I0(add_out[25]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[21]),
        .O(D[25]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[26]_i_1 
       (.I0(\rem_reg[30] [17]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[22]),
        .O(D[26]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[27]_i_1 
       (.I0(\rem_reg[30] [18]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[23]),
        .O(D[27]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[2]_i_1 
       (.I0(\rem_reg[30] [2]),
        .I1(\quo_reg[27]_1 ),
        .I2(\quo_reg[2] ),
        .O(D[2]));
  LUT3 #(
    .INIT(8'h8B)) 
    \quo[3]_i_1 
       (.I0(\rem_reg[30] [3]),
        .I1(\quo_reg[27]_1 ),
        .I2(O),
        .O(D[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[4]_i_1 
       (.I0(\rem_reg[30] [4]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[0]),
        .O(D[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[5]_i_1 
       (.I0(\rem_reg[30] [5]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[1]),
        .O(D[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[6]_i_1 
       (.I0(\rem_reg[30] [6]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[2]),
        .O(D[6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[7]_i_1 
       (.I0(\rem_reg[30] [7]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[3]),
        .O(D[7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[8]_i_1 
       (.I0(\rem_reg[30] [8]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[4]),
        .O(D[8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[9]_i_1 
       (.I0(\rem_reg[30] [9]),
        .I1(\quo_reg[27]_1 ),
        .I2(Q[5]),
        .O(D[9]));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[16]_i_1 
       (.I0(rst_n),
        .I1(add_out[16]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[16] ),
        .O(rst_n_8));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[17]_i_1 
       (.I0(rst_n),
        .I1(add_out[17]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[17] ),
        .O(rst_n_7));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[18]_i_1 
       (.I0(rst_n),
        .I1(add_out[18]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[18] ),
        .O(rst_n_6));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[20]_i_1 
       (.I0(rst_n),
        .I1(add_out[20]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[20] ),
        .O(rst_n_5));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[21]_i_1 
       (.I0(rst_n),
        .I1(add_out[21]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[21] ),
        .O(rst_n_4));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[22]_i_1 
       (.I0(rst_n),
        .I1(add_out[22]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[22] ),
        .O(rst_n_3));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[23]_i_1 
       (.I0(rst_n),
        .I1(add_out[23]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[23]_1 ),
        .O(rst_n_2));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[24]_i_1 
       (.I0(rst_n),
        .I1(add_out[24]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[24] ),
        .O(rst_n_1));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[25]_i_1 
       (.I0(rst_n),
        .I1(add_out[25]),
        .I2(\remden_reg[25] ),
        .I3(\remden_reg[25]_0 ),
        .O(rst_n_0));
endmodule

module niho_div_ctl
   (dctl_long_f,
    dctl_sign_f,
    div_crdy_reg_0,
    \sr_reg[8] ,
    \dctl_stat_reg[3] ,
    div_crdy_reg_1,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \dctl_stat_reg[2] ,
    \dctl_stat_reg[1] ,
    E,
    D,
    div_crdy_reg_2,
    \dctl_stat_reg[2]_0 ,
    \rem_reg[3] ,
    \dso_reg[31] ,
    S,
    div_crdy_reg_3,
    crdy_0,
    rst_n_0,
    div_crdy_reg_4,
    \rem_reg[30] ,
    \rem_reg[27] ,
    \rem_reg[23] ,
    \rem_reg[19] ,
    \rem_reg[15] ,
    \rem_reg[11] ,
    \rem_reg[7] ,
    \rem_reg[27]_0 ,
    \rem_reg[23]_0 ,
    \rem_reg[19]_0 ,
    \rem_reg[15]_0 ,
    \rem_reg[11]_0 ,
    \rem_reg[7]_0 ,
    rst_n_1,
    rst_n_2,
    rst_n_3,
    rst_n_4,
    rst_n_5,
    rst_n_6,
    rst_n_7,
    rst_n_8,
    rst_n_9,
    rst_n_10,
    rst_n_11,
    rst_n_12,
    rst_n_13,
    rst_n_14,
    rst_n_15,
    rst_n_16,
    rst_n_17,
    rst_n_18,
    rst_n_19,
    rst_n_20,
    rst_n_21,
    rst_n_22,
    rst_n_23,
    rst_n_24,
    rst_n_25,
    rst_n_26,
    rst_n_27,
    rst_n_28,
    rst_n_29,
    \remden_reg[28] ,
    \remden_reg[28]_0 ,
    \remden_reg[28]_1 ,
    \remden_reg[28]_2 ,
    rst_n_30,
    rst_n_31,
    rst_n_32,
    rst_n_33,
    rst_n_34,
    rst_n_35,
    rst_n_36,
    rst_n_37,
    \rem_reg[31] ,
    \sr_reg[8]_11 ,
    p_0_in,
    fdiv_rem_msb_f_reg,
    clk,
    dctl_sign,
    \remden_reg[31] ,
    abus_0,
    rgf_sr_nh,
    \remden_reg[15] ,
    \remden_reg[14] ,
    \remden_reg[13] ,
    \remden_reg[12] ,
    \remden_reg[11] ,
    \remden_reg[10] ,
    \remden_reg[9] ,
    \remden_reg[8] ,
    \remden_reg[7] ,
    \remden_reg[6] ,
    \remden_reg[5] ,
    \remden_reg[4] ,
    Q,
    add_out0_carry__6,
    add_out0_carry__2_i_11,
    add_out0_carry__2_i_9,
    add_out0_carry__4_i_10,
    add_out0_carry__4_i_9,
    add_out0_carry__5_i_12,
    add_out0_carry__5_i_10,
    DI,
    add_out0_carry__6_i_9,
    add_out0_carry__6_i_10,
    add_out0_carry__5_i_11,
    add_out0_carry__4_i_11,
    add_out0_carry__4_i_12,
    add_out0_carry__3_i_9,
    add_out0_carry__3_i_10,
    add_out0_carry__3_i_11,
    add_out0_carry__3_i_12,
    add_out0_carry__2_i_12,
    \rem_reg[31]_0 ,
    add_out0_carry__2_i_10,
    \remden_reg[31]_0 ,
    den2,
    \dctl_stat_reg[3]_0 ,
    chg_quo_sgn_reg,
    \dctl_stat_reg[2]_1 ,
    chg_rem_sgn0,
    crdy,
    \bcmd[2]_INST_0_i_1 ,
    rst_n,
    out,
    \niho_dsp_a[32]_INST_0_i_12 ,
    fdiv_rem,
    \dso_reg[19] ,
    \dso_reg[19]_0 ,
    \dso_reg[19]_1 ,
    \dso_reg[19]_2 ,
    \dso_reg[23] ,
    \dso_reg[23]_0 ,
    \dso_reg[23]_1 ,
    \dso_reg[23]_2 ,
    \dso_reg[27] ,
    \dso_reg[27]_0 ,
    \dso_reg[27]_1 ,
    \dso_reg[27]_2 ,
    \dso_reg[31]_0 ,
    \dso_reg[31]_1 ,
    \dso_reg[31]_2 ,
    \dso_reg[31]_3 ,
    \remden_reg[31]_1 ,
    \remden_reg[29] ,
    \remden_reg[30] ,
    \remden_reg[19] ,
    bbus_0);
  output dctl_long_f;
  output dctl_sign_f;
  output div_crdy_reg_0;
  output \sr_reg[8] ;
  output \dctl_stat_reg[3] ;
  output div_crdy_reg_1;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \dctl_stat_reg[2] ;
  output \dctl_stat_reg[1] ;
  output [0:0]E;
  output [3:0]D;
  output [0:0]div_crdy_reg_2;
  output [0:0]\dctl_stat_reg[2]_0 ;
  output [3:0]\rem_reg[3] ;
  output [3:0]\dso_reg[31] ;
  output [3:0]S;
  output div_crdy_reg_3;
  output crdy_0;
  output rst_n_0;
  output div_crdy_reg_4;
  output [2:0]\rem_reg[30] ;
  output [3:0]\rem_reg[27] ;
  output [3:0]\rem_reg[23] ;
  output [3:0]\rem_reg[19] ;
  output [3:0]\rem_reg[15] ;
  output [3:0]\rem_reg[11] ;
  output [3:0]\rem_reg[7] ;
  output [3:0]\rem_reg[27]_0 ;
  output [3:0]\rem_reg[23]_0 ;
  output [3:0]\rem_reg[19]_0 ;
  output [3:0]\rem_reg[15]_0 ;
  output [3:0]\rem_reg[11]_0 ;
  output [3:0]\rem_reg[7]_0 ;
  output rst_n_1;
  output rst_n_2;
  output rst_n_3;
  output rst_n_4;
  output rst_n_5;
  output rst_n_6;
  output rst_n_7;
  output rst_n_8;
  output rst_n_9;
  output rst_n_10;
  output rst_n_11;
  output rst_n_12;
  output rst_n_13;
  output rst_n_14;
  output rst_n_15;
  output rst_n_16;
  output rst_n_17;
  output rst_n_18;
  output rst_n_19;
  output rst_n_20;
  output rst_n_21;
  output rst_n_22;
  output rst_n_23;
  output rst_n_24;
  output rst_n_25;
  output rst_n_26;
  output rst_n_27;
  output rst_n_28;
  output rst_n_29;
  output \remden_reg[28] ;
  output \remden_reg[28]_0 ;
  output \remden_reg[28]_1 ;
  output \remden_reg[28]_2 ;
  output rst_n_30;
  output rst_n_31;
  output rst_n_32;
  output rst_n_33;
  output rst_n_34;
  output rst_n_35;
  output rst_n_36;
  output rst_n_37;
  output [31:0]\rem_reg[31] ;
  output [31:0]\sr_reg[8]_11 ;
  input p_0_in;
  input [0:0]fdiv_rem_msb_f_reg;
  input clk;
  input dctl_sign;
  input [20:0]\remden_reg[31] ;
  input [15:0]abus_0;
  input rgf_sr_nh;
  input \remden_reg[15] ;
  input \remden_reg[14] ;
  input \remden_reg[13] ;
  input \remden_reg[12] ;
  input \remden_reg[11] ;
  input \remden_reg[10] ;
  input \remden_reg[9] ;
  input \remden_reg[8] ;
  input \remden_reg[7] ;
  input \remden_reg[6] ;
  input \remden_reg[5] ;
  input \remden_reg[4] ;
  input [31:0]Q;
  input [31:0]add_out0_carry__6;
  input add_out0_carry__2_i_11;
  input add_out0_carry__2_i_9;
  input add_out0_carry__4_i_10;
  input add_out0_carry__4_i_9;
  input add_out0_carry__5_i_12;
  input add_out0_carry__5_i_10;
  input [0:0]DI;
  input [0:0]add_out0_carry__6_i_9;
  input add_out0_carry__6_i_10;
  input add_out0_carry__5_i_11;
  input add_out0_carry__4_i_11;
  input add_out0_carry__4_i_12;
  input add_out0_carry__3_i_9;
  input add_out0_carry__3_i_10;
  input add_out0_carry__3_i_11;
  input add_out0_carry__3_i_12;
  input add_out0_carry__2_i_12;
  input [31:0]\rem_reg[31]_0 ;
  input add_out0_carry__2_i_10;
  input \remden_reg[31]_0 ;
  input [0:0]den2;
  input \dctl_stat_reg[3]_0 ;
  input chg_quo_sgn_reg;
  input \dctl_stat_reg[2]_1 ;
  input chg_rem_sgn0;
  input crdy;
  input \bcmd[2]_INST_0_i_1 ;
  input rst_n;
  input [0:0]out;
  input [0:0]\niho_dsp_a[32]_INST_0_i_12 ;
  input [31:0]fdiv_rem;
  input \dso_reg[19] ;
  input \dso_reg[19]_0 ;
  input \dso_reg[19]_1 ;
  input \dso_reg[19]_2 ;
  input \dso_reg[23] ;
  input \dso_reg[23]_0 ;
  input \dso_reg[23]_1 ;
  input \dso_reg[23]_2 ;
  input \dso_reg[27] ;
  input \dso_reg[27]_0 ;
  input \dso_reg[27]_1 ;
  input \dso_reg[27]_2 ;
  input \dso_reg[31]_0 ;
  input \dso_reg[31]_1 ;
  input \dso_reg[31]_2 ;
  input \dso_reg[31]_3 ;
  input \remden_reg[31]_1 ;
  input \remden_reg[29] ;
  input \remden_reg[30] ;
  input \remden_reg[19] ;
  input [15:0]bbus_0;

  wire \<const1> ;
  wire [3:0]D;
  wire [0:0]DI;
  wire [0:0]E;
  wire [31:0]Q;
  wire [3:0]S;
  wire [15:0]abus_0;
  wire add_out0_carry__2_i_10;
  wire add_out0_carry__2_i_11;
  wire add_out0_carry__2_i_12;
  wire add_out0_carry__2_i_9;
  wire add_out0_carry__3_i_10;
  wire add_out0_carry__3_i_11;
  wire add_out0_carry__3_i_12;
  wire add_out0_carry__3_i_9;
  wire add_out0_carry__4_i_10;
  wire add_out0_carry__4_i_11;
  wire add_out0_carry__4_i_12;
  wire add_out0_carry__4_i_9;
  wire add_out0_carry__5_i_10;
  wire add_out0_carry__5_i_11;
  wire add_out0_carry__5_i_12;
  wire [31:0]add_out0_carry__6;
  wire add_out0_carry__6_i_10;
  wire [0:0]add_out0_carry__6_i_9;
  wire [15:0]bbus_0;
  wire \bcmd[2]_INST_0_i_1 ;
  wire chg_quo_sgn_reg;
  wire chg_rem_sgn0;
  wire clk;
  wire crdy;
  wire crdy_0;
  wire dctl_long;
  wire dctl_long_f;
  wire dctl_sign;
  wire dctl_sign_f;
  wire \dctl_stat_reg[1] ;
  wire \dctl_stat_reg[2] ;
  wire [0:0]\dctl_stat_reg[2]_0 ;
  wire \dctl_stat_reg[2]_1 ;
  wire \dctl_stat_reg[3] ;
  wire \dctl_stat_reg[3]_0 ;
  wire [0:0]den2;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  wire [0:0]div_crdy_reg_2;
  wire div_crdy_reg_3;
  wire div_crdy_reg_4;
  wire \dso_reg[19] ;
  wire \dso_reg[19]_0 ;
  wire \dso_reg[19]_1 ;
  wire \dso_reg[19]_2 ;
  wire \dso_reg[23] ;
  wire \dso_reg[23]_0 ;
  wire \dso_reg[23]_1 ;
  wire \dso_reg[23]_2 ;
  wire \dso_reg[27] ;
  wire \dso_reg[27]_0 ;
  wire \dso_reg[27]_1 ;
  wire \dso_reg[27]_2 ;
  wire [3:0]\dso_reg[31] ;
  wire \dso_reg[31]_0 ;
  wire \dso_reg[31]_1 ;
  wire \dso_reg[31]_2 ;
  wire \dso_reg[31]_3 ;
  wire [31:0]fdiv_rem;
  wire [0:0]fdiv_rem_msb_f_reg;
  wire fsm_n_35;
  wire [0:0]\niho_dsp_a[32]_INST_0_i_12 ;
  wire [0:0]out;
  wire p_0_in;
  wire [3:0]\rem_reg[11] ;
  wire [3:0]\rem_reg[11]_0 ;
  wire [3:0]\rem_reg[15] ;
  wire [3:0]\rem_reg[15]_0 ;
  wire [3:0]\rem_reg[19] ;
  wire [3:0]\rem_reg[19]_0 ;
  wire [3:0]\rem_reg[23] ;
  wire [3:0]\rem_reg[23]_0 ;
  wire [3:0]\rem_reg[27] ;
  wire [3:0]\rem_reg[27]_0 ;
  wire [2:0]\rem_reg[30] ;
  wire [31:0]\rem_reg[31] ;
  wire [31:0]\rem_reg[31]_0 ;
  wire [3:0]\rem_reg[3] ;
  wire [3:0]\rem_reg[7] ;
  wire [3:0]\rem_reg[7]_0 ;
  wire \remden[64]_i_6_n_0 ;
  wire \remden_reg[10] ;
  wire \remden_reg[11] ;
  wire \remden_reg[12] ;
  wire \remden_reg[13] ;
  wire \remden_reg[14] ;
  wire \remden_reg[15] ;
  wire \remden_reg[19] ;
  wire \remden_reg[28] ;
  wire \remden_reg[28]_0 ;
  wire \remden_reg[28]_1 ;
  wire \remden_reg[28]_2 ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire [20:0]\remden_reg[31] ;
  wire \remden_reg[31]_0 ;
  wire \remden_reg[31]_1 ;
  wire \remden_reg[4] ;
  wire \remden_reg[5] ;
  wire \remden_reg[6] ;
  wire \remden_reg[7] ;
  wire \remden_reg[8] ;
  wire \remden_reg[9] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_1;
  wire rst_n_10;
  wire rst_n_11;
  wire rst_n_12;
  wire rst_n_13;
  wire rst_n_14;
  wire rst_n_15;
  wire rst_n_16;
  wire rst_n_17;
  wire rst_n_18;
  wire rst_n_19;
  wire rst_n_2;
  wire rst_n_20;
  wire rst_n_21;
  wire rst_n_22;
  wire rst_n_23;
  wire rst_n_24;
  wire rst_n_25;
  wire rst_n_26;
  wire rst_n_27;
  wire rst_n_28;
  wire rst_n_29;
  wire rst_n_3;
  wire rst_n_30;
  wire rst_n_31;
  wire rst_n_32;
  wire rst_n_33;
  wire rst_n_34;
  wire rst_n_35;
  wire rst_n_36;
  wire rst_n_37;
  wire rst_n_4;
  wire rst_n_5;
  wire rst_n_6;
  wire rst_n_7;
  wire rst_n_8;
  wire rst_n_9;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire [31:0]\sr_reg[8]_11 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'h07)) 
    \bcmd[2]_INST_0_i_3 
       (.I0(div_crdy_reg_0),
        .I1(crdy),
        .I2(\bcmd[2]_INST_0_i_1 ),
        .O(div_crdy_reg_3));
  LUT4 #(
    .INIT(16'h0080)) 
    \ccmd[0]_INST_0_i_16 
       (.I0(div_crdy_reg_0),
        .I1(crdy),
        .I2(out),
        .I3(\niho_dsp_a[32]_INST_0_i_12 ),
        .O(div_crdy_reg_4));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[3]_INST_0_i_14 
       (.I0(crdy),
        .I1(div_crdy_reg_0),
        .O(crdy_0));
  FDRE dctl_long_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_long),
        .Q(dctl_long_f),
        .R(p_0_in));
  FDRE dctl_sign_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_sign),
        .Q(dctl_sign_f),
        .R(p_0_in));
  FDSE div_crdy_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fsm_n_35),
        .Q(div_crdy_reg_0),
        .S(p_0_in));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_4 
       (.I0(div_crdy_reg_0),
        .I1(\dctl_stat_reg[2]_1 ),
        .O(div_crdy_reg_1));
  niho_div_fsm fsm
       (.D(D),
        .DI(DI),
        .E(E),
        .Q(Q),
        .S(S),
        .abus_0(abus_0),
        .add_out0_carry__2_i_10_0(add_out0_carry__2_i_10),
        .add_out0_carry__2_i_11_0(add_out0_carry__2_i_11),
        .add_out0_carry__2_i_12_0(add_out0_carry__2_i_12),
        .add_out0_carry__2_i_9_0(add_out0_carry__2_i_9),
        .add_out0_carry__3_i_10_0(add_out0_carry__3_i_10),
        .add_out0_carry__3_i_11_0(add_out0_carry__3_i_11),
        .add_out0_carry__3_i_12_0(add_out0_carry__3_i_12),
        .add_out0_carry__3_i_9_0(add_out0_carry__3_i_9),
        .add_out0_carry__4_i_10_0(add_out0_carry__4_i_10),
        .add_out0_carry__4_i_11_0(add_out0_carry__4_i_11),
        .add_out0_carry__4_i_12_0(add_out0_carry__4_i_12),
        .add_out0_carry__4_i_9_0(add_out0_carry__4_i_9),
        .add_out0_carry__5_i_10_0(add_out0_carry__5_i_10),
        .add_out0_carry__5_i_11_0(add_out0_carry__5_i_11),
        .add_out0_carry__5_i_12_0(add_out0_carry__5_i_12),
        .add_out0_carry__6(add_out0_carry__6),
        .add_out0_carry__6_i_10_0(add_out0_carry__6_i_10),
        .add_out0_carry__6_i_9_0(add_out0_carry__6_i_9),
        .bbus_0(bbus_0),
        .chg_quo_sgn_reg_0(chg_quo_sgn_reg),
        .chg_rem_sgn0(chg_rem_sgn0),
        .clk(clk),
        .dctl_long(dctl_long),
        .dctl_long_f_reg(dctl_long_f),
        .dctl_long_f_reg_0(div_crdy_reg_0),
        .dctl_sign(dctl_sign),
        .\dctl_stat_reg[1]_0 (\dctl_stat_reg[1] ),
        .\dctl_stat_reg[2]_0 (\dctl_stat_reg[2] ),
        .\dctl_stat_reg[2]_1 (\dctl_stat_reg[2]_0 ),
        .\dctl_stat_reg[2]_2 (\dctl_stat_reg[2]_1 ),
        .\dctl_stat_reg[3]_0 (\dctl_stat_reg[3] ),
        .\dctl_stat_reg[3]_1 (\dctl_stat_reg[3]_0 ),
        .den2(den2),
        .div_crdy_reg(div_crdy_reg_2),
        .div_crdy_reg_0(fsm_n_35),
        .\dso_reg[19] (\dso_reg[19] ),
        .\dso_reg[19]_0 (\dso_reg[19]_0 ),
        .\dso_reg[19]_1 (\dso_reg[19]_1 ),
        .\dso_reg[19]_2 (\dso_reg[19]_2 ),
        .\dso_reg[23] (\dso_reg[23] ),
        .\dso_reg[23]_0 (\dso_reg[23]_0 ),
        .\dso_reg[23]_1 (\dso_reg[23]_1 ),
        .\dso_reg[23]_2 (\dso_reg[23]_2 ),
        .\dso_reg[27] (\dso_reg[27] ),
        .\dso_reg[27]_0 (\dso_reg[27]_0 ),
        .\dso_reg[27]_1 (\dso_reg[27]_1 ),
        .\dso_reg[27]_2 (\dso_reg[27]_2 ),
        .\dso_reg[31] (\dso_reg[31] ),
        .\dso_reg[31]_0 (\dso_reg[31]_0 ),
        .\dso_reg[31]_1 (\dso_reg[31]_1 ),
        .\dso_reg[31]_2 (\dso_reg[31]_2 ),
        .\dso_reg[31]_3 (\dso_reg[31]_3 ),
        .fdiv_rem(fdiv_rem),
        .fdiv_rem_msb_f_reg_0(fdiv_rem_msb_f_reg),
        .p_0_in(p_0_in),
        .\rem_reg[11] (\rem_reg[11] ),
        .\rem_reg[11]_0 (\rem_reg[11]_0 ),
        .\rem_reg[15] (\rem_reg[15] ),
        .\rem_reg[15]_0 (\rem_reg[15]_0 ),
        .\rem_reg[19] (\rem_reg[19] ),
        .\rem_reg[19]_0 (\rem_reg[19]_0 ),
        .\rem_reg[23] (\rem_reg[23] ),
        .\rem_reg[23]_0 (\rem_reg[23]_0 ),
        .\rem_reg[27] (\rem_reg[27] ),
        .\rem_reg[27]_0 (\rem_reg[27]_0 ),
        .\rem_reg[30] (\rem_reg[30] ),
        .\rem_reg[31] (\rem_reg[31] ),
        .\rem_reg[31]_0 (\rem_reg[31]_0 ),
        .\rem_reg[3] (\rem_reg[3] ),
        .\rem_reg[7] (\rem_reg[7] ),
        .\rem_reg[7]_0 (\rem_reg[7]_0 ),
        .\remden_reg[0] (div_crdy_reg_1),
        .\remden_reg[10] (\remden_reg[10] ),
        .\remden_reg[11] (\remden_reg[11] ),
        .\remden_reg[12] (\remden_reg[12] ),
        .\remden_reg[13] (\remden_reg[13] ),
        .\remden_reg[14] (\remden_reg[14] ),
        .\remden_reg[15] (\remden_reg[15] ),
        .\remden_reg[19] (\remden_reg[19] ),
        .\remden_reg[28] (\remden_reg[28] ),
        .\remden_reg[28]_0 (\remden_reg[28]_0 ),
        .\remden_reg[28]_1 (\remden_reg[28]_1 ),
        .\remden_reg[28]_2 (\remden_reg[28]_2 ),
        .\remden_reg[29] (\remden_reg[29] ),
        .\remden_reg[30] (\remden_reg[30] ),
        .\remden_reg[31] (\remden_reg[31] ),
        .\remden_reg[31]_0 (\remden_reg[31]_0 ),
        .\remden_reg[31]_1 (\remden_reg[31]_1 ),
        .\remden_reg[4] (\remden_reg[4] ),
        .\remden_reg[5] (\remden_reg[5] ),
        .\remden_reg[64] (\remden[64]_i_6_n_0 ),
        .\remden_reg[6] (\remden_reg[6] ),
        .\remden_reg[7] (\remden_reg[7] ),
        .\remden_reg[8] (\remden_reg[8] ),
        .\remden_reg[9] (\remden_reg[9] ),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .rst_n_0(rst_n_0),
        .rst_n_1(rst_n_1),
        .rst_n_10(rst_n_10),
        .rst_n_11(rst_n_11),
        .rst_n_12(rst_n_12),
        .rst_n_13(rst_n_13),
        .rst_n_14(rst_n_14),
        .rst_n_15(rst_n_15),
        .rst_n_16(rst_n_16),
        .rst_n_17(rst_n_17),
        .rst_n_18(rst_n_18),
        .rst_n_19(rst_n_19),
        .rst_n_2(rst_n_2),
        .rst_n_20(rst_n_20),
        .rst_n_21(rst_n_21),
        .rst_n_22(rst_n_22),
        .rst_n_23(rst_n_23),
        .rst_n_24(rst_n_24),
        .rst_n_25(rst_n_25),
        .rst_n_26(rst_n_26),
        .rst_n_27(rst_n_27),
        .rst_n_28(rst_n_28),
        .rst_n_29(rst_n_29),
        .rst_n_3(rst_n_3),
        .rst_n_30(rst_n_30),
        .rst_n_31(rst_n_31),
        .rst_n_32(rst_n_32),
        .rst_n_33(rst_n_33),
        .rst_n_34(rst_n_34),
        .rst_n_35(rst_n_35),
        .rst_n_36(rst_n_36),
        .rst_n_37(rst_n_37),
        .rst_n_4(rst_n_4),
        .rst_n_5(rst_n_5),
        .rst_n_6(rst_n_6),
        .rst_n_7(rst_n_7),
        .rst_n_8(rst_n_8),
        .rst_n_9(rst_n_9),
        .\sr_reg[8] (\sr_reg[8] ),
        .\sr_reg[8]_0 (\sr_reg[8]_0 ),
        .\sr_reg[8]_1 (\sr_reg[8]_1 ),
        .\sr_reg[8]_10 (\sr_reg[8]_10 ),
        .\sr_reg[8]_11 (\sr_reg[8]_11 ),
        .\sr_reg[8]_2 (\sr_reg[8]_2 ),
        .\sr_reg[8]_3 (\sr_reg[8]_3 ),
        .\sr_reg[8]_4 (\sr_reg[8]_4 ),
        .\sr_reg[8]_5 (\sr_reg[8]_5 ),
        .\sr_reg[8]_6 (\sr_reg[8]_6 ),
        .\sr_reg[8]_7 (\sr_reg[8]_7 ),
        .\sr_reg[8]_8 (\sr_reg[8]_8 ),
        .\sr_reg[8]_9 (\sr_reg[8]_9 ));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_6 
       (.I0(div_crdy_reg_1),
        .I1(rst_n),
        .O(\remden[64]_i_6_n_0 ));
endmodule

module niho_div_fdiv
   (O,
    rem2_carry__7_i_1_0,
    rem1_carry__7_i_1_0,
    fdiv_rem,
    rem0_carry__7_i_1_0,
    p_1_in5_in,
    DI,
    S,
    rem2_carry__0_0,
    rem2_carry__0_1,
    rem2_carry__1_0,
    rem2_carry__1_1,
    rem2_carry__2_0,
    rem2_carry__2_1,
    rem2_carry__3_0,
    rem2_carry__3_1,
    rem2_carry__4_0,
    rem2_carry__4_1,
    rem2_carry__5_0,
    rem2_carry__5_1,
    rem2_carry__6_0,
    rem2_carry__6_1,
    \quo_reg[3] ,
    rem1_carry_0,
    rem1_carry_1,
    rem0_carry_0,
    rem0_carry_1,
    \remden_reg[35] ,
    \remden_reg[35]_0 ,
    Q);
  output [0:0]O;
  output [0:0]rem2_carry__7_i_1_0;
  output [0:0]rem1_carry__7_i_1_0;
  output [31:0]fdiv_rem;
  output [0:0]rem0_carry__7_i_1_0;
  input [0:0]p_1_in5_in;
  input [3:0]DI;
  input [3:0]S;
  input [3:0]rem2_carry__0_0;
  input [3:0]rem2_carry__0_1;
  input [3:0]rem2_carry__1_0;
  input [3:0]rem2_carry__1_1;
  input [3:0]rem2_carry__2_0;
  input [3:0]rem2_carry__2_1;
  input [3:0]rem2_carry__3_0;
  input [3:0]rem2_carry__3_1;
  input [3:0]rem2_carry__4_0;
  input [3:0]rem2_carry__4_1;
  input [3:0]rem2_carry__5_0;
  input [3:0]rem2_carry__5_1;
  input [3:0]rem2_carry__6_0;
  input [3:0]rem2_carry__6_1;
  input [0:0]\quo_reg[3] ;
  input [0:0]rem1_carry_0;
  input [0:0]rem1_carry_1;
  input [0:0]rem0_carry_0;
  input [0:0]rem0_carry_1;
  input \remden_reg[35] ;
  input [0:0]\remden_reg[35]_0 ;
  input [30:0]Q;

  wire \<const0> ;
  wire [3:0]DI;
  wire [0:0]O;
  wire [30:0]Q;
  wire [3:0]S;
  wire [31:0]fdiv_rem;
  wire [0:0]p_1_in3_in;
  wire [0:0]p_1_in5_in;
  wire [0:0]\quo_reg[3] ;
  wire [0:0]rem0_carry_0;
  wire [0:0]rem0_carry_1;
  wire rem0_carry__0_i_1_n_0;
  wire rem0_carry__0_i_2_n_0;
  wire rem0_carry__0_i_3_n_0;
  wire rem0_carry__0_i_4_n_0;
  wire rem0_carry__0_n_0;
  wire rem0_carry__0_n_1;
  wire rem0_carry__0_n_2;
  wire rem0_carry__0_n_3;
  wire rem0_carry__1_i_1_n_0;
  wire rem0_carry__1_i_2_n_0;
  wire rem0_carry__1_i_3_n_0;
  wire rem0_carry__1_i_4_n_0;
  wire rem0_carry__1_n_0;
  wire rem0_carry__1_n_1;
  wire rem0_carry__1_n_2;
  wire rem0_carry__1_n_3;
  wire rem0_carry__2_i_1_n_0;
  wire rem0_carry__2_i_2_n_0;
  wire rem0_carry__2_i_3_n_0;
  wire rem0_carry__2_i_4_n_0;
  wire rem0_carry__2_n_0;
  wire rem0_carry__2_n_1;
  wire rem0_carry__2_n_2;
  wire rem0_carry__2_n_3;
  wire rem0_carry__3_i_1_n_0;
  wire rem0_carry__3_i_2_n_0;
  wire rem0_carry__3_i_3_n_0;
  wire rem0_carry__3_i_4_n_0;
  wire rem0_carry__3_n_0;
  wire rem0_carry__3_n_1;
  wire rem0_carry__3_n_2;
  wire rem0_carry__3_n_3;
  wire rem0_carry__4_i_1_n_0;
  wire rem0_carry__4_i_2_n_0;
  wire rem0_carry__4_i_3_n_0;
  wire rem0_carry__4_i_4_n_0;
  wire rem0_carry__4_n_0;
  wire rem0_carry__4_n_1;
  wire rem0_carry__4_n_2;
  wire rem0_carry__4_n_3;
  wire rem0_carry__5_i_1_n_0;
  wire rem0_carry__5_i_2_n_0;
  wire rem0_carry__5_i_3_n_0;
  wire rem0_carry__5_i_4_n_0;
  wire rem0_carry__5_n_0;
  wire rem0_carry__5_n_1;
  wire rem0_carry__5_n_2;
  wire rem0_carry__5_n_3;
  wire rem0_carry__6_i_1_n_0;
  wire rem0_carry__6_i_2_n_0;
  wire rem0_carry__6_i_3_n_0;
  wire rem0_carry__6_i_4_n_0;
  wire rem0_carry__6_n_0;
  wire rem0_carry__6_n_1;
  wire rem0_carry__6_n_2;
  wire rem0_carry__6_n_3;
  wire [0:0]rem0_carry__7_i_1_0;
  wire rem0_carry__7_i_1_n_0;
  wire rem0_carry_i_1_n_0;
  wire rem0_carry_i_2_n_0;
  wire rem0_carry_i_3_n_0;
  wire rem0_carry_i_4_n_0;
  wire rem0_carry_n_0;
  wire rem0_carry_n_1;
  wire rem0_carry_n_2;
  wire rem0_carry_n_3;
  wire [32:1]rem1;
  wire [0:0]rem1_carry_0;
  wire [0:0]rem1_carry_1;
  wire rem1_carry__0_i_1_n_0;
  wire rem1_carry__0_i_2_n_0;
  wire rem1_carry__0_i_3_n_0;
  wire rem1_carry__0_i_4_n_0;
  wire rem1_carry__0_n_0;
  wire rem1_carry__0_n_1;
  wire rem1_carry__0_n_2;
  wire rem1_carry__0_n_3;
  wire rem1_carry__1_i_1_n_0;
  wire rem1_carry__1_i_2_n_0;
  wire rem1_carry__1_i_3_n_0;
  wire rem1_carry__1_i_4_n_0;
  wire rem1_carry__1_n_0;
  wire rem1_carry__1_n_1;
  wire rem1_carry__1_n_2;
  wire rem1_carry__1_n_3;
  wire rem1_carry__2_i_1_n_0;
  wire rem1_carry__2_i_2_n_0;
  wire rem1_carry__2_i_3_n_0;
  wire rem1_carry__2_i_4_n_0;
  wire rem1_carry__2_n_0;
  wire rem1_carry__2_n_1;
  wire rem1_carry__2_n_2;
  wire rem1_carry__2_n_3;
  wire rem1_carry__3_i_1_n_0;
  wire rem1_carry__3_i_2_n_0;
  wire rem1_carry__3_i_3_n_0;
  wire rem1_carry__3_i_4_n_0;
  wire rem1_carry__3_n_0;
  wire rem1_carry__3_n_1;
  wire rem1_carry__3_n_2;
  wire rem1_carry__3_n_3;
  wire rem1_carry__4_i_1_n_0;
  wire rem1_carry__4_i_2_n_0;
  wire rem1_carry__4_i_3_n_0;
  wire rem1_carry__4_i_4_n_0;
  wire rem1_carry__4_n_0;
  wire rem1_carry__4_n_1;
  wire rem1_carry__4_n_2;
  wire rem1_carry__4_n_3;
  wire rem1_carry__5_i_1_n_0;
  wire rem1_carry__5_i_2_n_0;
  wire rem1_carry__5_i_3_n_0;
  wire rem1_carry__5_i_4_n_0;
  wire rem1_carry__5_n_0;
  wire rem1_carry__5_n_1;
  wire rem1_carry__5_n_2;
  wire rem1_carry__5_n_3;
  wire rem1_carry__6_i_1_n_0;
  wire rem1_carry__6_i_2_n_0;
  wire rem1_carry__6_i_3_n_0;
  wire rem1_carry__6_i_4_n_0;
  wire rem1_carry__6_n_0;
  wire rem1_carry__6_n_1;
  wire rem1_carry__6_n_2;
  wire rem1_carry__6_n_3;
  wire [0:0]rem1_carry__7_i_1_0;
  wire rem1_carry__7_i_1_n_0;
  wire rem1_carry_i_1_n_0;
  wire rem1_carry_i_2_n_0;
  wire rem1_carry_i_3_n_0;
  wire rem1_carry_i_4_n_0;
  wire rem1_carry_n_0;
  wire rem1_carry_n_1;
  wire rem1_carry_n_2;
  wire rem1_carry_n_3;
  wire [32:1]rem2;
  wire [3:0]rem2_carry__0_0;
  wire [3:0]rem2_carry__0_1;
  wire rem2_carry__0_i_1_n_0;
  wire rem2_carry__0_i_2_n_0;
  wire rem2_carry__0_i_3_n_0;
  wire rem2_carry__0_i_4_n_0;
  wire rem2_carry__0_n_0;
  wire rem2_carry__0_n_1;
  wire rem2_carry__0_n_2;
  wire rem2_carry__0_n_3;
  wire [3:0]rem2_carry__1_0;
  wire [3:0]rem2_carry__1_1;
  wire rem2_carry__1_i_1_n_0;
  wire rem2_carry__1_i_2_n_0;
  wire rem2_carry__1_i_3_n_0;
  wire rem2_carry__1_i_4_n_0;
  wire rem2_carry__1_n_0;
  wire rem2_carry__1_n_1;
  wire rem2_carry__1_n_2;
  wire rem2_carry__1_n_3;
  wire [3:0]rem2_carry__2_0;
  wire [3:0]rem2_carry__2_1;
  wire rem2_carry__2_i_1_n_0;
  wire rem2_carry__2_i_2_n_0;
  wire rem2_carry__2_i_3_n_0;
  wire rem2_carry__2_i_4_n_0;
  wire rem2_carry__2_n_0;
  wire rem2_carry__2_n_1;
  wire rem2_carry__2_n_2;
  wire rem2_carry__2_n_3;
  wire [3:0]rem2_carry__3_0;
  wire [3:0]rem2_carry__3_1;
  wire rem2_carry__3_i_1_n_0;
  wire rem2_carry__3_i_2_n_0;
  wire rem2_carry__3_i_3_n_0;
  wire rem2_carry__3_i_4_n_0;
  wire rem2_carry__3_n_0;
  wire rem2_carry__3_n_1;
  wire rem2_carry__3_n_2;
  wire rem2_carry__3_n_3;
  wire [3:0]rem2_carry__4_0;
  wire [3:0]rem2_carry__4_1;
  wire rem2_carry__4_i_1_n_0;
  wire rem2_carry__4_i_2_n_0;
  wire rem2_carry__4_i_3_n_0;
  wire rem2_carry__4_i_4_n_0;
  wire rem2_carry__4_n_0;
  wire rem2_carry__4_n_1;
  wire rem2_carry__4_n_2;
  wire rem2_carry__4_n_3;
  wire [3:0]rem2_carry__5_0;
  wire [3:0]rem2_carry__5_1;
  wire rem2_carry__5_i_1_n_0;
  wire rem2_carry__5_i_2_n_0;
  wire rem2_carry__5_i_3_n_0;
  wire rem2_carry__5_i_4_n_0;
  wire rem2_carry__5_n_0;
  wire rem2_carry__5_n_1;
  wire rem2_carry__5_n_2;
  wire rem2_carry__5_n_3;
  wire [3:0]rem2_carry__6_0;
  wire [3:0]rem2_carry__6_1;
  wire rem2_carry__6_i_1_n_0;
  wire rem2_carry__6_i_2_n_0;
  wire rem2_carry__6_i_3_n_0;
  wire rem2_carry__6_i_4_n_0;
  wire rem2_carry__6_n_0;
  wire rem2_carry__6_n_1;
  wire rem2_carry__6_n_2;
  wire rem2_carry__6_n_3;
  wire [0:0]rem2_carry__7_i_1_0;
  wire rem2_carry__7_i_1_n_0;
  wire rem2_carry_i_2_n_0;
  wire rem2_carry_i_3_n_0;
  wire rem2_carry_i_4_n_0;
  wire rem2_carry_n_0;
  wire rem2_carry_n_1;
  wire rem2_carry_n_2;
  wire rem2_carry_n_3;
  wire [32:1]rem3;
  wire rem3_carry__0_n_0;
  wire rem3_carry__0_n_1;
  wire rem3_carry__0_n_2;
  wire rem3_carry__0_n_3;
  wire rem3_carry__1_n_0;
  wire rem3_carry__1_n_1;
  wire rem3_carry__1_n_2;
  wire rem3_carry__1_n_3;
  wire rem3_carry__2_n_0;
  wire rem3_carry__2_n_1;
  wire rem3_carry__2_n_2;
  wire rem3_carry__2_n_3;
  wire rem3_carry__3_n_0;
  wire rem3_carry__3_n_1;
  wire rem3_carry__3_n_2;
  wire rem3_carry__3_n_3;
  wire rem3_carry__4_n_0;
  wire rem3_carry__4_n_1;
  wire rem3_carry__4_n_2;
  wire rem3_carry__4_n_3;
  wire rem3_carry__5_n_0;
  wire rem3_carry__5_n_1;
  wire rem3_carry__5_n_2;
  wire rem3_carry__5_n_3;
  wire rem3_carry__6_n_0;
  wire rem3_carry__6_n_1;
  wire rem3_carry__6_n_2;
  wire rem3_carry__6_n_3;
  wire rem3_carry_n_0;
  wire rem3_carry_n_1;
  wire rem3_carry_n_2;
  wire rem3_carry_n_3;
  wire \remden_reg[35] ;
  wire [0:0]\remden_reg[35]_0 ;

  GND GND
       (.G(\<const0> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry
       (.CI(\<const0> ),
        .CO({rem0_carry_n_0,rem0_carry_n_1,rem0_carry_n_2,rem0_carry_n_3}),
        .CYINIT(rem0_carry_i_1_n_0),
        .DI({rem1[3:1],\remden_reg[35] }),
        .O(fdiv_rem[3:0]),
        .S({rem0_carry_i_2_n_0,rem0_carry_i_3_n_0,rem0_carry_i_4_n_0,\remden_reg[35]_0 }));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__0
       (.CI(rem0_carry_n_0),
        .CO({rem0_carry__0_n_0,rem0_carry__0_n_1,rem0_carry__0_n_2,rem0_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1[7:4]),
        .O(fdiv_rem[7:4]),
        .S({rem0_carry__0_i_1_n_0,rem0_carry__0_i_2_n_0,rem0_carry__0_i_3_n_0,rem0_carry__0_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_1
       (.I0(rem1[7]),
        .I1(Q[6]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_2
       (.I0(rem1[6]),
        .I1(Q[5]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_3
       (.I0(rem1[5]),
        .I1(Q[4]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__0_i_4
       (.I0(rem1[4]),
        .I1(Q[3]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__0_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__1
       (.CI(rem0_carry__0_n_0),
        .CO({rem0_carry__1_n_0,rem0_carry__1_n_1,rem0_carry__1_n_2,rem0_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1[11:8]),
        .O(fdiv_rem[11:8]),
        .S({rem0_carry__1_i_1_n_0,rem0_carry__1_i_2_n_0,rem0_carry__1_i_3_n_0,rem0_carry__1_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_1
       (.I0(rem1[11]),
        .I1(Q[10]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_2
       (.I0(rem1[10]),
        .I1(Q[9]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_3
       (.I0(rem1[9]),
        .I1(Q[8]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__1_i_4
       (.I0(rem1[8]),
        .I1(Q[7]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__1_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__2
       (.CI(rem0_carry__1_n_0),
        .CO({rem0_carry__2_n_0,rem0_carry__2_n_1,rem0_carry__2_n_2,rem0_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1[15:12]),
        .O(fdiv_rem[15:12]),
        .S({rem0_carry__2_i_1_n_0,rem0_carry__2_i_2_n_0,rem0_carry__2_i_3_n_0,rem0_carry__2_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_1
       (.I0(rem1[15]),
        .I1(rem1_carry__7_i_1_0),
        .I2(Q[14]),
        .O(rem0_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_2
       (.I0(rem1[14]),
        .I1(Q[13]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_3
       (.I0(rem1[13]),
        .I1(Q[12]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__2_i_4
       (.I0(rem1[12]),
        .I1(Q[11]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__2_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__3
       (.CI(rem0_carry__2_n_0),
        .CO({rem0_carry__3_n_0,rem0_carry__3_n_1,rem0_carry__3_n_2,rem0_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1[19:16]),
        .O(fdiv_rem[19:16]),
        .S({rem0_carry__3_i_1_n_0,rem0_carry__3_i_2_n_0,rem0_carry__3_i_3_n_0,rem0_carry__3_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_1
       (.I0(rem1[19]),
        .I1(Q[18]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_2
       (.I0(rem1[18]),
        .I1(Q[17]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_3
       (.I0(rem1[17]),
        .I1(Q[16]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__3_i_4
       (.I0(rem1[16]),
        .I1(Q[15]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__3_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__4
       (.CI(rem0_carry__3_n_0),
        .CO({rem0_carry__4_n_0,rem0_carry__4_n_1,rem0_carry__4_n_2,rem0_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1[23:20]),
        .O(fdiv_rem[23:20]),
        .S({rem0_carry__4_i_1_n_0,rem0_carry__4_i_2_n_0,rem0_carry__4_i_3_n_0,rem0_carry__4_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_1
       (.I0(rem1[23]),
        .I1(Q[22]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_2
       (.I0(rem1[22]),
        .I1(Q[21]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_3
       (.I0(rem1[21]),
        .I1(Q[20]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__4_i_4
       (.I0(rem1[20]),
        .I1(Q[19]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__4_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__5
       (.CI(rem0_carry__4_n_0),
        .CO({rem0_carry__5_n_0,rem0_carry__5_n_1,rem0_carry__5_n_2,rem0_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1[27:24]),
        .O(fdiv_rem[27:24]),
        .S({rem0_carry__5_i_1_n_0,rem0_carry__5_i_2_n_0,rem0_carry__5_i_3_n_0,rem0_carry__5_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_1
       (.I0(rem1[27]),
        .I1(Q[26]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_2
       (.I0(rem1[26]),
        .I1(Q[25]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_3
       (.I0(rem1[25]),
        .I1(Q[24]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__5_i_4
       (.I0(rem1[24]),
        .I1(Q[23]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__5_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__6
       (.CI(rem0_carry__5_n_0),
        .CO({rem0_carry__6_n_0,rem0_carry__6_n_1,rem0_carry__6_n_2,rem0_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem1[31:28]),
        .O(fdiv_rem[31:28]),
        .S({rem0_carry__6_i_1_n_0,rem0_carry__6_i_2_n_0,rem0_carry__6_i_3_n_0,rem0_carry__6_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_1
       (.I0(rem1[31]),
        .I1(rem1_carry__7_i_1_0),
        .I2(Q[30]),
        .O(rem0_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_2
       (.I0(rem1[30]),
        .I1(Q[29]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_3
       (.I0(rem1[29]),
        .I1(Q[28]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry__6_i_4
       (.I0(rem1[28]),
        .I1(Q[27]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry__6_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem0_carry__7
       (.CI(rem0_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(rem0_carry__7_i_1_0),
        .S({\<const0> ,\<const0> ,\<const0> ,rem0_carry__7_i_1_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem0_carry__7_i_1
       (.I0(rem1_carry__7_i_1_0),
        .I1(rem1[32]),
        .O(rem0_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem0_carry_i_1
       (.I0(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_2
       (.I0(rem1[3]),
        .I1(Q[2]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_3
       (.I0(rem1[2]),
        .I1(Q[1]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_4
       (.I0(rem1[1]),
        .I1(Q[0]),
        .I2(rem1_carry__7_i_1_0),
        .O(rem0_carry_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry
       (.CI(\<const0> ),
        .CO({rem1_carry_n_0,rem1_carry_n_1,rem1_carry_n_2,rem1_carry_n_3}),
        .CYINIT(rem1_carry_i_1_n_0),
        .DI({rem2[3:1],rem0_carry_0}),
        .O(rem1[4:1]),
        .S({rem1_carry_i_2_n_0,rem1_carry_i_3_n_0,rem1_carry_i_4_n_0,rem0_carry_1}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__0
       (.CI(rem1_carry_n_0),
        .CO({rem1_carry__0_n_0,rem1_carry__0_n_1,rem1_carry__0_n_2,rem1_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2[7:4]),
        .O(rem1[8:5]),
        .S({rem1_carry__0_i_1_n_0,rem1_carry__0_i_2_n_0,rem1_carry__0_i_3_n_0,rem1_carry__0_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_1
       (.I0(rem2[7]),
        .I1(Q[6]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_2
       (.I0(rem2[6]),
        .I1(Q[5]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_3
       (.I0(rem2[5]),
        .I1(Q[4]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__0_i_4
       (.I0(rem2[4]),
        .I1(Q[3]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__0_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__1
       (.CI(rem1_carry__0_n_0),
        .CO({rem1_carry__1_n_0,rem1_carry__1_n_1,rem1_carry__1_n_2,rem1_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2[11:8]),
        .O(rem1[12:9]),
        .S({rem1_carry__1_i_1_n_0,rem1_carry__1_i_2_n_0,rem1_carry__1_i_3_n_0,rem1_carry__1_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_1
       (.I0(rem2[11]),
        .I1(Q[10]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_2
       (.I0(rem2[10]),
        .I1(Q[9]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_3
       (.I0(rem2[9]),
        .I1(Q[8]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__1_i_4
       (.I0(rem2[8]),
        .I1(Q[7]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__1_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__2
       (.CI(rem1_carry__1_n_0),
        .CO({rem1_carry__2_n_0,rem1_carry__2_n_1,rem1_carry__2_n_2,rem1_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2[15:12]),
        .O(rem1[16:13]),
        .S({rem1_carry__2_i_1_n_0,rem1_carry__2_i_2_n_0,rem1_carry__2_i_3_n_0,rem1_carry__2_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_1
       (.I0(rem2[15]),
        .I1(rem2_carry__7_i_1_0),
        .I2(Q[14]),
        .O(rem1_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_2
       (.I0(rem2[14]),
        .I1(Q[13]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_3
       (.I0(rem2[13]),
        .I1(Q[12]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__2_i_4
       (.I0(rem2[12]),
        .I1(Q[11]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__2_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__3
       (.CI(rem1_carry__2_n_0),
        .CO({rem1_carry__3_n_0,rem1_carry__3_n_1,rem1_carry__3_n_2,rem1_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2[19:16]),
        .O(rem1[20:17]),
        .S({rem1_carry__3_i_1_n_0,rem1_carry__3_i_2_n_0,rem1_carry__3_i_3_n_0,rem1_carry__3_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_1
       (.I0(rem2[19]),
        .I1(Q[18]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_2
       (.I0(rem2[18]),
        .I1(Q[17]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_3
       (.I0(rem2[17]),
        .I1(Q[16]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__3_i_4
       (.I0(rem2[16]),
        .I1(Q[15]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__3_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__4
       (.CI(rem1_carry__3_n_0),
        .CO({rem1_carry__4_n_0,rem1_carry__4_n_1,rem1_carry__4_n_2,rem1_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2[23:20]),
        .O(rem1[24:21]),
        .S({rem1_carry__4_i_1_n_0,rem1_carry__4_i_2_n_0,rem1_carry__4_i_3_n_0,rem1_carry__4_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_1
       (.I0(rem2[23]),
        .I1(Q[22]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_2
       (.I0(rem2[22]),
        .I1(Q[21]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_3
       (.I0(rem2[21]),
        .I1(Q[20]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__4_i_4
       (.I0(rem2[20]),
        .I1(Q[19]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__4_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__5
       (.CI(rem1_carry__4_n_0),
        .CO({rem1_carry__5_n_0,rem1_carry__5_n_1,rem1_carry__5_n_2,rem1_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2[27:24]),
        .O(rem1[28:25]),
        .S({rem1_carry__5_i_1_n_0,rem1_carry__5_i_2_n_0,rem1_carry__5_i_3_n_0,rem1_carry__5_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_1
       (.I0(rem2[27]),
        .I1(Q[26]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_2
       (.I0(rem2[26]),
        .I1(Q[25]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_3
       (.I0(rem2[25]),
        .I1(Q[24]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__5_i_4
       (.I0(rem2[24]),
        .I1(Q[23]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__5_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__6
       (.CI(rem1_carry__5_n_0),
        .CO({rem1_carry__6_n_0,rem1_carry__6_n_1,rem1_carry__6_n_2,rem1_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2[31:28]),
        .O(rem1[32:29]),
        .S({rem1_carry__6_i_1_n_0,rem1_carry__6_i_2_n_0,rem1_carry__6_i_3_n_0,rem1_carry__6_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_1
       (.I0(rem2[31]),
        .I1(rem2_carry__7_i_1_0),
        .I2(Q[30]),
        .O(rem1_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_2
       (.I0(rem2[30]),
        .I1(Q[29]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_3
       (.I0(rem2[29]),
        .I1(Q[28]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry__6_i_4
       (.I0(rem2[28]),
        .I1(Q[27]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry__6_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem1_carry__7
       (.CI(rem1_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(rem1_carry__7_i_1_0),
        .S({\<const0> ,\<const0> ,\<const0> ,rem1_carry__7_i_1_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem1_carry__7_i_1
       (.I0(rem2_carry__7_i_1_0),
        .I1(rem2[32]),
        .O(rem1_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem1_carry_i_1
       (.I0(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_2
       (.I0(rem2[3]),
        .I1(Q[2]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_3
       (.I0(rem2[2]),
        .I1(Q[1]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_4
       (.I0(rem2[1]),
        .I1(Q[0]),
        .I2(rem2_carry__7_i_1_0),
        .O(rem1_carry_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry
       (.CI(\<const0> ),
        .CO({rem2_carry_n_0,rem2_carry_n_1,rem2_carry_n_2,rem2_carry_n_3}),
        .CYINIT(p_1_in3_in),
        .DI({rem3[3:1],rem1_carry_0}),
        .O(rem2[4:1]),
        .S({rem2_carry_i_2_n_0,rem2_carry_i_3_n_0,rem2_carry_i_4_n_0,rem1_carry_1}));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__0
       (.CI(rem2_carry_n_0),
        .CO({rem2_carry__0_n_0,rem2_carry__0_n_1,rem2_carry__0_n_2,rem2_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3[7:4]),
        .O(rem2[8:5]),
        .S({rem2_carry__0_i_1_n_0,rem2_carry__0_i_2_n_0,rem2_carry__0_i_3_n_0,rem2_carry__0_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_1
       (.I0(rem3[7]),
        .I1(Q[6]),
        .I2(O),
        .O(rem2_carry__0_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_2
       (.I0(rem3[6]),
        .I1(Q[5]),
        .I2(O),
        .O(rem2_carry__0_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_3
       (.I0(rem3[5]),
        .I1(Q[4]),
        .I2(O),
        .O(rem2_carry__0_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__0_i_4
       (.I0(rem3[4]),
        .I1(Q[3]),
        .I2(O),
        .O(rem2_carry__0_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__1
       (.CI(rem2_carry__0_n_0),
        .CO({rem2_carry__1_n_0,rem2_carry__1_n_1,rem2_carry__1_n_2,rem2_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3[11:8]),
        .O(rem2[12:9]),
        .S({rem2_carry__1_i_1_n_0,rem2_carry__1_i_2_n_0,rem2_carry__1_i_3_n_0,rem2_carry__1_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_1
       (.I0(rem3[11]),
        .I1(Q[10]),
        .I2(O),
        .O(rem2_carry__1_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_2
       (.I0(rem3[10]),
        .I1(Q[9]),
        .I2(O),
        .O(rem2_carry__1_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_3
       (.I0(rem3[9]),
        .I1(Q[8]),
        .I2(O),
        .O(rem2_carry__1_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__1_i_4
       (.I0(rem3[8]),
        .I1(Q[7]),
        .I2(O),
        .O(rem2_carry__1_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__2
       (.CI(rem2_carry__1_n_0),
        .CO({rem2_carry__2_n_0,rem2_carry__2_n_1,rem2_carry__2_n_2,rem2_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3[15:12]),
        .O(rem2[16:13]),
        .S({rem2_carry__2_i_1_n_0,rem2_carry__2_i_2_n_0,rem2_carry__2_i_3_n_0,rem2_carry__2_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_1
       (.I0(rem3[15]),
        .I1(O),
        .I2(Q[14]),
        .O(rem2_carry__2_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_2
       (.I0(rem3[14]),
        .I1(Q[13]),
        .I2(O),
        .O(rem2_carry__2_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_3
       (.I0(rem3[13]),
        .I1(Q[12]),
        .I2(O),
        .O(rem2_carry__2_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__2_i_4
       (.I0(rem3[12]),
        .I1(Q[11]),
        .I2(O),
        .O(rem2_carry__2_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__3
       (.CI(rem2_carry__2_n_0),
        .CO({rem2_carry__3_n_0,rem2_carry__3_n_1,rem2_carry__3_n_2,rem2_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3[19:16]),
        .O(rem2[20:17]),
        .S({rem2_carry__3_i_1_n_0,rem2_carry__3_i_2_n_0,rem2_carry__3_i_3_n_0,rem2_carry__3_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_1
       (.I0(rem3[19]),
        .I1(Q[18]),
        .I2(O),
        .O(rem2_carry__3_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_2
       (.I0(rem3[18]),
        .I1(Q[17]),
        .I2(O),
        .O(rem2_carry__3_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_3
       (.I0(rem3[17]),
        .I1(Q[16]),
        .I2(O),
        .O(rem2_carry__3_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__3_i_4
       (.I0(rem3[16]),
        .I1(Q[15]),
        .I2(O),
        .O(rem2_carry__3_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__4
       (.CI(rem2_carry__3_n_0),
        .CO({rem2_carry__4_n_0,rem2_carry__4_n_1,rem2_carry__4_n_2,rem2_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3[23:20]),
        .O(rem2[24:21]),
        .S({rem2_carry__4_i_1_n_0,rem2_carry__4_i_2_n_0,rem2_carry__4_i_3_n_0,rem2_carry__4_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_1
       (.I0(rem3[23]),
        .I1(Q[22]),
        .I2(O),
        .O(rem2_carry__4_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_2
       (.I0(rem3[22]),
        .I1(Q[21]),
        .I2(O),
        .O(rem2_carry__4_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_3
       (.I0(rem3[21]),
        .I1(Q[20]),
        .I2(O),
        .O(rem2_carry__4_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__4_i_4
       (.I0(rem3[20]),
        .I1(Q[19]),
        .I2(O),
        .O(rem2_carry__4_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__5
       (.CI(rem2_carry__4_n_0),
        .CO({rem2_carry__5_n_0,rem2_carry__5_n_1,rem2_carry__5_n_2,rem2_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3[27:24]),
        .O(rem2[28:25]),
        .S({rem2_carry__5_i_1_n_0,rem2_carry__5_i_2_n_0,rem2_carry__5_i_3_n_0,rem2_carry__5_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_1
       (.I0(rem3[27]),
        .I1(Q[26]),
        .I2(O),
        .O(rem2_carry__5_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_2
       (.I0(rem3[26]),
        .I1(Q[25]),
        .I2(O),
        .O(rem2_carry__5_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_3
       (.I0(rem3[25]),
        .I1(Q[24]),
        .I2(O),
        .O(rem2_carry__5_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__5_i_4
       (.I0(rem3[24]),
        .I1(Q[23]),
        .I2(O),
        .O(rem2_carry__5_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__6
       (.CI(rem2_carry__5_n_0),
        .CO({rem2_carry__6_n_0,rem2_carry__6_n_1,rem2_carry__6_n_2,rem2_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem3[31:28]),
        .O(rem2[32:29]),
        .S({rem2_carry__6_i_1_n_0,rem2_carry__6_i_2_n_0,rem2_carry__6_i_3_n_0,rem2_carry__6_i_4_n_0}));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_1
       (.I0(rem3[31]),
        .I1(O),
        .I2(Q[30]),
        .O(rem2_carry__6_i_1_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_2
       (.I0(rem3[30]),
        .I1(Q[29]),
        .I2(O),
        .O(rem2_carry__6_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_3
       (.I0(rem3[29]),
        .I1(Q[28]),
        .I2(O),
        .O(rem2_carry__6_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry__6_i_4
       (.I0(rem3[28]),
        .I1(Q[27]),
        .I2(O),
        .O(rem2_carry__6_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem2_carry__7
       (.CI(rem2_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(rem2_carry__7_i_1_0),
        .S({\<const0> ,\<const0> ,\<const0> ,rem2_carry__7_i_1_n_0}));
  LUT2 #(
    .INIT(4'h9)) 
    rem2_carry__7_i_1
       (.I0(O),
        .I1(rem3[32]),
        .O(rem2_carry__7_i_1_n_0));
  LUT1 #(
    .INIT(2'h1)) 
    rem2_carry_i_1
       (.I0(O),
        .O(p_1_in3_in));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_2
       (.I0(rem3[3]),
        .I1(Q[2]),
        .I2(O),
        .O(rem2_carry_i_2_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_3
       (.I0(rem3[2]),
        .I1(Q[1]),
        .I2(O),
        .O(rem2_carry_i_3_n_0));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_4
       (.I0(rem3[1]),
        .I1(Q[0]),
        .I2(O),
        .O(rem2_carry_i_4_n_0));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry
       (.CI(\<const0> ),
        .CO({rem3_carry_n_0,rem3_carry_n_1,rem3_carry_n_2,rem3_carry_n_3}),
        .CYINIT(p_1_in5_in),
        .DI(DI),
        .O(rem3[4:1]),
        .S(S));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__0
       (.CI(rem3_carry_n_0),
        .CO({rem3_carry__0_n_0,rem3_carry__0_n_1,rem3_carry__0_n_2,rem3_carry__0_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2_carry__0_0),
        .O(rem3[8:5]),
        .S(rem2_carry__0_1));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__1
       (.CI(rem3_carry__0_n_0),
        .CO({rem3_carry__1_n_0,rem3_carry__1_n_1,rem3_carry__1_n_2,rem3_carry__1_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2_carry__1_0),
        .O(rem3[12:9]),
        .S(rem2_carry__1_1));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__2
       (.CI(rem3_carry__1_n_0),
        .CO({rem3_carry__2_n_0,rem3_carry__2_n_1,rem3_carry__2_n_2,rem3_carry__2_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2_carry__2_0),
        .O(rem3[16:13]),
        .S(rem2_carry__2_1));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__3
       (.CI(rem3_carry__2_n_0),
        .CO({rem3_carry__3_n_0,rem3_carry__3_n_1,rem3_carry__3_n_2,rem3_carry__3_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2_carry__3_0),
        .O(rem3[20:17]),
        .S(rem2_carry__3_1));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__4
       (.CI(rem3_carry__3_n_0),
        .CO({rem3_carry__4_n_0,rem3_carry__4_n_1,rem3_carry__4_n_2,rem3_carry__4_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2_carry__4_0),
        .O(rem3[24:21]),
        .S(rem2_carry__4_1));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__5
       (.CI(rem3_carry__4_n_0),
        .CO({rem3_carry__5_n_0,rem3_carry__5_n_1,rem3_carry__5_n_2,rem3_carry__5_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2_carry__5_0),
        .O(rem3[28:25]),
        .S(rem2_carry__5_1));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__6
       (.CI(rem3_carry__5_n_0),
        .CO({rem3_carry__6_n_0,rem3_carry__6_n_1,rem3_carry__6_n_2,rem3_carry__6_n_3}),
        .CYINIT(\<const0> ),
        .DI(rem2_carry__6_0),
        .O(rem3[32:29]),
        .S(rem2_carry__6_1));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 rem3_carry__7
       (.CI(rem3_carry__6_n_0),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(O),
        .S({\<const0> ,\<const0> ,\<const0> ,\quo_reg[3] }));
endmodule

module niho_div_fsm
   (\sr_reg[8] ,
    \dctl_stat_reg[3]_0 ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \dctl_stat_reg[2]_0 ,
    \dctl_stat_reg[1]_0 ,
    E,
    D,
    div_crdy_reg,
    dctl_long,
    \dctl_stat_reg[2]_1 ,
    \rem_reg[3] ,
    \dso_reg[31] ,
    S,
    div_crdy_reg_0,
    rst_n_0,
    \rem_reg[30] ,
    \rem_reg[27] ,
    \rem_reg[23] ,
    \rem_reg[19] ,
    \rem_reg[15] ,
    \rem_reg[11] ,
    \rem_reg[7] ,
    \rem_reg[27]_0 ,
    \rem_reg[23]_0 ,
    \rem_reg[19]_0 ,
    \rem_reg[15]_0 ,
    \rem_reg[11]_0 ,
    \rem_reg[7]_0 ,
    rst_n_1,
    rst_n_2,
    rst_n_3,
    rst_n_4,
    rst_n_5,
    rst_n_6,
    rst_n_7,
    rst_n_8,
    rst_n_9,
    rst_n_10,
    rst_n_11,
    rst_n_12,
    rst_n_13,
    rst_n_14,
    rst_n_15,
    rst_n_16,
    rst_n_17,
    rst_n_18,
    rst_n_19,
    rst_n_20,
    rst_n_21,
    rst_n_22,
    rst_n_23,
    rst_n_24,
    rst_n_25,
    rst_n_26,
    rst_n_27,
    rst_n_28,
    rst_n_29,
    \remden_reg[28] ,
    \remden_reg[28]_0 ,
    \remden_reg[28]_1 ,
    \remden_reg[28]_2 ,
    rst_n_30,
    rst_n_31,
    rst_n_32,
    rst_n_33,
    rst_n_34,
    rst_n_35,
    rst_n_36,
    rst_n_37,
    \rem_reg[31] ,
    \sr_reg[8]_11 ,
    p_0_in,
    fdiv_rem_msb_f_reg_0,
    clk,
    \remden_reg[31] ,
    abus_0,
    rgf_sr_nh,
    \remden_reg[15] ,
    \remden_reg[0] ,
    \remden_reg[14] ,
    \remden_reg[13] ,
    \remden_reg[12] ,
    \remden_reg[11] ,
    \remden_reg[10] ,
    \remden_reg[9] ,
    \remden_reg[8] ,
    \remden_reg[7] ,
    \remden_reg[6] ,
    \remden_reg[5] ,
    \remden_reg[4] ,
    dctl_sign,
    Q,
    add_out0_carry__6,
    add_out0_carry__2_i_11_0,
    add_out0_carry__2_i_9_0,
    add_out0_carry__4_i_10_0,
    add_out0_carry__4_i_9_0,
    add_out0_carry__5_i_12_0,
    add_out0_carry__5_i_10_0,
    DI,
    add_out0_carry__6_i_9_0,
    add_out0_carry__6_i_10_0,
    add_out0_carry__5_i_11_0,
    add_out0_carry__4_i_11_0,
    add_out0_carry__4_i_12_0,
    add_out0_carry__3_i_9_0,
    add_out0_carry__3_i_10_0,
    add_out0_carry__3_i_11_0,
    add_out0_carry__3_i_12_0,
    add_out0_carry__2_i_12_0,
    \rem_reg[31]_0 ,
    add_out0_carry__2_i_10_0,
    \remden_reg[31]_0 ,
    dctl_long_f_reg,
    dctl_long_f_reg_0,
    den2,
    \dctl_stat_reg[3]_1 ,
    chg_quo_sgn_reg_0,
    \dctl_stat_reg[2]_2 ,
    \remden_reg[64] ,
    chg_rem_sgn0,
    rst_n,
    fdiv_rem,
    \dso_reg[19] ,
    \dso_reg[19]_0 ,
    \dso_reg[19]_1 ,
    \dso_reg[19]_2 ,
    \dso_reg[23] ,
    \dso_reg[23]_0 ,
    \dso_reg[23]_1 ,
    \dso_reg[23]_2 ,
    \dso_reg[27] ,
    \dso_reg[27]_0 ,
    \dso_reg[27]_1 ,
    \dso_reg[27]_2 ,
    \dso_reg[31]_0 ,
    \dso_reg[31]_1 ,
    \dso_reg[31]_2 ,
    \dso_reg[31]_3 ,
    \remden_reg[31]_1 ,
    \remden_reg[29] ,
    \remden_reg[30] ,
    \remden_reg[19] ,
    bbus_0);
  output \sr_reg[8] ;
  output \dctl_stat_reg[3]_0 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \dctl_stat_reg[2]_0 ;
  output \dctl_stat_reg[1]_0 ;
  output [0:0]E;
  output [3:0]D;
  output [0:0]div_crdy_reg;
  output dctl_long;
  output [0:0]\dctl_stat_reg[2]_1 ;
  output [3:0]\rem_reg[3] ;
  output [3:0]\dso_reg[31] ;
  output [3:0]S;
  output div_crdy_reg_0;
  output rst_n_0;
  output [2:0]\rem_reg[30] ;
  output [3:0]\rem_reg[27] ;
  output [3:0]\rem_reg[23] ;
  output [3:0]\rem_reg[19] ;
  output [3:0]\rem_reg[15] ;
  output [3:0]\rem_reg[11] ;
  output [3:0]\rem_reg[7] ;
  output [3:0]\rem_reg[27]_0 ;
  output [3:0]\rem_reg[23]_0 ;
  output [3:0]\rem_reg[19]_0 ;
  output [3:0]\rem_reg[15]_0 ;
  output [3:0]\rem_reg[11]_0 ;
  output [3:0]\rem_reg[7]_0 ;
  output rst_n_1;
  output rst_n_2;
  output rst_n_3;
  output rst_n_4;
  output rst_n_5;
  output rst_n_6;
  output rst_n_7;
  output rst_n_8;
  output rst_n_9;
  output rst_n_10;
  output rst_n_11;
  output rst_n_12;
  output rst_n_13;
  output rst_n_14;
  output rst_n_15;
  output rst_n_16;
  output rst_n_17;
  output rst_n_18;
  output rst_n_19;
  output rst_n_20;
  output rst_n_21;
  output rst_n_22;
  output rst_n_23;
  output rst_n_24;
  output rst_n_25;
  output rst_n_26;
  output rst_n_27;
  output rst_n_28;
  output rst_n_29;
  output \remden_reg[28] ;
  output \remden_reg[28]_0 ;
  output \remden_reg[28]_1 ;
  output \remden_reg[28]_2 ;
  output rst_n_30;
  output rst_n_31;
  output rst_n_32;
  output rst_n_33;
  output rst_n_34;
  output rst_n_35;
  output rst_n_36;
  output rst_n_37;
  output [31:0]\rem_reg[31] ;
  output [31:0]\sr_reg[8]_11 ;
  input p_0_in;
  input [0:0]fdiv_rem_msb_f_reg_0;
  input clk;
  input [20:0]\remden_reg[31] ;
  input [15:0]abus_0;
  input rgf_sr_nh;
  input \remden_reg[15] ;
  input \remden_reg[0] ;
  input \remden_reg[14] ;
  input \remden_reg[13] ;
  input \remden_reg[12] ;
  input \remden_reg[11] ;
  input \remden_reg[10] ;
  input \remden_reg[9] ;
  input \remden_reg[8] ;
  input \remden_reg[7] ;
  input \remden_reg[6] ;
  input \remden_reg[5] ;
  input \remden_reg[4] ;
  input dctl_sign;
  input [31:0]Q;
  input [31:0]add_out0_carry__6;
  input add_out0_carry__2_i_11_0;
  input add_out0_carry__2_i_9_0;
  input add_out0_carry__4_i_10_0;
  input add_out0_carry__4_i_9_0;
  input add_out0_carry__5_i_12_0;
  input add_out0_carry__5_i_10_0;
  input [0:0]DI;
  input [0:0]add_out0_carry__6_i_9_0;
  input add_out0_carry__6_i_10_0;
  input add_out0_carry__5_i_11_0;
  input add_out0_carry__4_i_11_0;
  input add_out0_carry__4_i_12_0;
  input add_out0_carry__3_i_9_0;
  input add_out0_carry__3_i_10_0;
  input add_out0_carry__3_i_11_0;
  input add_out0_carry__3_i_12_0;
  input add_out0_carry__2_i_12_0;
  input [31:0]\rem_reg[31]_0 ;
  input add_out0_carry__2_i_10_0;
  input \remden_reg[31]_0 ;
  input dctl_long_f_reg;
  input dctl_long_f_reg_0;
  input [0:0]den2;
  input \dctl_stat_reg[3]_1 ;
  input chg_quo_sgn_reg_0;
  input \dctl_stat_reg[2]_2 ;
  input \remden_reg[64] ;
  input chg_rem_sgn0;
  input rst_n;
  input [31:0]fdiv_rem;
  input \dso_reg[19] ;
  input \dso_reg[19]_0 ;
  input \dso_reg[19]_1 ;
  input \dso_reg[19]_2 ;
  input \dso_reg[23] ;
  input \dso_reg[23]_0 ;
  input \dso_reg[23]_1 ;
  input \dso_reg[23]_2 ;
  input \dso_reg[27] ;
  input \dso_reg[27]_0 ;
  input \dso_reg[27]_1 ;
  input \dso_reg[27]_2 ;
  input \dso_reg[31]_0 ;
  input \dso_reg[31]_1 ;
  input \dso_reg[31]_2 ;
  input \dso_reg[31]_3 ;
  input \remden_reg[31]_1 ;
  input \remden_reg[29] ;
  input \remden_reg[30] ;
  input \remden_reg[19] ;
  input [15:0]bbus_0;

  wire \<const0> ;
  wire \<const1> ;
  wire [3:0]D;
  wire [0:0]DI;
  wire [0:0]E;
  wire [31:0]Q;
  wire [3:0]S;
  wire [15:0]abus_0;
  wire add_out0_carry__0_i_13_n_0;
  wire add_out0_carry__0_i_14_n_0;
  wire add_out0_carry__0_i_15_n_0;
  wire add_out0_carry__0_i_16_n_0;
  wire add_out0_carry__1_i_13_n_0;
  wire add_out0_carry__1_i_14_n_0;
  wire add_out0_carry__1_i_15_n_0;
  wire add_out0_carry__1_i_16_n_0;
  wire add_out0_carry__2_i_10_0;
  wire add_out0_carry__2_i_11_0;
  wire add_out0_carry__2_i_12_0;
  wire add_out0_carry__2_i_13_n_0;
  wire add_out0_carry__2_i_14_n_0;
  wire add_out0_carry__2_i_15_n_0;
  wire add_out0_carry__2_i_16_n_0;
  wire add_out0_carry__2_i_9_0;
  wire add_out0_carry__3_i_10_0;
  wire add_out0_carry__3_i_11_0;
  wire add_out0_carry__3_i_12_0;
  wire add_out0_carry__3_i_13_n_0;
  wire add_out0_carry__3_i_14_n_0;
  wire add_out0_carry__3_i_15_n_0;
  wire add_out0_carry__3_i_16_n_0;
  wire add_out0_carry__3_i_9_0;
  wire add_out0_carry__4_i_10_0;
  wire add_out0_carry__4_i_11_0;
  wire add_out0_carry__4_i_12_0;
  wire add_out0_carry__4_i_13_n_0;
  wire add_out0_carry__4_i_14_n_0;
  wire add_out0_carry__4_i_15_n_0;
  wire add_out0_carry__4_i_16_n_0;
  wire add_out0_carry__4_i_9_0;
  wire add_out0_carry__5_i_10_0;
  wire add_out0_carry__5_i_11_0;
  wire add_out0_carry__5_i_12_0;
  wire add_out0_carry__5_i_13_n_0;
  wire add_out0_carry__5_i_14_n_0;
  wire add_out0_carry__5_i_15_n_0;
  wire add_out0_carry__5_i_16_n_0;
  wire [31:0]add_out0_carry__6;
  wire add_out0_carry__6_i_10_0;
  wire add_out0_carry__6_i_11_n_0;
  wire add_out0_carry__6_i_12_n_0;
  wire add_out0_carry__6_i_13_n_0;
  wire [0:0]add_out0_carry__6_i_9_0;
  wire add_out0_carry_i_10_n_0;
  wire add_out0_carry_i_15_n_0;
  wire add_out0_carry_i_16_n_0;
  wire add_out0_carry_i_17_n_0;
  wire add_out0_carry_i_18_n_0;
  wire add_out0_carry_i_19_n_0;
  wire add_out0_carry_i_20_n_0;
  wire add_out0_carry_i_21_n_0;
  wire add_out0_carry_i_9_n_0;
  wire [15:0]bbus_0;
  wire chg_quo_sgn;
  wire chg_quo_sgn_i_1_n_0;
  wire chg_quo_sgn_reg_0;
  wire chg_rem_sgn;
  wire chg_rem_sgn0;
  wire chg_rem_sgn_i_1_n_0;
  wire clk;
  wire dctl_long;
  wire dctl_long_f_reg;
  wire dctl_long_f_reg_0;
  wire [3:0]dctl_next;
  wire dctl_sign;
  wire [3:0]dctl_stat;
  wire \dctl_stat[0]_i_2_n_0 ;
  wire \dctl_stat[0]_i_3_n_0 ;
  wire \dctl_stat[1]_i_2_n_0 ;
  wire \dctl_stat[1]_i_3_n_0 ;
  wire \dctl_stat[3]_i_4_n_0 ;
  wire \dctl_stat[3]_i_5_n_0 ;
  wire \dctl_stat_reg[1]_0 ;
  wire \dctl_stat_reg[2]_0 ;
  wire [0:0]\dctl_stat_reg[2]_1 ;
  wire \dctl_stat_reg[2]_2 ;
  wire \dctl_stat_reg[3]_0 ;
  wire \dctl_stat_reg[3]_1 ;
  wire [0:0]den2;
  wire div_crdy_i_2_n_0;
  wire div_crdy_i_3_n_0;
  wire div_crdy_i_4_n_0;
  wire [0:0]div_crdy_reg;
  wire div_crdy_reg_0;
  wire \dso[11]_i_10_n_0 ;
  wire \dso[11]_i_11_n_0 ;
  wire \dso[11]_i_12_n_0 ;
  wire \dso[11]_i_13_n_0 ;
  wire \dso[11]_i_2_n_0 ;
  wire \dso[11]_i_3_n_0 ;
  wire \dso[11]_i_4_n_0 ;
  wire \dso[11]_i_5_n_0 ;
  wire \dso[11]_i_6_n_0 ;
  wire \dso[11]_i_7_n_0 ;
  wire \dso[11]_i_8_n_0 ;
  wire \dso[11]_i_9_n_0 ;
  wire \dso[15]_i_10_n_0 ;
  wire \dso[15]_i_11_n_0 ;
  wire \dso[15]_i_12_n_0 ;
  wire \dso[15]_i_13_n_0 ;
  wire \dso[15]_i_14_n_0 ;
  wire \dso[15]_i_2_n_0 ;
  wire \dso[15]_i_3_n_0 ;
  wire \dso[15]_i_4_n_0 ;
  wire \dso[15]_i_5_n_0 ;
  wire \dso[15]_i_6_n_0 ;
  wire \dso[15]_i_7_n_0 ;
  wire \dso[15]_i_8_n_0 ;
  wire \dso[15]_i_9_n_0 ;
  wire \dso[19]_i_10_n_0 ;
  wire \dso[19]_i_11_n_0 ;
  wire \dso[19]_i_12_n_0 ;
  wire \dso[19]_i_13_n_0 ;
  wire \dso[19]_i_2_n_0 ;
  wire \dso[19]_i_3_n_0 ;
  wire \dso[19]_i_4_n_0 ;
  wire \dso[19]_i_5_n_0 ;
  wire \dso[19]_i_6_n_0 ;
  wire \dso[19]_i_7_n_0 ;
  wire \dso[19]_i_8_n_0 ;
  wire \dso[19]_i_9_n_0 ;
  wire \dso[23]_i_10_n_0 ;
  wire \dso[23]_i_11_n_0 ;
  wire \dso[23]_i_12_n_0 ;
  wire \dso[23]_i_13_n_0 ;
  wire \dso[23]_i_2_n_0 ;
  wire \dso[23]_i_3_n_0 ;
  wire \dso[23]_i_4_n_0 ;
  wire \dso[23]_i_5_n_0 ;
  wire \dso[23]_i_6_n_0 ;
  wire \dso[23]_i_7_n_0 ;
  wire \dso[23]_i_8_n_0 ;
  wire \dso[23]_i_9_n_0 ;
  wire \dso[27]_i_10_n_0 ;
  wire \dso[27]_i_11_n_0 ;
  wire \dso[27]_i_12_n_0 ;
  wire \dso[27]_i_13_n_0 ;
  wire \dso[27]_i_2_n_0 ;
  wire \dso[27]_i_3_n_0 ;
  wire \dso[27]_i_4_n_0 ;
  wire \dso[27]_i_5_n_0 ;
  wire \dso[27]_i_6_n_0 ;
  wire \dso[27]_i_7_n_0 ;
  wire \dso[27]_i_8_n_0 ;
  wire \dso[27]_i_9_n_0 ;
  wire \dso[31]_i_10_n_0 ;
  wire \dso[31]_i_11_n_0 ;
  wire \dso[31]_i_12_n_0 ;
  wire \dso[31]_i_13_n_0 ;
  wire \dso[31]_i_14_n_0 ;
  wire \dso[31]_i_15_n_0 ;
  wire \dso[31]_i_16_n_0 ;
  wire \dso[31]_i_3_n_0 ;
  wire \dso[31]_i_5_n_0 ;
  wire \dso[31]_i_6_n_0 ;
  wire \dso[31]_i_7_n_0 ;
  wire \dso[31]_i_8_n_0 ;
  wire \dso[31]_i_9_n_0 ;
  wire \dso[3]_i_10_n_0 ;
  wire \dso[3]_i_11_n_0 ;
  wire \dso[3]_i_12_n_0 ;
  wire \dso[3]_i_13_n_0 ;
  wire \dso[3]_i_2_n_0 ;
  wire \dso[3]_i_3_n_0 ;
  wire \dso[3]_i_4_n_0 ;
  wire \dso[3]_i_5_n_0 ;
  wire \dso[3]_i_6_n_0 ;
  wire \dso[3]_i_7_n_0 ;
  wire \dso[3]_i_8_n_0 ;
  wire \dso[3]_i_9_n_0 ;
  wire \dso[7]_i_10_n_0 ;
  wire \dso[7]_i_11_n_0 ;
  wire \dso[7]_i_12_n_0 ;
  wire \dso[7]_i_13_n_0 ;
  wire \dso[7]_i_2_n_0 ;
  wire \dso[7]_i_3_n_0 ;
  wire \dso[7]_i_4_n_0 ;
  wire \dso[7]_i_5_n_0 ;
  wire \dso[7]_i_6_n_0 ;
  wire \dso[7]_i_7_n_0 ;
  wire \dso[7]_i_8_n_0 ;
  wire \dso[7]_i_9_n_0 ;
  wire \dso_reg[11]_i_1_n_0 ;
  wire \dso_reg[11]_i_1_n_1 ;
  wire \dso_reg[11]_i_1_n_2 ;
  wire \dso_reg[11]_i_1_n_3 ;
  wire \dso_reg[15]_i_1_n_0 ;
  wire \dso_reg[15]_i_1_n_1 ;
  wire \dso_reg[15]_i_1_n_2 ;
  wire \dso_reg[15]_i_1_n_3 ;
  wire \dso_reg[19] ;
  wire \dso_reg[19]_0 ;
  wire \dso_reg[19]_1 ;
  wire \dso_reg[19]_2 ;
  wire \dso_reg[19]_i_1_n_0 ;
  wire \dso_reg[19]_i_1_n_1 ;
  wire \dso_reg[19]_i_1_n_2 ;
  wire \dso_reg[19]_i_1_n_3 ;
  wire \dso_reg[23] ;
  wire \dso_reg[23]_0 ;
  wire \dso_reg[23]_1 ;
  wire \dso_reg[23]_2 ;
  wire \dso_reg[23]_i_1_n_0 ;
  wire \dso_reg[23]_i_1_n_1 ;
  wire \dso_reg[23]_i_1_n_2 ;
  wire \dso_reg[23]_i_1_n_3 ;
  wire \dso_reg[27] ;
  wire \dso_reg[27]_0 ;
  wire \dso_reg[27]_1 ;
  wire \dso_reg[27]_2 ;
  wire \dso_reg[27]_i_1_n_0 ;
  wire \dso_reg[27]_i_1_n_1 ;
  wire \dso_reg[27]_i_1_n_2 ;
  wire \dso_reg[27]_i_1_n_3 ;
  wire [3:0]\dso_reg[31] ;
  wire \dso_reg[31]_0 ;
  wire \dso_reg[31]_1 ;
  wire \dso_reg[31]_2 ;
  wire \dso_reg[31]_3 ;
  wire \dso_reg[31]_i_2_n_1 ;
  wire \dso_reg[31]_i_2_n_2 ;
  wire \dso_reg[31]_i_2_n_3 ;
  wire \dso_reg[3]_i_1_n_0 ;
  wire \dso_reg[3]_i_1_n_1 ;
  wire \dso_reg[3]_i_1_n_2 ;
  wire \dso_reg[3]_i_1_n_3 ;
  wire \dso_reg[7]_i_1_n_0 ;
  wire \dso_reg[7]_i_1_n_1 ;
  wire \dso_reg[7]_i_1_n_2 ;
  wire \dso_reg[7]_i_1_n_3 ;
  wire [31:0]fdiv_rem;
  wire fdiv_rem_msb_f;
  wire [0:0]fdiv_rem_msb_f_reg_0;
  wire p_0_in;
  wire [31:0]p_0_out;
  wire \quo[31]_i_4_n_0 ;
  wire \quo[31]_i_5_n_0 ;
  wire \rem[11]_i_2_n_0 ;
  wire \rem[11]_i_3_n_0 ;
  wire \rem[11]_i_4_n_0 ;
  wire \rem[11]_i_5_n_0 ;
  wire \rem[11]_i_6_n_0 ;
  wire \rem[11]_i_7_n_0 ;
  wire \rem[11]_i_8_n_0 ;
  wire \rem[11]_i_9_n_0 ;
  wire \rem[15]_i_2_n_0 ;
  wire \rem[15]_i_3_n_0 ;
  wire \rem[15]_i_4_n_0 ;
  wire \rem[15]_i_5_n_0 ;
  wire \rem[15]_i_6_n_0 ;
  wire \rem[15]_i_7_n_0 ;
  wire \rem[15]_i_8_n_0 ;
  wire \rem[15]_i_9_n_0 ;
  wire \rem[19]_i_2_n_0 ;
  wire \rem[19]_i_3_n_0 ;
  wire \rem[19]_i_4_n_0 ;
  wire \rem[19]_i_5_n_0 ;
  wire \rem[19]_i_6_n_0 ;
  wire \rem[19]_i_7_n_0 ;
  wire \rem[19]_i_8_n_0 ;
  wire \rem[19]_i_9_n_0 ;
  wire \rem[23]_i_2_n_0 ;
  wire \rem[23]_i_3_n_0 ;
  wire \rem[23]_i_4_n_0 ;
  wire \rem[23]_i_5_n_0 ;
  wire \rem[23]_i_6_n_0 ;
  wire \rem[23]_i_7_n_0 ;
  wire \rem[23]_i_8_n_0 ;
  wire \rem[23]_i_9_n_0 ;
  wire \rem[27]_i_2_n_0 ;
  wire \rem[27]_i_3_n_0 ;
  wire \rem[27]_i_4_n_0 ;
  wire \rem[27]_i_5_n_0 ;
  wire \rem[27]_i_6_n_0 ;
  wire \rem[27]_i_7_n_0 ;
  wire \rem[27]_i_8_n_0 ;
  wire \rem[27]_i_9_n_0 ;
  wire \rem[31]_i_10_n_0 ;
  wire \rem[31]_i_11_n_0 ;
  wire \rem[31]_i_3_n_0 ;
  wire \rem[31]_i_4_n_0 ;
  wire \rem[31]_i_5_n_0 ;
  wire \rem[31]_i_6_n_0 ;
  wire \rem[31]_i_7_n_0 ;
  wire \rem[31]_i_8_n_0 ;
  wire \rem[31]_i_9_n_0 ;
  wire \rem[3]_i_2_n_0 ;
  wire \rem[3]_i_3_n_0 ;
  wire \rem[3]_i_4_n_0 ;
  wire \rem[3]_i_5_n_0 ;
  wire \rem[3]_i_6_n_0 ;
  wire \rem[3]_i_7_n_0 ;
  wire \rem[3]_i_8_n_0 ;
  wire \rem[3]_i_9_n_0 ;
  wire \rem[7]_i_2_n_0 ;
  wire \rem[7]_i_3_n_0 ;
  wire \rem[7]_i_4_n_0 ;
  wire \rem[7]_i_5_n_0 ;
  wire \rem[7]_i_6_n_0 ;
  wire \rem[7]_i_7_n_0 ;
  wire \rem[7]_i_8_n_0 ;
  wire \rem[7]_i_9_n_0 ;
  wire [3:0]\rem_reg[11] ;
  wire [3:0]\rem_reg[11]_0 ;
  wire \rem_reg[11]_i_1_n_0 ;
  wire \rem_reg[11]_i_1_n_1 ;
  wire \rem_reg[11]_i_1_n_2 ;
  wire \rem_reg[11]_i_1_n_3 ;
  wire [3:0]\rem_reg[15] ;
  wire [3:0]\rem_reg[15]_0 ;
  wire \rem_reg[15]_i_1_n_0 ;
  wire \rem_reg[15]_i_1_n_1 ;
  wire \rem_reg[15]_i_1_n_2 ;
  wire \rem_reg[15]_i_1_n_3 ;
  wire [3:0]\rem_reg[19] ;
  wire [3:0]\rem_reg[19]_0 ;
  wire \rem_reg[19]_i_1_n_0 ;
  wire \rem_reg[19]_i_1_n_1 ;
  wire \rem_reg[19]_i_1_n_2 ;
  wire \rem_reg[19]_i_1_n_3 ;
  wire [3:0]\rem_reg[23] ;
  wire [3:0]\rem_reg[23]_0 ;
  wire \rem_reg[23]_i_1_n_0 ;
  wire \rem_reg[23]_i_1_n_1 ;
  wire \rem_reg[23]_i_1_n_2 ;
  wire \rem_reg[23]_i_1_n_3 ;
  wire [3:0]\rem_reg[27] ;
  wire [3:0]\rem_reg[27]_0 ;
  wire \rem_reg[27]_i_1_n_0 ;
  wire \rem_reg[27]_i_1_n_1 ;
  wire \rem_reg[27]_i_1_n_2 ;
  wire \rem_reg[27]_i_1_n_3 ;
  wire [2:0]\rem_reg[30] ;
  wire [31:0]\rem_reg[31] ;
  wire [31:0]\rem_reg[31]_0 ;
  wire \rem_reg[31]_i_2_n_1 ;
  wire \rem_reg[31]_i_2_n_2 ;
  wire \rem_reg[31]_i_2_n_3 ;
  wire [3:0]\rem_reg[3] ;
  wire \rem_reg[3]_i_1_n_0 ;
  wire \rem_reg[3]_i_1_n_1 ;
  wire \rem_reg[3]_i_1_n_2 ;
  wire \rem_reg[3]_i_1_n_3 ;
  wire [3:0]\rem_reg[7] ;
  wire [3:0]\rem_reg[7]_0 ;
  wire \rem_reg[7]_i_1_n_0 ;
  wire \rem_reg[7]_i_1_n_1 ;
  wire \rem_reg[7]_i_1_n_2 ;
  wire \rem_reg[7]_i_1_n_3 ;
  wire \remden[64]_i_3_n_0 ;
  wire \remden[64]_i_4_n_0 ;
  wire \remden[64]_i_7_n_0 ;
  wire \remden_reg[0] ;
  wire \remden_reg[10] ;
  wire \remden_reg[11] ;
  wire \remden_reg[12] ;
  wire \remden_reg[13] ;
  wire \remden_reg[14] ;
  wire \remden_reg[15] ;
  wire \remden_reg[19] ;
  wire \remden_reg[28] ;
  wire \remden_reg[28]_0 ;
  wire \remden_reg[28]_1 ;
  wire \remden_reg[28]_2 ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire [20:0]\remden_reg[31] ;
  wire \remden_reg[31]_0 ;
  wire \remden_reg[31]_1 ;
  wire \remden_reg[4] ;
  wire \remden_reg[5] ;
  wire \remden_reg[64] ;
  wire \remden_reg[6] ;
  wire \remden_reg[7] ;
  wire \remden_reg[8] ;
  wire \remden_reg[9] ;
  wire rgf_sr_nh;
  wire rst_n;
  wire rst_n_0;
  wire rst_n_1;
  wire rst_n_10;
  wire rst_n_11;
  wire rst_n_12;
  wire rst_n_13;
  wire rst_n_14;
  wire rst_n_15;
  wire rst_n_16;
  wire rst_n_17;
  wire rst_n_18;
  wire rst_n_19;
  wire rst_n_2;
  wire rst_n_20;
  wire rst_n_21;
  wire rst_n_22;
  wire rst_n_23;
  wire rst_n_24;
  wire rst_n_25;
  wire rst_n_26;
  wire rst_n_27;
  wire rst_n_28;
  wire rst_n_29;
  wire rst_n_3;
  wire rst_n_30;
  wire rst_n_31;
  wire rst_n_32;
  wire rst_n_33;
  wire rst_n_34;
  wire rst_n_35;
  wire rst_n_36;
  wire rst_n_37;
  wire rst_n_4;
  wire rst_n_5;
  wire rst_n_6;
  wire rst_n_7;
  wire rst_n_8;
  wire rst_n_9;
  wire set_sgn;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire [31:0]\sr_reg[8]_11 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [7]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[7] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_14_n_0),
        .I3(\rem_reg[31]_0 [6]),
        .I4(add_out0_carry__6[6]),
        .O(p_0_out[6]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_15_n_0),
        .I3(\rem_reg[31]_0 [5]),
        .I4(add_out0_carry__6[5]),
        .O(p_0_out[5]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_16_n_0),
        .I3(\rem_reg[31]_0 [4]),
        .I4(add_out0_carry__6[4]),
        .O(p_0_out[4]));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__0_i_13
       (.I0(Q[7]),
        .I1(add_out0_carry__6[7]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\remden_reg[11] ),
        .O(add_out0_carry__0_i_13_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__0_i_14
       (.I0(\remden_reg[10] ),
        .I1(Q[6]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(add_out0_carry__6[6]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__0_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__0_i_15
       (.I0(add_out0_carry__6[5]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\dctl_stat_reg[2]_0 ),
        .I3(Q[5]),
        .I4(\remden_reg[9] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__0_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__0_i_16
       (.I0(Q[4]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[4]),
        .I4(\remden_reg[8] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__0_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [6]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[7] [2]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [5]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[7] [1]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__0_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [4]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[7] [0]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [7]),
        .I4(p_0_out[7]),
        .O(\rem_reg[7]_0 [3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [6]),
        .I4(p_0_out[6]),
        .O(\rem_reg[7]_0 [2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [5]),
        .I4(p_0_out[5]),
        .O(\rem_reg[7]_0 [1]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__0_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [4]),
        .I4(p_0_out[4]),
        .O(\rem_reg[7]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__0_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__0_i_13_n_0),
        .I3(\rem_reg[31]_0 [7]),
        .I4(add_out0_carry__6[7]),
        .O(p_0_out[7]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [11]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[11] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_14_n_0),
        .I3(\rem_reg[31]_0 [10]),
        .I4(add_out0_carry__6[10]),
        .O(p_0_out[10]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_15_n_0),
        .I3(\rem_reg[31]_0 [9]),
        .I4(add_out0_carry__6[9]),
        .O(p_0_out[9]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_16_n_0),
        .I3(\rem_reg[31]_0 [8]),
        .I4(add_out0_carry__6[8]),
        .O(p_0_out[8]));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__1_i_13
       (.I0(Q[11]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[11]),
        .I4(\remden_reg[15] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__1_i_13_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__1_i_14
       (.I0(Q[10]),
        .I1(add_out0_carry__6[10]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\remden_reg[14] ),
        .O(add_out0_carry__1_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__1_i_15
       (.I0(add_out0_carry__6[9]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\dctl_stat_reg[2]_0 ),
        .I3(Q[9]),
        .I4(\remden_reg[13] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__1_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__1_i_16
       (.I0(Q[8]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[8]),
        .I4(\remden_reg[12] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__1_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [10]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[11] [2]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [9]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[11] [1]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__1_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [8]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[11] [0]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [11]),
        .I4(p_0_out[11]),
        .O(\rem_reg[11]_0 [3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [10]),
        .I4(p_0_out[10]),
        .O(\rem_reg[11]_0 [2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [9]),
        .I4(p_0_out[9]),
        .O(\rem_reg[11]_0 [1]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__1_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [8]),
        .I4(p_0_out[8]),
        .O(\rem_reg[11]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__1_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__1_i_13_n_0),
        .I3(\rem_reg[31]_0 [11]),
        .I4(add_out0_carry__6[11]),
        .O(p_0_out[11]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [15]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[15] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_14_n_0),
        .I3(\rem_reg[31]_0 [14]),
        .I4(add_out0_carry__6[14]),
        .O(p_0_out[14]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_15_n_0),
        .I3(\rem_reg[31]_0 [13]),
        .I4(add_out0_carry__6[13]),
        .O(p_0_out[13]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_16_n_0),
        .I3(\rem_reg[31]_0 [12]),
        .I4(add_out0_carry__6[12]),
        .O(p_0_out[12]));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__2_i_13
       (.I0(Q[15]),
        .I1(add_out0_carry__6[15]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(add_out0_carry__2_i_9_0),
        .O(add_out0_carry__2_i_13_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__2_i_14
       (.I0(Q[14]),
        .I1(add_out0_carry__6[14]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(add_out0_carry__2_i_10_0),
        .O(add_out0_carry__2_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__2_i_15
       (.I0(Q[13]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[13]),
        .I4(add_out0_carry__2_i_11_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__2_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__2_i_16
       (.I0(Q[12]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[12]),
        .I4(add_out0_carry__2_i_12_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__2_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [14]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[15] [2]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [13]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[15] [1]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__2_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [12]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[15] [0]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [15]),
        .I4(p_0_out[15]),
        .O(\rem_reg[15]_0 [3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [14]),
        .I4(p_0_out[14]),
        .O(\rem_reg[15]_0 [2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [13]),
        .I4(p_0_out[13]),
        .O(\rem_reg[15]_0 [1]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__2_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [12]),
        .I4(p_0_out[12]),
        .O(\rem_reg[15]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__2_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__2_i_13_n_0),
        .I3(\rem_reg[31]_0 [15]),
        .I4(add_out0_carry__6[15]),
        .O(p_0_out[15]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [19]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[19] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_14_n_0),
        .I3(\rem_reg[31]_0 [18]),
        .I4(add_out0_carry__6[18]),
        .O(p_0_out[18]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_15_n_0),
        .I3(\rem_reg[31]_0 [17]),
        .I4(add_out0_carry__6[17]),
        .O(p_0_out[17]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_16_n_0),
        .I3(\rem_reg[31]_0 [16]),
        .I4(add_out0_carry__6[16]),
        .O(p_0_out[16]));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__3_i_13
       (.I0(add_out0_carry__3_i_9_0),
        .I1(Q[19]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(add_out0_carry__6[19]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__3_i_13_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__3_i_14
       (.I0(Q[18]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[18]),
        .I4(add_out0_carry__3_i_10_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__3_i_14_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__3_i_15
       (.I0(Q[17]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[17]),
        .I4(add_out0_carry__3_i_11_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__3_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__3_i_16
       (.I0(Q[16]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[16]),
        .I4(add_out0_carry__3_i_12_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__3_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [18]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[19] [2]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [17]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[19] [1]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__3_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [16]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[19] [0]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [19]),
        .I4(p_0_out[19]),
        .O(\rem_reg[19]_0 [3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [18]),
        .I4(p_0_out[18]),
        .O(\rem_reg[19]_0 [2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [17]),
        .I4(p_0_out[17]),
        .O(\rem_reg[19]_0 [1]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__3_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [16]),
        .I4(p_0_out[16]),
        .O(\rem_reg[19]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__3_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__3_i_13_n_0),
        .I3(\rem_reg[31]_0 [19]),
        .I4(add_out0_carry__6[19]),
        .O(p_0_out[19]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [23]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[23] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_14_n_0),
        .I3(\rem_reg[31]_0 [22]),
        .I4(add_out0_carry__6[22]),
        .O(p_0_out[22]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_15_n_0),
        .I3(\rem_reg[31]_0 [21]),
        .I4(add_out0_carry__6[21]),
        .O(p_0_out[21]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_16_n_0),
        .I3(\rem_reg[31]_0 [20]),
        .I4(add_out0_carry__6[20]),
        .O(p_0_out[20]));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__4_i_13
       (.I0(Q[23]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[23]),
        .I4(add_out0_carry__4_i_9_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__4_i_13_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__4_i_14
       (.I0(add_out0_carry__4_i_10_0),
        .I1(Q[22]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(add_out0_carry__6[22]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_14_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__4_i_15
       (.I0(Q[21]),
        .I1(add_out0_carry__6[21]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(add_out0_carry__4_i_11_0),
        .O(add_out0_carry__4_i_15_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__4_i_16
       (.I0(add_out0_carry__4_i_12_0),
        .I1(Q[20]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(add_out0_carry__6[20]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__4_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [22]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[23] [2]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [21]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[23] [1]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__4_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [20]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[23] [0]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [23]),
        .I4(p_0_out[23]),
        .O(\rem_reg[23]_0 [3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [22]),
        .I4(p_0_out[22]),
        .O(\rem_reg[23]_0 [2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [21]),
        .I4(p_0_out[21]),
        .O(\rem_reg[23]_0 [1]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__4_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [20]),
        .I4(p_0_out[20]),
        .O(\rem_reg[23]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__4_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__4_i_13_n_0),
        .I3(\rem_reg[31]_0 [23]),
        .I4(add_out0_carry__6[23]),
        .O(p_0_out[23]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [27]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[27] [3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_14_n_0),
        .I3(\rem_reg[31]_0 [26]),
        .I4(add_out0_carry__6[26]),
        .O(p_0_out[26]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_15_n_0),
        .I3(\rem_reg[31]_0 [25]),
        .I4(add_out0_carry__6[25]),
        .O(p_0_out[25]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_16_n_0),
        .I3(\rem_reg[31]_0 [24]),
        .I4(add_out0_carry__6[24]),
        .O(p_0_out[24]));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__5_i_13
       (.I0(Q[27]),
        .I1(add_out0_carry__6[27]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\remden_reg[31]_0 ),
        .O(add_out0_carry__5_i_13_n_0));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__5_i_14
       (.I0(add_out0_carry__5_i_10_0),
        .I1(Q[26]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(add_out0_carry__6[26]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__5_i_14_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__5_i_15
       (.I0(Q[25]),
        .I1(add_out0_carry__6[25]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(add_out0_carry__5_i_11_0),
        .O(add_out0_carry__5_i_15_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__5_i_16
       (.I0(Q[24]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[24]),
        .I4(add_out0_carry__5_i_12_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__5_i_16_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [26]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[27] [2]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [25]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[27] [1]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__5_i_4
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [24]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[27] [0]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [27]),
        .I4(p_0_out[27]),
        .O(\rem_reg[27]_0 [3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [26]),
        .I4(p_0_out[26]),
        .O(\rem_reg[27]_0 [2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [25]),
        .I4(p_0_out[25]),
        .O(\rem_reg[27]_0 [1]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__5_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [24]),
        .I4(p_0_out[24]),
        .O(\rem_reg[27]_0 [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__5_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__5_i_13_n_0),
        .I3(\rem_reg[31]_0 [27]),
        .I4(add_out0_carry__6[27]),
        .O(p_0_out[27]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__6_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [30]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[30] [2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_10
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__6_i_13_n_0),
        .I3(\rem_reg[31]_0 [28]),
        .I4(add_out0_carry__6[28]),
        .O(p_0_out[28]));
  LUT5 #(
    .INIT(32'h303F5050)) 
    add_out0_carry__6_i_11
       (.I0(DI),
        .I1(Q[30]),
        .I2(add_out0_carry_i_9_n_0),
        .I3(add_out0_carry__6[30]),
        .I4(add_out0_carry_i_10_n_0),
        .O(add_out0_carry__6_i_11_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry__6_i_12
       (.I0(Q[29]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[29]),
        .I4(add_out0_carry__6_i_9_0),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry__6_i_12_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry__6_i_13
       (.I0(Q[28]),
        .I1(add_out0_carry__6[28]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(add_out0_carry__6_i_10_0),
        .O(add_out0_carry__6_i_13_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__6_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [29]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[30] [1]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry__6_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [28]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[30] [0]));
  LUT6 #(
    .INIT(64'h30305050B5BA50FF)) 
    add_out0_carry__6_i_4
       (.I0(add_out0_carry__6[31]),
        .I1(Q[31]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [31]),
        .I4(add_out0_carry_i_9_n_0),
        .I5(\rem[31]_i_3_n_0 ),
        .O(\dso_reg[31] [3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__6_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [30]),
        .I4(p_0_out[30]),
        .O(\dso_reg[31] [2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__6_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [29]),
        .I4(p_0_out[29]),
        .O(\dso_reg[31] [1]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry__6_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [28]),
        .I4(p_0_out[28]),
        .O(\dso_reg[31] [0]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_8
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__6_i_11_n_0),
        .I3(\rem_reg[31]_0 [30]),
        .I4(add_out0_carry__6[30]),
        .O(p_0_out[30]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry__6_i_9
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry__6_i_12_n_0),
        .I3(\rem_reg[31]_0 [29]),
        .I4(add_out0_carry__6[29]),
        .O(p_0_out[29]));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry_i_1
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [3]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[3] [3]));
  LUT6 #(
    .INIT(64'h04FF000004000000)) 
    add_out0_carry_i_10
       (.I0(dctl_stat[2]),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[1]),
        .I4(dctl_stat[3]),
        .I5(add_out0_carry_i_16_n_0),
        .O(add_out0_carry_i_10_n_0));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_11
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_17_n_0),
        .I3(\rem_reg[31]_0 [3]),
        .I4(add_out0_carry__6[3]),
        .O(p_0_out[3]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_12
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_18_n_0),
        .I3(\rem_reg[31]_0 [2]),
        .I4(add_out0_carry__6[2]),
        .O(p_0_out[2]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_13
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_19_n_0),
        .I3(\rem_reg[31]_0 [1]),
        .I4(add_out0_carry__6[1]),
        .O(p_0_out[1]));
  LUT5 #(
    .INIT(32'hE4F5A0B1)) 
    add_out0_carry_i_14
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(add_out0_carry_i_9_n_0),
        .I2(add_out0_carry_i_20_n_0),
        .I3(\rem_reg[31]_0 [0]),
        .I4(add_out0_carry__6[0]),
        .O(p_0_out[0]));
  LUT6 #(
    .INIT(64'hF0FF7070F0FF707F)) 
    add_out0_carry_i_15
       (.I0(dctl_sign),
        .I1(den2),
        .I2(dctl_stat[0]),
        .I3(chg_quo_sgn),
        .I4(dctl_stat[1]),
        .I5(fdiv_rem_msb_f),
        .O(add_out0_carry_i_15_n_0));
  LUT6 #(
    .INIT(64'h0000F0002200F0FF)) 
    add_out0_carry_i_16
       (.I0(dctl_sign),
        .I1(den2),
        .I2(add_out0_carry_i_21_n_0),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[0]),
        .I5(chg_quo_sgn_reg_0),
        .O(add_out0_carry_i_16_n_0));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry_i_17
       (.I0(add_out0_carry__6[3]),
        .I1(\dso[31]_i_3_n_0 ),
        .I2(\dctl_stat_reg[2]_0 ),
        .I3(Q[3]),
        .I4(\remden_reg[7] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry_i_17_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry_i_18
       (.I0(Q[2]),
        .I1(add_out0_carry__6[2]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\remden_reg[6] ),
        .O(add_out0_carry_i_18_n_0));
  LUT5 #(
    .INIT(32'h50305F30)) 
    add_out0_carry_i_19
       (.I0(Q[1]),
        .I1(add_out0_carry__6[1]),
        .I2(add_out0_carry_i_10_n_0),
        .I3(add_out0_carry_i_9_n_0),
        .I4(\remden_reg[5] ),
        .O(add_out0_carry_i_19_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry_i_2
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [2]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[3] [2]));
  LUT6 #(
    .INIT(64'h44F444F444F4FFFF)) 
    add_out0_carry_i_20
       (.I0(Q[0]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(\dso[31]_i_3_n_0 ),
        .I3(add_out0_carry__6[0]),
        .I4(\remden_reg[4] ),
        .I5(\remden[64]_i_7_n_0 ),
        .O(add_out0_carry_i_20_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    add_out0_carry_i_21
       (.I0(chg_quo_sgn),
        .I1(fdiv_rem_msb_f),
        .O(add_out0_carry_i_21_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    add_out0_carry_i_3
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [1]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\rem_reg[3] [1]));
  LUT4 #(
    .INIT(16'hFCBB)) 
    add_out0_carry_i_4
       (.I0(add_out0_carry_i_10_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [0]),
        .I3(add_out0_carry_i_9_n_0),
        .O(\rem_reg[3] [0]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry_i_5
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [3]),
        .I4(p_0_out[3]),
        .O(S[3]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry_i_6
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [2]),
        .I4(p_0_out[2]),
        .O(S[2]));
  LUT5 #(
    .INIT(32'hFDFF0200)) 
    add_out0_carry_i_7
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(add_out0_carry_i_10_n_0),
        .I3(\rem_reg[31]_0 [1]),
        .I4(p_0_out[1]),
        .O(S[1]));
  LUT5 #(
    .INIT(32'h0252FDAD)) 
    add_out0_carry_i_8
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem_reg[31]_0 [0]),
        .I2(\rem[31]_i_3_n_0 ),
        .I3(add_out0_carry_i_10_n_0),
        .I4(p_0_out[0]),
        .O(S[0]));
  LUT4 #(
    .INIT(16'h0028)) 
    add_out0_carry_i_9
       (.I0(dctl_stat[3]),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[1]),
        .I3(add_out0_carry_i_15_n_0),
        .O(add_out0_carry_i_9_n_0));
  LUT5 #(
    .INIT(32'h82FF8200)) 
    chg_quo_sgn_i_1
       (.I0(dctl_sign),
        .I1(chg_quo_sgn_reg_0),
        .I2(den2),
        .I3(set_sgn),
        .I4(chg_quo_sgn),
        .O(chg_quo_sgn_i_1_n_0));
  FDRE chg_quo_sgn_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_quo_sgn_i_1_n_0),
        .Q(chg_quo_sgn),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'hEFFFFFFF20000000)) 
    chg_rem_sgn_i_1
       (.I0(chg_rem_sgn0),
        .I1(dctl_stat[1]),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[3]),
        .I5(chg_rem_sgn),
        .O(chg_rem_sgn_i_1_n_0));
  FDRE chg_rem_sgn_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(chg_rem_sgn_i_1_n_0),
        .Q(chg_rem_sgn),
        .R(p_0_in));
  LUT3 #(
    .INIT(8'hB8)) 
    dctl_long_f_i_1
       (.I0(rgf_sr_nh),
        .I1(dctl_long_f_reg_0),
        .I2(dctl_long_f_reg),
        .O(dctl_long));
  LUT6 #(
    .INIT(64'h4F4F5F5F404F5050)) 
    \dctl_stat[0]_i_1 
       (.I0(dctl_stat[0]),
        .I1(\dctl_stat[1]_i_3_n_0 ),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .I5(\dctl_stat[0]_i_2_n_0 ),
        .O(dctl_next[0]));
  LUT6 #(
    .INIT(64'h007F007F0000007F)) 
    \dctl_stat[0]_i_2 
       (.I0(den2),
        .I1(dctl_sign),
        .I2(dctl_stat[0]),
        .I3(\dctl_stat[0]_i_3_n_0 ),
        .I4(\dctl_stat_reg[2]_2 ),
        .I5(dctl_stat[2]),
        .O(\dctl_stat[0]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00FFD700)) 
    \dctl_stat[0]_i_3 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .I2(fdiv_rem_msb_f),
        .I3(dctl_stat[3]),
        .I4(dctl_stat[0]),
        .O(\dctl_stat[0]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0F300B38)) 
    \dctl_stat[1]_i_1 
       (.I0(\dctl_stat[1]_i_2_n_0 ),
        .I1(dctl_stat[3]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[1]),
        .I4(\dctl_stat[1]_i_3_n_0 ),
        .O(dctl_next[1]));
  LUT5 #(
    .INIT(32'h0C080800)) 
    \dctl_stat[1]_i_2 
       (.I0(fdiv_rem_msb_f),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[1]),
        .I3(chg_quo_sgn),
        .I4(chg_rem_sgn),
        .O(\dctl_stat[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \dctl_stat[1]_i_3 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[2]),
        .O(\dctl_stat[1]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0000FFC1)) 
    \dctl_stat[2]_i_1 
       (.I0(\dctl_stat_reg[2]_2 ),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .O(dctl_next[2]));
  LUT6 #(
    .INIT(64'hF4F4F4F4F4FFF4F4)) 
    \dctl_stat[3]_i_1 
       (.I0(\dctl_stat_reg[3]_1 ),
        .I1(set_sgn),
        .I2(\dctl_stat[3]_i_4_n_0 ),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[3]),
        .I5(\dctl_stat[3]_i_5_n_0 ),
        .O(dctl_next[3]));
  LUT4 #(
    .INIT(16'h4000)) 
    \dctl_stat[3]_i_3 
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[3]),
        .O(set_sgn));
  LUT6 #(
    .INIT(64'h00000000F5000003)) 
    \dctl_stat[3]_i_4 
       (.I0(dctl_long),
        .I1(\dctl_stat_reg[2]_2 ),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[1]),
        .I4(dctl_stat[0]),
        .I5(dctl_stat[3]),
        .O(\dctl_stat[3]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF00AFF3AFF3AFFFA)) 
    \dctl_stat[3]_i_5 
       (.I0(chg_quo_sgn_reg_0),
        .I1(fdiv_rem_msb_f),
        .I2(dctl_stat[2]),
        .I3(dctl_stat[1]),
        .I4(chg_quo_sgn),
        .I5(chg_rem_sgn),
        .O(\dctl_stat[3]_i_5_n_0 ));
  FDRE \dctl_stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[0]),
        .Q(dctl_stat[0]),
        .R(p_0_in));
  FDRE \dctl_stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[1]),
        .Q(dctl_stat[1]),
        .R(p_0_in));
  FDRE \dctl_stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[2]),
        .Q(dctl_stat[2]),
        .R(p_0_in));
  FDRE \dctl_stat_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(dctl_next[3]),
        .Q(dctl_stat[3]),
        .R(p_0_in));
  LUT3 #(
    .INIT(8'hC8)) 
    div_crdy_i_1
       (.I0(div_crdy_i_2_n_0),
        .I1(\dctl_stat_reg[2]_2 ),
        .I2(dctl_long_f_reg_0),
        .O(div_crdy_reg_0));
  LUT5 #(
    .INIT(32'hFFFF5700)) 
    div_crdy_i_2
       (.I0(dctl_sign),
        .I1(chg_rem_sgn),
        .I2(chg_quo_sgn),
        .I3(div_crdy_i_3_n_0),
        .I4(div_crdy_i_4_n_0),
        .O(div_crdy_i_2_n_0));
  LUT5 #(
    .INIT(32'h08000808)) 
    div_crdy_i_3
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[2]),
        .I4(dctl_long),
        .O(div_crdy_i_3_n_0));
  LUT6 #(
    .INIT(64'h000000F000700000)) 
    div_crdy_i_4
       (.I0(fdiv_rem_msb_f),
        .I1(chg_quo_sgn),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[2]),
        .I5(dctl_stat[1]),
        .O(div_crdy_i_4_n_0));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [11]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [10]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [9]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[11]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [8]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[11]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_2 
       (.I0(p_0_out[11]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_3 
       (.I0(p_0_out[10]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_4 
       (.I0(p_0_out[9]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[11]_i_5 
       (.I0(p_0_out[8]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_6 
       (.I0(p_0_out[11]),
        .I1(\dso[11]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [11]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[11]),
        .O(\dso[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_7 
       (.I0(p_0_out[10]),
        .I1(\dso[11]_i_11_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [10]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[10]),
        .O(\dso[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_8 
       (.I0(p_0_out[9]),
        .I1(\dso[11]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [9]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[9]),
        .O(\dso[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[11]_i_9 
       (.I0(p_0_out[8]),
        .I1(\dso[11]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [8]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[8]),
        .O(\dso[11]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [15]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hE2FF)) 
    \dso[15]_i_11 
       (.I0(dctl_long_f_reg),
        .I1(dctl_long_f_reg_0),
        .I2(rgf_sr_nh),
        .I3(\dso[31]_i_3_n_0 ),
        .O(\dso[15]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [14]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [13]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[15]_i_14 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [12]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[15]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_2 
       (.I0(p_0_out[15]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_3 
       (.I0(p_0_out[14]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_4 
       (.I0(p_0_out[13]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[15]_i_5 
       (.I0(p_0_out[12]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_6 
       (.I0(p_0_out[15]),
        .I1(\dso[15]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [15]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[15]),
        .O(\dso[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_7 
       (.I0(p_0_out[14]),
        .I1(\dso[15]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [14]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[14]),
        .O(\dso[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_8 
       (.I0(p_0_out[13]),
        .I1(\dso[15]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [13]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[13]),
        .O(\dso[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[15]_i_9 
       (.I0(p_0_out[12]),
        .I1(\dso[15]_i_14_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [12]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[12]),
        .O(\dso[15]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [19]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [18]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [17]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[19]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [16]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[19]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_2 
       (.I0(p_0_out[19]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_3 
       (.I0(p_0_out[18]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_4 
       (.I0(p_0_out[17]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[19]_i_5 
       (.I0(p_0_out[16]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_6 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[19]),
        .I3(\dso[19]_i_10_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[19]_2 ),
        .O(\dso[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_7 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[18]),
        .I3(\dso[19]_i_11_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[19]_1 ),
        .O(\dso[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_8 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[17]),
        .I3(\dso[19]_i_12_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[19]_0 ),
        .O(\dso[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[19]_i_9 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[16]),
        .I3(\dso[19]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[19] ),
        .O(\dso[19]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [23]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [22]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [21]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[23]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [20]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[23]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_2 
       (.I0(p_0_out[23]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_3 
       (.I0(p_0_out[22]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_4 
       (.I0(p_0_out[21]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[23]_i_5 
       (.I0(p_0_out[20]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_6 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[23]),
        .I3(\dso[23]_i_10_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[23]_2 ),
        .O(\dso[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_7 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[22]),
        .I3(\dso[23]_i_11_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[23]_1 ),
        .O(\dso[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_8 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[21]),
        .I3(\dso[23]_i_12_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[23]_0 ),
        .O(\dso[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[23]_i_9 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[20]),
        .I3(\dso[23]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[23] ),
        .O(\dso[23]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [27]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [26]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [25]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[27]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [24]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[27]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_2 
       (.I0(p_0_out[27]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_3 
       (.I0(p_0_out[26]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_4 
       (.I0(p_0_out[25]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[27]_i_5 
       (.I0(p_0_out[24]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_6 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[27]),
        .I3(\dso[27]_i_10_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[27]_2 ),
        .O(\dso[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_7 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[26]),
        .I3(\dso[27]_i_11_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[27]_1 ),
        .O(\dso[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_8 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[25]),
        .I3(\dso[27]_i_12_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[27]_0 ),
        .O(\dso[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[27]_i_9 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[24]),
        .I3(\dso[27]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[27] ),
        .O(\dso[27]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \dso[31]_i_1 
       (.I0(\dso[31]_i_3_n_0 ),
        .I1(\remden_reg[0] ),
        .O(div_crdy_reg));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_10 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[29]),
        .I3(\dso[31]_i_15_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[31]_1 ),
        .O(\dso[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_11 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[28]),
        .I3(\dso[31]_i_16_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[31]_0 ),
        .O(\dso[31]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h1DFF)) 
    \dso[31]_i_12 
       (.I0(dctl_long_f_reg),
        .I1(dctl_long_f_reg_0),
        .I2(rgf_sr_nh),
        .I3(\dso[31]_i_3_n_0 ),
        .O(\dso[31]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [31]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_14 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [30]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_15 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [29]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[31]_i_16 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [28]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[31]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_3 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(add_out0_carry_i_9_n_0),
        .O(\dso[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_5 
       (.I0(p_0_out[30]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_6 
       (.I0(p_0_out[29]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[31]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[31]_i_7 
       (.I0(p_0_out[28]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_8 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[31]),
        .I3(\dso[31]_i_13_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[31]_3 ),
        .O(\dso[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000FF088880FF0)) 
    \dso[31]_i_9 
       (.I0(\remden_reg[0] ),
        .I1(rgf_sr_nh),
        .I2(p_0_out[30]),
        .I3(\dso[31]_i_14_n_0 ),
        .I4(\dso[31]_i_12_n_0 ),
        .I5(\dso_reg[31]_2 ),
        .O(\dso[31]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[3]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [3]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[3]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[3]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [2]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[3]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[3]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [1]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[3]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'hFCBB)) 
    \dso[3]_i_13 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [0]),
        .I3(add_out0_carry_i_9_n_0),
        .O(\dso[3]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_2 
       (.I0(p_0_out[3]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_3 
       (.I0(p_0_out[2]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_4 
       (.I0(p_0_out[1]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[3]_i_5 
       (.I0(p_0_out[0]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_6 
       (.I0(p_0_out[3]),
        .I1(\dso[3]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [3]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[3]),
        .O(\dso[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_7 
       (.I0(p_0_out[2]),
        .I1(\dso[3]_i_11_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [2]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[2]),
        .O(\dso[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_8 
       (.I0(p_0_out[1]),
        .I1(\dso[3]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [1]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[1]),
        .O(\dso[3]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[3]_i_9 
       (.I0(p_0_out[0]),
        .I1(\dso[3]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [0]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[0]),
        .O(\dso[3]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [7]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_11 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [6]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_12 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [5]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_12_n_0 ));
  LUT4 #(
    .INIT(16'h0020)) 
    \dso[7]_i_13 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(\rem_reg[31]_0 [4]),
        .I3(add_out0_carry_i_10_n_0),
        .O(\dso[7]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_2 
       (.I0(p_0_out[7]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_3 
       (.I0(p_0_out[6]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_4 
       (.I0(p_0_out[5]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \dso[7]_i_5 
       (.I0(p_0_out[4]),
        .I1(\dso[31]_i_12_n_0 ),
        .O(\dso[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_6 
       (.I0(p_0_out[7]),
        .I1(\dso[7]_i_10_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [7]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[7]),
        .O(\dso[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_7 
       (.I0(p_0_out[6]),
        .I1(\dso[7]_i_11_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [6]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[6]),
        .O(\dso[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_8 
       (.I0(p_0_out[5]),
        .I1(\dso[7]_i_12_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [5]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[5]),
        .O(\dso[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hF6F6F6060606F606)) 
    \dso[7]_i_9 
       (.I0(p_0_out[4]),
        .I1(\dso[7]_i_13_n_0 ),
        .I2(\dso[31]_i_12_n_0 ),
        .I3(\remden_reg[31] [4]),
        .I4(\dso[15]_i_11_n_0 ),
        .I5(bbus_0[4]),
        .O(\dso[7]_i_9_n_0 ));
  CARRY4 \dso_reg[11]_i_1 
       (.CI(\dso_reg[7]_i_1_n_0 ),
        .CO({\dso_reg[11]_i_1_n_0 ,\dso_reg[11]_i_1_n_1 ,\dso_reg[11]_i_1_n_2 ,\dso_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[11]_i_2_n_0 ,\dso[11]_i_3_n_0 ,\dso[11]_i_4_n_0 ,\dso[11]_i_5_n_0 }),
        .O(\sr_reg[8]_11 [11:8]),
        .S({\dso[11]_i_6_n_0 ,\dso[11]_i_7_n_0 ,\dso[11]_i_8_n_0 ,\dso[11]_i_9_n_0 }));
  CARRY4 \dso_reg[15]_i_1 
       (.CI(\dso_reg[11]_i_1_n_0 ),
        .CO({\dso_reg[15]_i_1_n_0 ,\dso_reg[15]_i_1_n_1 ,\dso_reg[15]_i_1_n_2 ,\dso_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[15]_i_2_n_0 ,\dso[15]_i_3_n_0 ,\dso[15]_i_4_n_0 ,\dso[15]_i_5_n_0 }),
        .O(\sr_reg[8]_11 [15:12]),
        .S({\dso[15]_i_6_n_0 ,\dso[15]_i_7_n_0 ,\dso[15]_i_8_n_0 ,\dso[15]_i_9_n_0 }));
  CARRY4 \dso_reg[19]_i_1 
       (.CI(\dso_reg[15]_i_1_n_0 ),
        .CO({\dso_reg[19]_i_1_n_0 ,\dso_reg[19]_i_1_n_1 ,\dso_reg[19]_i_1_n_2 ,\dso_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[19]_i_2_n_0 ,\dso[19]_i_3_n_0 ,\dso[19]_i_4_n_0 ,\dso[19]_i_5_n_0 }),
        .O(\sr_reg[8]_11 [19:16]),
        .S({\dso[19]_i_6_n_0 ,\dso[19]_i_7_n_0 ,\dso[19]_i_8_n_0 ,\dso[19]_i_9_n_0 }));
  CARRY4 \dso_reg[23]_i_1 
       (.CI(\dso_reg[19]_i_1_n_0 ),
        .CO({\dso_reg[23]_i_1_n_0 ,\dso_reg[23]_i_1_n_1 ,\dso_reg[23]_i_1_n_2 ,\dso_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[23]_i_2_n_0 ,\dso[23]_i_3_n_0 ,\dso[23]_i_4_n_0 ,\dso[23]_i_5_n_0 }),
        .O(\sr_reg[8]_11 [23:20]),
        .S({\dso[23]_i_6_n_0 ,\dso[23]_i_7_n_0 ,\dso[23]_i_8_n_0 ,\dso[23]_i_9_n_0 }));
  CARRY4 \dso_reg[27]_i_1 
       (.CI(\dso_reg[23]_i_1_n_0 ),
        .CO({\dso_reg[27]_i_1_n_0 ,\dso_reg[27]_i_1_n_1 ,\dso_reg[27]_i_1_n_2 ,\dso_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[27]_i_2_n_0 ,\dso[27]_i_3_n_0 ,\dso[27]_i_4_n_0 ,\dso[27]_i_5_n_0 }),
        .O(\sr_reg[8]_11 [27:24]),
        .S({\dso[27]_i_6_n_0 ,\dso[27]_i_7_n_0 ,\dso[27]_i_8_n_0 ,\dso[27]_i_9_n_0 }));
  CARRY4 \dso_reg[31]_i_2 
       (.CI(\dso_reg[27]_i_1_n_0 ),
        .CO({\dso_reg[31]_i_2_n_1 ,\dso_reg[31]_i_2_n_2 ,\dso_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\dso[31]_i_5_n_0 ,\dso[31]_i_6_n_0 ,\dso[31]_i_7_n_0 }),
        .O(\sr_reg[8]_11 [31:28]),
        .S({\dso[31]_i_8_n_0 ,\dso[31]_i_9_n_0 ,\dso[31]_i_10_n_0 ,\dso[31]_i_11_n_0 }));
  CARRY4 \dso_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\dso_reg[3]_i_1_n_0 ,\dso_reg[3]_i_1_n_1 ,\dso_reg[3]_i_1_n_2 ,\dso_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[3]_i_2_n_0 ,\dso[3]_i_3_n_0 ,\dso[3]_i_4_n_0 ,\dso[3]_i_5_n_0 }),
        .O(\sr_reg[8]_11 [3:0]),
        .S({\dso[3]_i_6_n_0 ,\dso[3]_i_7_n_0 ,\dso[3]_i_8_n_0 ,\dso[3]_i_9_n_0 }));
  CARRY4 \dso_reg[7]_i_1 
       (.CI(\dso_reg[3]_i_1_n_0 ),
        .CO({\dso_reg[7]_i_1_n_0 ,\dso_reg[7]_i_1_n_1 ,\dso_reg[7]_i_1_n_2 ,\dso_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\dso[7]_i_2_n_0 ,\dso[7]_i_3_n_0 ,\dso[7]_i_4_n_0 ,\dso[7]_i_5_n_0 }),
        .O(\sr_reg[8]_11 [7:4]),
        .S({\dso[7]_i_6_n_0 ,\dso[7]_i_7_n_0 ,\dso[7]_i_8_n_0 ,\dso[7]_i_9_n_0 }));
  FDRE fdiv_rem_msb_f_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fdiv_rem_msb_f_reg_0),
        .Q(fdiv_rem_msb_f),
        .R(p_0_in));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[28]_i_1 
       (.I0(\remden_reg[31] [17]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(Q[24]),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[29]_i_1 
       (.I0(\remden_reg[31] [18]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(Q[25]),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[30]_i_1 
       (.I0(\remden_reg[31] [19]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(Q[26]),
        .O(D[2]));
  LUT6 #(
    .INIT(64'hEFEFEFEFEFEFEFEE)) 
    \quo[31]_i_1 
       (.I0(\dctl_stat_reg[2]_0 ),
        .I1(\quo[31]_i_4_n_0 ),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[1]),
        .I5(dctl_stat[0]),
        .O(E));
  LUT3 #(
    .INIT(8'hB8)) 
    \quo[31]_i_2 
       (.I0(\remden_reg[31] [20]),
        .I1(\dctl_stat_reg[2]_0 ),
        .I2(Q[27]),
        .O(D[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \quo[31]_i_3 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(add_out0_carry_i_9_n_0),
        .O(\dctl_stat_reg[2]_0 ));
  LUT6 #(
    .INIT(64'h0022202232323232)) 
    \quo[31]_i_4 
       (.I0(dctl_stat[0]),
        .I1(\quo[31]_i_5_n_0 ),
        .I2(chg_quo_sgn_reg_0),
        .I3(dctl_sign),
        .I4(den2),
        .I5(dctl_stat[2]),
        .O(\quo[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \quo[31]_i_5 
       (.I0(dctl_stat[1]),
        .I1(dctl_stat[3]),
        .O(\quo[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_2 
       (.I0(p_0_out[11]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_3 
       (.I0(p_0_out[10]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_4 
       (.I0(p_0_out[9]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[11]_i_5 
       (.I0(p_0_out[8]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[11]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[11]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [11]),
        .I5(fdiv_rem[11]),
        .O(\rem[11]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[10]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [10]),
        .I5(fdiv_rem[10]),
        .O(\rem[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[9]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [9]),
        .I5(fdiv_rem[9]),
        .O(\rem[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[11]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[8]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [8]),
        .I5(fdiv_rem[8]),
        .O(\rem[11]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_2 
       (.I0(p_0_out[15]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_3 
       (.I0(p_0_out[14]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_4 
       (.I0(p_0_out[13]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[15]_i_5 
       (.I0(p_0_out[12]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[15]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[15]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [15]),
        .I5(fdiv_rem[15]),
        .O(\rem[15]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[14]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [14]),
        .I5(fdiv_rem[14]),
        .O(\rem[15]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[13]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [13]),
        .I5(fdiv_rem[13]),
        .O(\rem[15]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[15]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[12]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [12]),
        .I5(fdiv_rem[12]),
        .O(\rem[15]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_2 
       (.I0(p_0_out[19]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_3 
       (.I0(p_0_out[18]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_4 
       (.I0(p_0_out[17]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[19]_i_5 
       (.I0(p_0_out[16]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[19]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[19]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [19]),
        .I5(fdiv_rem[19]),
        .O(\rem[19]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[18]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [18]),
        .I5(fdiv_rem[18]),
        .O(\rem[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[17]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [17]),
        .I5(fdiv_rem[17]),
        .O(\rem[19]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[19]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[16]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [16]),
        .I5(fdiv_rem[16]),
        .O(\rem[19]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_2 
       (.I0(p_0_out[23]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_3 
       (.I0(p_0_out[22]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_4 
       (.I0(p_0_out[21]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[23]_i_5 
       (.I0(p_0_out[20]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[23]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[23]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [23]),
        .I5(fdiv_rem[23]),
        .O(\rem[23]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[22]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [22]),
        .I5(fdiv_rem[22]),
        .O(\rem[23]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[21]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [21]),
        .I5(fdiv_rem[21]),
        .O(\rem[23]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[23]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[20]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [20]),
        .I5(fdiv_rem[20]),
        .O(\rem[23]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_2 
       (.I0(p_0_out[27]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_3 
       (.I0(p_0_out[26]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_4 
       (.I0(p_0_out[25]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[27]_i_5 
       (.I0(p_0_out[24]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[27]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[27]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [27]),
        .I5(fdiv_rem[27]),
        .O(\rem[27]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[26]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [26]),
        .I5(fdiv_rem[26]),
        .O(\rem[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[25]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [25]),
        .I5(fdiv_rem[25]),
        .O(\rem[27]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[27]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[24]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [24]),
        .I5(fdiv_rem[24]),
        .O(\rem[27]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0D000000FFFFFFFF)) 
    \rem[31]_i_1 
       (.I0(dctl_long),
        .I1(dctl_stat[2]),
        .I2(dctl_stat[3]),
        .I3(dctl_stat[0]),
        .I4(dctl_stat[1]),
        .I5(\rem[31]_i_3_n_0 ),
        .O(\dctl_stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_10 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[28]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [28]),
        .I5(fdiv_rem[28]),
        .O(\rem[31]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_11 
       (.I0(chg_rem_sgn),
        .I1(chg_quo_sgn),
        .O(\rem[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h3F110FFF33110011)) 
    \rem[31]_i_12 
       (.I0(\rem_reg[31]_0 [31]),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(Q[31]),
        .I3(add_out0_carry_i_9_n_0),
        .I4(add_out0_carry__6[31]),
        .I5(add_out0_carry_i_10_n_0),
        .O(p_0_out[31]));
  LUT6 #(
    .INIT(64'hFD77FD77FD7FFF7F)) 
    \rem[31]_i_3 
       (.I0(dctl_stat[3]),
        .I1(dctl_stat[1]),
        .I2(dctl_stat[0]),
        .I3(dctl_stat[2]),
        .I4(fdiv_rem_msb_f),
        .I5(\rem[31]_i_11_n_0 ),
        .O(\rem[31]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_4 
       (.I0(p_0_out[30]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_5 
       (.I0(p_0_out[29]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[31]_i_6 
       (.I0(p_0_out[28]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[31]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [31]),
        .I5(fdiv_rem[31]),
        .O(\rem[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[30]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [30]),
        .I5(fdiv_rem[30]),
        .O(\rem[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[31]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[29]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [29]),
        .I5(fdiv_rem[29]),
        .O(\rem[31]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_2 
       (.I0(p_0_out[3]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_3 
       (.I0(p_0_out[2]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_4 
       (.I0(p_0_out[1]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[3]_i_5 
       (.I0(p_0_out[0]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[3]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[3]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[3]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [3]),
        .I5(fdiv_rem[3]),
        .O(\rem[3]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[3]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[2]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [2]),
        .I5(fdiv_rem[2]),
        .O(\rem[3]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[3]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[1]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [1]),
        .I5(fdiv_rem[1]),
        .O(\rem[3]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFF590059)) 
    \rem[3]_i_9 
       (.I0(p_0_out[0]),
        .I1(add_out0_carry_i_9_n_0),
        .I2(\rem_reg[31]_0 [0]),
        .I3(\rem[31]_i_3_n_0 ),
        .I4(fdiv_rem[0]),
        .O(\rem[3]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_2 
       (.I0(p_0_out[7]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_3 
       (.I0(p_0_out[6]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_4 
       (.I0(p_0_out[5]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \rem[7]_i_5 
       (.I0(p_0_out[4]),
        .I1(\rem[31]_i_3_n_0 ),
        .O(\rem[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_6 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[7]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [7]),
        .I5(fdiv_rem[7]),
        .O(\rem[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_7 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[6]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [6]),
        .I5(fdiv_rem[6]),
        .O(\rem[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_8 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[5]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [5]),
        .I5(fdiv_rem[5]),
        .O(\rem[7]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFCDEFCFC30123030)) 
    \rem[7]_i_9 
       (.I0(add_out0_carry_i_9_n_0),
        .I1(\rem[31]_i_3_n_0 ),
        .I2(p_0_out[4]),
        .I3(add_out0_carry_i_10_n_0),
        .I4(\rem_reg[31]_0 [4]),
        .I5(fdiv_rem[4]),
        .O(\rem[7]_i_9_n_0 ));
  CARRY4 \rem_reg[11]_i_1 
       (.CI(\rem_reg[7]_i_1_n_0 ),
        .CO({\rem_reg[11]_i_1_n_0 ,\rem_reg[11]_i_1_n_1 ,\rem_reg[11]_i_1_n_2 ,\rem_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[11]_i_2_n_0 ,\rem[11]_i_3_n_0 ,\rem[11]_i_4_n_0 ,\rem[11]_i_5_n_0 }),
        .O(\rem_reg[31] [11:8]),
        .S({\rem[11]_i_6_n_0 ,\rem[11]_i_7_n_0 ,\rem[11]_i_8_n_0 ,\rem[11]_i_9_n_0 }));
  CARRY4 \rem_reg[15]_i_1 
       (.CI(\rem_reg[11]_i_1_n_0 ),
        .CO({\rem_reg[15]_i_1_n_0 ,\rem_reg[15]_i_1_n_1 ,\rem_reg[15]_i_1_n_2 ,\rem_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[15]_i_2_n_0 ,\rem[15]_i_3_n_0 ,\rem[15]_i_4_n_0 ,\rem[15]_i_5_n_0 }),
        .O(\rem_reg[31] [15:12]),
        .S({\rem[15]_i_6_n_0 ,\rem[15]_i_7_n_0 ,\rem[15]_i_8_n_0 ,\rem[15]_i_9_n_0 }));
  CARRY4 \rem_reg[19]_i_1 
       (.CI(\rem_reg[15]_i_1_n_0 ),
        .CO({\rem_reg[19]_i_1_n_0 ,\rem_reg[19]_i_1_n_1 ,\rem_reg[19]_i_1_n_2 ,\rem_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[19]_i_2_n_0 ,\rem[19]_i_3_n_0 ,\rem[19]_i_4_n_0 ,\rem[19]_i_5_n_0 }),
        .O(\rem_reg[31] [19:16]),
        .S({\rem[19]_i_6_n_0 ,\rem[19]_i_7_n_0 ,\rem[19]_i_8_n_0 ,\rem[19]_i_9_n_0 }));
  CARRY4 \rem_reg[23]_i_1 
       (.CI(\rem_reg[19]_i_1_n_0 ),
        .CO({\rem_reg[23]_i_1_n_0 ,\rem_reg[23]_i_1_n_1 ,\rem_reg[23]_i_1_n_2 ,\rem_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[23]_i_2_n_0 ,\rem[23]_i_3_n_0 ,\rem[23]_i_4_n_0 ,\rem[23]_i_5_n_0 }),
        .O(\rem_reg[31] [23:20]),
        .S({\rem[23]_i_6_n_0 ,\rem[23]_i_7_n_0 ,\rem[23]_i_8_n_0 ,\rem[23]_i_9_n_0 }));
  CARRY4 \rem_reg[27]_i_1 
       (.CI(\rem_reg[23]_i_1_n_0 ),
        .CO({\rem_reg[27]_i_1_n_0 ,\rem_reg[27]_i_1_n_1 ,\rem_reg[27]_i_1_n_2 ,\rem_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[27]_i_2_n_0 ,\rem[27]_i_3_n_0 ,\rem[27]_i_4_n_0 ,\rem[27]_i_5_n_0 }),
        .O(\rem_reg[31] [27:24]),
        .S({\rem[27]_i_6_n_0 ,\rem[27]_i_7_n_0 ,\rem[27]_i_8_n_0 ,\rem[27]_i_9_n_0 }));
  CARRY4 \rem_reg[31]_i_2 
       (.CI(\rem_reg[27]_i_1_n_0 ),
        .CO({\rem_reg[31]_i_2_n_1 ,\rem_reg[31]_i_2_n_2 ,\rem_reg[31]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\rem[31]_i_4_n_0 ,\rem[31]_i_5_n_0 ,\rem[31]_i_6_n_0 }),
        .O(\rem_reg[31] [31:28]),
        .S({\rem[31]_i_7_n_0 ,\rem[31]_i_8_n_0 ,\rem[31]_i_9_n_0 ,\rem[31]_i_10_n_0 }));
  CARRY4 \rem_reg[3]_i_1 
       (.CI(\<const0> ),
        .CO({\rem_reg[3]_i_1_n_0 ,\rem_reg[3]_i_1_n_1 ,\rem_reg[3]_i_1_n_2 ,\rem_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[3]_i_2_n_0 ,\rem[3]_i_3_n_0 ,\rem[3]_i_4_n_0 ,\rem[3]_i_5_n_0 }),
        .O(\rem_reg[31] [3:0]),
        .S({\rem[3]_i_6_n_0 ,\rem[3]_i_7_n_0 ,\rem[3]_i_8_n_0 ,\rem[3]_i_9_n_0 }));
  CARRY4 \rem_reg[7]_i_1 
       (.CI(\rem_reg[3]_i_1_n_0 ),
        .CO({\rem_reg[7]_i_1_n_0 ,\rem_reg[7]_i_1_n_1 ,\rem_reg[7]_i_1_n_2 ,\rem_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\rem[7]_i_2_n_0 ,\rem[7]_i_3_n_0 ,\rem[7]_i_4_n_0 ,\rem[7]_i_5_n_0 }),
        .O(\rem_reg[31] [7:4]),
        .S({\rem[7]_i_6_n_0 ,\rem[7]_i_7_n_0 ,\rem[7]_i_8_n_0 ,\rem[7]_i_9_n_0 }));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[0]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[0] ),
        .I2(rgf_sr_nh),
        .I3(\remden_reg[31] [0]),
        .I4(\dctl_stat_reg[3]_0 ),
        .I5(abus_0[0]),
        .O(rst_n_37));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[10]_i_1 
       (.I0(\remden_reg[31] [10]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[10]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[10] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_4 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[11]_i_1 
       (.I0(\remden_reg[31] [11]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[11]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[11] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[12]_i_1 
       (.I0(\remden_reg[31] [12]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[12]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[12] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[13]_i_1 
       (.I0(\remden_reg[31] [13]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[13]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[13] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[14]_i_1 
       (.I0(\remden_reg[31] [14]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[14]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[14] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[15]_i_1 
       (.I0(\dctl_stat_reg[1]_0 ),
        .I1(rst_n),
        .O(rst_n_0));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[15]_i_2 
       (.I0(\remden_reg[31] [15]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[15]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[15] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8] ));
  LUT4 #(
    .INIT(16'hA202)) 
    \remden[19]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[19] ),
        .I2(\dctl_stat_reg[3]_0 ),
        .I3(\remden_reg[31] [16]),
        .O(rst_n_33));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[1]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[0] ),
        .I2(rgf_sr_nh),
        .I3(\remden_reg[31] [1]),
        .I4(\dctl_stat_reg[3]_0 ),
        .I5(abus_0[1]),
        .O(rst_n_36));
  LUT4 #(
    .INIT(16'h8A80)) 
    \remden[29]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[31] [18]),
        .I2(\dctl_stat_reg[3]_0 ),
        .I3(\remden_reg[29] ),
        .O(rst_n_31));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[2]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[0] ),
        .I2(rgf_sr_nh),
        .I3(\remden_reg[31] [2]),
        .I4(\dctl_stat_reg[3]_0 ),
        .I5(abus_0[2]),
        .O(rst_n_35));
  LUT4 #(
    .INIT(16'hA202)) 
    \remden[30]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[30] ),
        .I2(\dctl_stat_reg[3]_0 ),
        .I3(\remden_reg[31] [19]),
        .O(rst_n_32));
  LUT6 #(
    .INIT(64'h8A8A80808A808A80)) 
    \remden[31]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[31] [20]),
        .I2(\dctl_stat_reg[3]_0 ),
        .I3(\remden_reg[31]_0 ),
        .I4(\remden_reg[31]_1 ),
        .I5(\remden_reg[0] ),
        .O(rst_n_30));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[32]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[0]),
        .I2(\remden_reg[64] ),
        .O(\remden_reg[28]_2 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[33]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[1]),
        .I2(\remden_reg[64] ),
        .O(\remden_reg[28]_1 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[34]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[2]),
        .I2(\remden_reg[64] ),
        .O(\remden_reg[28]_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[35]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[3]),
        .I2(\remden_reg[64] ),
        .O(\remden_reg[28] ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[36]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[4]),
        .I2(\remden_reg[64] ),
        .O(rst_n_29));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[37]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[5]),
        .I2(\remden_reg[64] ),
        .O(rst_n_28));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[38]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[6]),
        .I2(\remden_reg[64] ),
        .O(rst_n_27));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[39]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[7]),
        .I2(\remden_reg[64] ),
        .O(rst_n_26));
  LUT6 #(
    .INIT(64'hAA008080AA000000)) 
    \remden[3]_i_1 
       (.I0(rst_n),
        .I1(\remden_reg[0] ),
        .I2(rgf_sr_nh),
        .I3(\remden_reg[31] [3]),
        .I4(\dctl_stat_reg[3]_0 ),
        .I5(abus_0[3]),
        .O(rst_n_34));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[40]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[8]),
        .I2(\remden_reg[64] ),
        .O(rst_n_25));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[41]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[9]),
        .I2(\remden_reg[64] ),
        .O(rst_n_24));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[42]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[10]),
        .I2(\remden_reg[64] ),
        .O(rst_n_23));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[43]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[11]),
        .I2(\remden_reg[64] ),
        .O(rst_n_22));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[44]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[12]),
        .I2(\remden_reg[64] ),
        .O(rst_n_21));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[45]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[13]),
        .I2(\remden_reg[64] ),
        .O(rst_n_20));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[46]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[14]),
        .I2(\remden_reg[64] ),
        .O(rst_n_19));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[47]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[15]),
        .I2(\remden_reg[64] ),
        .O(rst_n_18));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[48]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[16]),
        .I2(\remden_reg[64] ),
        .O(rst_n_17));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[49]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[17]),
        .I2(\remden_reg[64] ),
        .O(rst_n_16));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[4]_i_1 
       (.I0(\remden_reg[31] [4]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[4]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[4] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_10 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[50]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[18]),
        .I2(\remden_reg[64] ),
        .O(rst_n_15));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[51]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[19]),
        .I2(\remden_reg[64] ),
        .O(rst_n_14));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[52]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[20]),
        .I2(\remden_reg[64] ),
        .O(rst_n_13));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[53]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[21]),
        .I2(\remden_reg[64] ),
        .O(rst_n_12));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[54]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[22]),
        .I2(\remden_reg[64] ),
        .O(rst_n_11));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[55]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[23]),
        .I2(\remden_reg[64] ),
        .O(rst_n_10));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[56]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[24]),
        .I2(\remden_reg[64] ),
        .O(rst_n_9));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[57]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[25]),
        .I2(\remden_reg[64] ),
        .O(rst_n_8));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[58]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[26]),
        .I2(\remden_reg[64] ),
        .O(rst_n_7));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[59]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[27]),
        .I2(\remden_reg[64] ),
        .O(rst_n_6));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[5]_i_1 
       (.I0(\remden_reg[31] [5]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[5]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[5] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_9 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[60]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[28]),
        .I2(\remden_reg[64] ),
        .O(rst_n_5));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[61]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[29]),
        .I2(\remden_reg[64] ),
        .O(rst_n_4));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[62]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[30]),
        .I2(\remden_reg[64] ),
        .O(rst_n_3));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[63]_i_1 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem[31]),
        .I2(\remden_reg[64] ),
        .O(rst_n_2));
  LUT4 #(
    .INIT(16'hFFF1)) 
    \remden[64]_i_1 
       (.I0(\remden[64]_i_3_n_0 ),
        .I1(dctl_stat[1]),
        .I2(\remden[64]_i_4_n_0 ),
        .I3(\dctl_stat_reg[3]_0 ),
        .O(\dctl_stat_reg[1]_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \remden[64]_i_2 
       (.I0(\dctl_stat_reg[3]_0 ),
        .I1(fdiv_rem_msb_f_reg_0),
        .I2(\remden_reg[64] ),
        .O(rst_n_1));
  LUT6 #(
    .INIT(64'hD5000055F5550055)) 
    \remden[64]_i_3 
       (.I0(dctl_stat[0]),
        .I1(den2),
        .I2(dctl_sign),
        .I3(dctl_stat[2]),
        .I4(dctl_stat[3]),
        .I5(chg_quo_sgn_reg_0),
        .O(\remden[64]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAABAAAFEAABAAABA)) 
    \remden[64]_i_4 
       (.I0(\remden_reg[64] ),
        .I1(dctl_stat[0]),
        .I2(dctl_stat[1]),
        .I3(dctl_stat[3]),
        .I4(dctl_stat[2]),
        .I5(dctl_long),
        .O(\remden[64]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \remden[64]_i_5 
       (.I0(\rem[31]_i_3_n_0 ),
        .I1(\remden[64]_i_7_n_0 ),
        .O(\dctl_stat_reg[3]_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \remden[64]_i_7 
       (.I0(add_out0_carry_i_10_n_0),
        .I1(add_out0_carry_i_9_n_0),
        .O(\remden[64]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[6]_i_1 
       (.I0(\remden_reg[31] [6]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[6]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[6] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_8 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[7]_i_1 
       (.I0(\remden_reg[31] [7]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[7]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[7] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_7 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[8]_i_1 
       (.I0(\remden_reg[31] [8]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(rgf_sr_nh),
        .I3(abus_0[8]),
        .I4(\remden_reg[8] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_6 ));
  LUT6 #(
    .INIT(64'hB888B888BBBB8888)) 
    \remden[9]_i_1 
       (.I0(\remden_reg[31] [9]),
        .I1(\dctl_stat_reg[3]_0 ),
        .I2(abus_0[9]),
        .I3(rgf_sr_nh),
        .I4(\remden_reg[9] ),
        .I5(\remden_reg[0] ),
        .O(\sr_reg[8]_5 ));
endmodule

module niho_div_reg_den
   (chg_rem_sgn0,
    DI,
    p_1_in5_in,
    S,
    \remden_reg[38]_0 ,
    \remden_reg[38]_1 ,
    \remden_reg[42]_0 ,
    \remden_reg[42]_1 ,
    \remden_reg[46]_0 ,
    \remden_reg[46]_1 ,
    \remden_reg[50]_0 ,
    \remden_reg[50]_1 ,
    \remden_reg[54]_0 ,
    \remden_reg[54]_1 ,
    \remden_reg[58]_0 ,
    \remden_reg[58]_1 ,
    \remden_reg[62]_0 ,
    \remden_reg[62]_1 ,
    \remden_reg[30]_0 ,
    \remden_reg[30]_1 ,
    \remden_reg[29]_0 ,
    \remden_reg[29]_1 ,
    \remden_reg[28]_0 ,
    \remden_reg[28]_1 ,
    \remden_reg[64]_0 ,
    \remden_reg[25]_0 ,
    \remden_reg[24]_0 ,
    \remden_reg[23]_0 ,
    \remden_reg[22]_0 ,
    \remden_reg[21]_0 ,
    \remden_reg[20]_0 ,
    \remden_reg[18]_0 ,
    \remden_reg[17]_0 ,
    \remden_reg[16]_0 ,
    \remden_reg[15]_0 ,
    \remden_reg[14]_0 ,
    \remden_reg[13]_0 ,
    \remden_reg[12]_0 ,
    \remden_reg[11]_0 ,
    \remden_reg[10]_0 ,
    \remden_reg[9]_0 ,
    \remden_reg[8]_0 ,
    \remden_reg[7]_0 ,
    \remden_reg[6]_0 ,
    \remden_reg[5]_0 ,
    \remden_reg[4]_0 ,
    \remden_reg[19]_0 ,
    \remden_reg[3]_0 ,
    \remden_reg[2]_0 ,
    \remden_reg[1]_0 ,
    \remden_reg[0]_0 ,
    \remden_reg[27]_0 ,
    \remden_reg[26]_0 ,
    dctl_sign,
    Q,
    O,
    rem1_carry,
    rem0_carry,
    \remden_reg[64]_1 ,
    \remden_reg[64]_2 ,
    clk,
    \remden_reg[63]_0 ,
    \remden_reg[62]_2 ,
    \remden_reg[61]_0 ,
    \remden_reg[60]_0 ,
    \remden_reg[59]_0 ,
    \remden_reg[58]_2 ,
    \remden_reg[57]_0 ,
    \remden_reg[56]_0 ,
    \remden_reg[55]_0 ,
    \remden_reg[54]_2 ,
    \remden_reg[53]_0 ,
    \remden_reg[52]_0 ,
    \remden_reg[51]_0 ,
    \remden_reg[50]_2 ,
    \remden_reg[49]_0 ,
    \remden_reg[48]_0 ,
    \remden_reg[47]_0 ,
    \remden_reg[46]_2 ,
    \remden_reg[45]_0 ,
    \remden_reg[44]_0 ,
    \remden_reg[43]_0 ,
    \remden_reg[42]_2 ,
    \remden_reg[41]_0 ,
    \remden_reg[40]_0 ,
    \remden_reg[39]_0 ,
    \remden_reg[38]_2 ,
    \remden_reg[37]_0 ,
    \remden_reg[36]_0 ,
    \remden_reg[35]_0 ,
    \remden_reg[34]_0 ,
    \remden_reg[33]_0 ,
    \remden_reg[32]_0 ,
    \remden_reg[31]_0 ,
    \remden_reg[29]_2 ,
    \remden_reg[25]_1 ,
    \remden_reg[24]_1 ,
    \remden_reg[23]_1 ,
    \remden_reg[22]_1 ,
    \remden_reg[21]_1 ,
    \remden_reg[20]_1 ,
    \remden_reg[18]_1 ,
    \remden_reg[17]_1 ,
    \remden_reg[16]_1 ,
    \remden_reg[4]_1 ,
    \remden_reg[15]_1 ,
    \remden_reg[14]_1 ,
    \remden_reg[13]_1 ,
    \remden_reg[12]_1 ,
    \remden_reg[11]_1 ,
    \remden_reg[10]_1 ,
    \remden_reg[9]_1 ,
    \remden_reg[8]_1 ,
    \remden_reg[7]_1 ,
    \remden_reg[6]_1 ,
    \remden_reg[5]_1 ,
    \remden_reg[4]_2 ,
    \remden_reg[30]_2 ,
    \remden_reg[19]_1 ,
    \remden_reg[3]_1 ,
    \remden_reg[2]_1 ,
    \remden_reg[1]_1 ,
    \remden_reg[0]_1 ,
    \remden_reg[28]_2 ,
    rst_n,
    \remden_reg[28]_3 ,
    \remden_reg[28]_4 ,
    \remden_reg[27]_1 ,
    \remden_reg[26]_1 );
  output chg_rem_sgn0;
  output [3:0]DI;
  output [0:0]p_1_in5_in;
  output [3:0]S;
  output [3:0]\remden_reg[38]_0 ;
  output [3:0]\remden_reg[38]_1 ;
  output [3:0]\remden_reg[42]_0 ;
  output [3:0]\remden_reg[42]_1 ;
  output [3:0]\remden_reg[46]_0 ;
  output [3:0]\remden_reg[46]_1 ;
  output [3:0]\remden_reg[50]_0 ;
  output [3:0]\remden_reg[50]_1 ;
  output [3:0]\remden_reg[54]_0 ;
  output [3:0]\remden_reg[54]_1 ;
  output [3:0]\remden_reg[58]_0 ;
  output [3:0]\remden_reg[58]_1 ;
  output [3:0]\remden_reg[62]_0 ;
  output [3:0]\remden_reg[62]_1 ;
  output [0:0]\remden_reg[30]_0 ;
  output [0:0]\remden_reg[30]_1 ;
  output [0:0]\remden_reg[29]_0 ;
  output [0:0]\remden_reg[29]_1 ;
  output [0:0]\remden_reg[28]_0 ;
  output \remden_reg[28]_1 ;
  output [0:0]\remden_reg[64]_0 ;
  output \remden_reg[25]_0 ;
  output \remden_reg[24]_0 ;
  output \remden_reg[23]_0 ;
  output \remden_reg[22]_0 ;
  output \remden_reg[21]_0 ;
  output \remden_reg[20]_0 ;
  output \remden_reg[18]_0 ;
  output \remden_reg[17]_0 ;
  output \remden_reg[16]_0 ;
  output \remden_reg[15]_0 ;
  output \remden_reg[14]_0 ;
  output \remden_reg[13]_0 ;
  output \remden_reg[12]_0 ;
  output \remden_reg[11]_0 ;
  output \remden_reg[10]_0 ;
  output \remden_reg[9]_0 ;
  output \remden_reg[8]_0 ;
  output \remden_reg[7]_0 ;
  output \remden_reg[6]_0 ;
  output \remden_reg[5]_0 ;
  output \remden_reg[4]_0 ;
  output \remden_reg[19]_0 ;
  output \remden_reg[3]_0 ;
  output \remden_reg[2]_0 ;
  output \remden_reg[1]_0 ;
  output \remden_reg[0]_0 ;
  output \remden_reg[27]_0 ;
  output \remden_reg[26]_0 ;
  input dctl_sign;
  input [31:0]Q;
  input [0:0]O;
  input [0:0]rem1_carry;
  input [0:0]rem0_carry;
  input \remden_reg[64]_1 ;
  input \remden_reg[64]_2 ;
  input clk;
  input \remden_reg[63]_0 ;
  input \remden_reg[62]_2 ;
  input \remden_reg[61]_0 ;
  input \remden_reg[60]_0 ;
  input \remden_reg[59]_0 ;
  input \remden_reg[58]_2 ;
  input \remden_reg[57]_0 ;
  input \remden_reg[56]_0 ;
  input \remden_reg[55]_0 ;
  input \remden_reg[54]_2 ;
  input \remden_reg[53]_0 ;
  input \remden_reg[52]_0 ;
  input \remden_reg[51]_0 ;
  input \remden_reg[50]_2 ;
  input \remden_reg[49]_0 ;
  input \remden_reg[48]_0 ;
  input \remden_reg[47]_0 ;
  input \remden_reg[46]_2 ;
  input \remden_reg[45]_0 ;
  input \remden_reg[44]_0 ;
  input \remden_reg[43]_0 ;
  input \remden_reg[42]_2 ;
  input \remden_reg[41]_0 ;
  input \remden_reg[40]_0 ;
  input \remden_reg[39]_0 ;
  input \remden_reg[38]_2 ;
  input \remden_reg[37]_0 ;
  input \remden_reg[36]_0 ;
  input \remden_reg[35]_0 ;
  input \remden_reg[34]_0 ;
  input \remden_reg[33]_0 ;
  input \remden_reg[32]_0 ;
  input \remden_reg[31]_0 ;
  input \remden_reg[29]_2 ;
  input \remden_reg[25]_1 ;
  input \remden_reg[24]_1 ;
  input \remden_reg[23]_1 ;
  input \remden_reg[22]_1 ;
  input \remden_reg[21]_1 ;
  input \remden_reg[20]_1 ;
  input \remden_reg[18]_1 ;
  input \remden_reg[17]_1 ;
  input \remden_reg[16]_1 ;
  input \remden_reg[4]_1 ;
  input \remden_reg[15]_1 ;
  input \remden_reg[14]_1 ;
  input \remden_reg[13]_1 ;
  input \remden_reg[12]_1 ;
  input \remden_reg[11]_1 ;
  input \remden_reg[10]_1 ;
  input \remden_reg[9]_1 ;
  input \remden_reg[8]_1 ;
  input \remden_reg[7]_1 ;
  input \remden_reg[6]_1 ;
  input \remden_reg[5]_1 ;
  input \remden_reg[4]_2 ;
  input \remden_reg[30]_2 ;
  input \remden_reg[19]_1 ;
  input \remden_reg[3]_1 ;
  input \remden_reg[2]_1 ;
  input \remden_reg[1]_1 ;
  input \remden_reg[0]_1 ;
  input \remden_reg[28]_2 ;
  input rst_n;
  input \remden_reg[28]_3 ;
  input [2:0]\remden_reg[28]_4 ;
  input \remden_reg[27]_1 ;
  input \remden_reg[26]_1 ;

  wire \<const0> ;
  wire \<const1> ;
  wire [3:0]DI;
  wire [0:0]O;
  wire [31:0]Q;
  wire [3:0]S;
  wire chg_rem_sgn0;
  wire clk;
  wire dctl_sign;
  wire [0:0]p_1_in5_in;
  wire [0:0]rem0_carry;
  wire [0:0]rem1_carry;
  wire \remden[26]_i_1_n_0 ;
  wire \remden[27]_i_1_n_0 ;
  wire \remden[28]_i_1_n_0 ;
  wire \remden_reg[0]_0 ;
  wire \remden_reg[0]_1 ;
  wire \remden_reg[10]_0 ;
  wire \remden_reg[10]_1 ;
  wire \remden_reg[11]_0 ;
  wire \remden_reg[11]_1 ;
  wire \remden_reg[12]_0 ;
  wire \remden_reg[12]_1 ;
  wire \remden_reg[13]_0 ;
  wire \remden_reg[13]_1 ;
  wire \remden_reg[14]_0 ;
  wire \remden_reg[14]_1 ;
  wire \remden_reg[15]_0 ;
  wire \remden_reg[15]_1 ;
  wire \remden_reg[16]_0 ;
  wire \remden_reg[16]_1 ;
  wire \remden_reg[17]_0 ;
  wire \remden_reg[17]_1 ;
  wire \remden_reg[18]_0 ;
  wire \remden_reg[18]_1 ;
  wire \remden_reg[19]_0 ;
  wire \remden_reg[19]_1 ;
  wire \remden_reg[1]_0 ;
  wire \remden_reg[1]_1 ;
  wire \remden_reg[20]_0 ;
  wire \remden_reg[20]_1 ;
  wire \remden_reg[21]_0 ;
  wire \remden_reg[21]_1 ;
  wire \remden_reg[22]_0 ;
  wire \remden_reg[22]_1 ;
  wire \remden_reg[23]_0 ;
  wire \remden_reg[23]_1 ;
  wire \remden_reg[24]_0 ;
  wire \remden_reg[24]_1 ;
  wire \remden_reg[25]_0 ;
  wire \remden_reg[25]_1 ;
  wire \remden_reg[26]_0 ;
  wire \remden_reg[26]_1 ;
  wire \remden_reg[27]_0 ;
  wire \remden_reg[27]_1 ;
  wire [0:0]\remden_reg[28]_0 ;
  wire \remden_reg[28]_1 ;
  wire \remden_reg[28]_2 ;
  wire \remden_reg[28]_3 ;
  wire [2:0]\remden_reg[28]_4 ;
  wire [0:0]\remden_reg[29]_0 ;
  wire [0:0]\remden_reg[29]_1 ;
  wire \remden_reg[29]_2 ;
  wire \remden_reg[2]_0 ;
  wire \remden_reg[2]_1 ;
  wire [0:0]\remden_reg[30]_0 ;
  wire [0:0]\remden_reg[30]_1 ;
  wire \remden_reg[30]_2 ;
  wire \remden_reg[31]_0 ;
  wire \remden_reg[32]_0 ;
  wire \remden_reg[33]_0 ;
  wire \remden_reg[34]_0 ;
  wire \remden_reg[35]_0 ;
  wire \remden_reg[36]_0 ;
  wire \remden_reg[37]_0 ;
  wire [3:0]\remden_reg[38]_0 ;
  wire [3:0]\remden_reg[38]_1 ;
  wire \remden_reg[38]_2 ;
  wire \remden_reg[39]_0 ;
  wire \remden_reg[3]_0 ;
  wire \remden_reg[3]_1 ;
  wire \remden_reg[40]_0 ;
  wire \remden_reg[41]_0 ;
  wire [3:0]\remden_reg[42]_0 ;
  wire [3:0]\remden_reg[42]_1 ;
  wire \remden_reg[42]_2 ;
  wire \remden_reg[43]_0 ;
  wire \remden_reg[44]_0 ;
  wire \remden_reg[45]_0 ;
  wire [3:0]\remden_reg[46]_0 ;
  wire [3:0]\remden_reg[46]_1 ;
  wire \remden_reg[46]_2 ;
  wire \remden_reg[47]_0 ;
  wire \remden_reg[48]_0 ;
  wire \remden_reg[49]_0 ;
  wire \remden_reg[4]_0 ;
  wire \remden_reg[4]_1 ;
  wire \remden_reg[4]_2 ;
  wire [3:0]\remden_reg[50]_0 ;
  wire [3:0]\remden_reg[50]_1 ;
  wire \remden_reg[50]_2 ;
  wire \remden_reg[51]_0 ;
  wire \remden_reg[52]_0 ;
  wire \remden_reg[53]_0 ;
  wire [3:0]\remden_reg[54]_0 ;
  wire [3:0]\remden_reg[54]_1 ;
  wire \remden_reg[54]_2 ;
  wire \remden_reg[55]_0 ;
  wire \remden_reg[56]_0 ;
  wire \remden_reg[57]_0 ;
  wire [3:0]\remden_reg[58]_0 ;
  wire [3:0]\remden_reg[58]_1 ;
  wire \remden_reg[58]_2 ;
  wire \remden_reg[59]_0 ;
  wire \remden_reg[5]_0 ;
  wire \remden_reg[5]_1 ;
  wire \remden_reg[60]_0 ;
  wire \remden_reg[61]_0 ;
  wire [3:0]\remden_reg[62]_0 ;
  wire [3:0]\remden_reg[62]_1 ;
  wire \remden_reg[62]_2 ;
  wire \remden_reg[63]_0 ;
  wire [0:0]\remden_reg[64]_0 ;
  wire \remden_reg[64]_1 ;
  wire \remden_reg[64]_2 ;
  wire \remden_reg[6]_0 ;
  wire \remden_reg[6]_1 ;
  wire \remden_reg[7]_0 ;
  wire \remden_reg[7]_1 ;
  wire \remden_reg[8]_0 ;
  wire \remden_reg[8]_1 ;
  wire \remden_reg[9]_0 ;
  wire \remden_reg[9]_1 ;
  wire \remden_reg_n_0_[63] ;
  wire \remden_reg_n_0_[64] ;
  wire rst_n;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    chg_rem_sgn_i_2
       (.I0(DI[0]),
        .I1(dctl_sign),
        .O(chg_rem_sgn0));
  LUT3 #(
    .INIT(8'h69)) 
    rem0_carry_i_5
       (.I0(\remden_reg[28]_1 ),
        .I1(Q[0]),
        .I2(rem0_carry),
        .O(\remden_reg[28]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem1_carry_i_5
       (.I0(\remden_reg[29]_1 ),
        .I1(Q[0]),
        .I2(rem1_carry),
        .O(\remden_reg[29]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem2_carry_i_5
       (.I0(\remden_reg[30]_1 ),
        .I1(Q[0]),
        .I2(O),
        .O(\remden_reg[30]_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_1
       (.I0(\remden_reg[38]_1 [3]),
        .I1(Q[7]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[38]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_2
       (.I0(\remden_reg[38]_1 [2]),
        .I1(Q[6]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[38]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_3
       (.I0(\remden_reg[38]_1 [1]),
        .I1(Q[5]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[38]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__0_i_4
       (.I0(\remden_reg[38]_1 [0]),
        .I1(Q[4]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[38]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_1
       (.I0(\remden_reg[42]_1 [3]),
        .I1(Q[11]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[42]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_2
       (.I0(\remden_reg[42]_1 [2]),
        .I1(Q[10]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[42]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_3
       (.I0(\remden_reg[42]_1 [1]),
        .I1(Q[9]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[42]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__1_i_4
       (.I0(\remden_reg[42]_1 [0]),
        .I1(Q[8]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[42]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_1
       (.I0(\remden_reg[46]_1 [3]),
        .I1(\remden_reg_n_0_[64] ),
        .I2(Q[15]),
        .O(\remden_reg[46]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_2
       (.I0(\remden_reg[46]_1 [2]),
        .I1(Q[14]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[46]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_3
       (.I0(\remden_reg[46]_1 [1]),
        .I1(Q[13]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[46]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__2_i_4
       (.I0(\remden_reg[46]_1 [0]),
        .I1(Q[12]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[46]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_1
       (.I0(\remden_reg[50]_1 [3]),
        .I1(Q[19]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[50]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_2
       (.I0(\remden_reg[50]_1 [2]),
        .I1(Q[18]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[50]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_3
       (.I0(\remden_reg[50]_1 [1]),
        .I1(Q[17]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[50]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__3_i_4
       (.I0(\remden_reg[50]_1 [0]),
        .I1(Q[16]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[50]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_1
       (.I0(\remden_reg[54]_1 [3]),
        .I1(Q[23]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[54]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_2
       (.I0(\remden_reg[54]_1 [2]),
        .I1(Q[22]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[54]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_3
       (.I0(\remden_reg[54]_1 [1]),
        .I1(Q[21]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[54]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__4_i_4
       (.I0(\remden_reg[54]_1 [0]),
        .I1(Q[20]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[54]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_1
       (.I0(\remden_reg[58]_1 [3]),
        .I1(Q[27]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[58]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_2
       (.I0(\remden_reg[58]_1 [2]),
        .I1(Q[26]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[58]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_3
       (.I0(\remden_reg[58]_1 [1]),
        .I1(Q[25]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[58]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__5_i_4
       (.I0(\remden_reg[58]_1 [0]),
        .I1(Q[24]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[58]_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_1
       (.I0(\remden_reg[62]_1 [3]),
        .I1(\remden_reg_n_0_[64] ),
        .I2(Q[31]),
        .O(\remden_reg[62]_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_2
       (.I0(\remden_reg[62]_1 [2]),
        .I1(Q[30]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[62]_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_3
       (.I0(\remden_reg[62]_1 [1]),
        .I1(Q[29]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[62]_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry__6_i_4
       (.I0(\remden_reg[62]_1 [0]),
        .I1(Q[28]),
        .I2(\remden_reg_n_0_[64] ),
        .O(\remden_reg[62]_0 [0]));
  LUT2 #(
    .INIT(4'h9)) 
    rem3_carry__7_i_1
       (.I0(\remden_reg_n_0_[64] ),
        .I1(\remden_reg_n_0_[63] ),
        .O(\remden_reg[64]_0 ));
  LUT1 #(
    .INIT(2'h1)) 
    rem3_carry_i_1
       (.I0(\remden_reg_n_0_[64] ),
        .O(p_1_in5_in));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_2
       (.I0(DI[3]),
        .I1(Q[3]),
        .I2(\remden_reg_n_0_[64] ),
        .O(S[3]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_3
       (.I0(DI[2]),
        .I1(Q[2]),
        .I2(\remden_reg_n_0_[64] ),
        .O(S[2]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_4
       (.I0(DI[1]),
        .I1(Q[1]),
        .I2(\remden_reg_n_0_[64] ),
        .O(S[1]));
  LUT3 #(
    .INIT(8'h69)) 
    rem3_carry_i_5
       (.I0(DI[0]),
        .I1(Q[0]),
        .I2(\remden_reg_n_0_[64] ),
        .O(S[0]));
  LUT6 #(
    .INIT(64'hC404FFFFC4040000)) 
    \remden[26]_i_1 
       (.I0(\remden_reg[26]_1 ),
        .I1(rst_n),
        .I2(\remden_reg[28]_3 ),
        .I3(\remden_reg[28]_4 [0]),
        .I4(\remden_reg[64]_1 ),
        .I5(\remden_reg[26]_0 ),
        .O(\remden[26]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hC404FFFFC4040000)) 
    \remden[27]_i_1 
       (.I0(\remden_reg[27]_1 ),
        .I1(rst_n),
        .I2(\remden_reg[28]_3 ),
        .I3(\remden_reg[28]_4 [1]),
        .I4(\remden_reg[64]_1 ),
        .I5(\remden_reg[27]_0 ),
        .O(\remden[27]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hC404FFFFC4040000)) 
    \remden[28]_i_1 
       (.I0(\remden_reg[28]_2 ),
        .I1(rst_n),
        .I2(\remden_reg[28]_3 ),
        .I3(\remden_reg[28]_4 [2]),
        .I4(\remden_reg[64]_1 ),
        .I5(\remden_reg[28]_1 ),
        .O(\remden[28]_i_1_n_0 ));
  FDRE \remden_reg[0] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[0]_1 ),
        .Q(\remden_reg[0]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[10] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[10]_1 ),
        .Q(\remden_reg[10]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[11] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[11]_1 ),
        .Q(\remden_reg[11]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[12] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[12]_1 ),
        .Q(\remden_reg[12]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[13] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[13]_1 ),
        .Q(\remden_reg[13]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[14] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[14]_1 ),
        .Q(\remden_reg[14]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[15] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[15]_1 ),
        .Q(\remden_reg[15]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[16] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[16]_1 ),
        .Q(\remden_reg[16]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[17] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[17]_1 ),
        .Q(\remden_reg[17]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[18] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[18]_1 ),
        .Q(\remden_reg[18]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[19] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[19]_1 ),
        .Q(\remden_reg[19]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[1] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[1]_1 ),
        .Q(\remden_reg[1]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[20] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[20]_1 ),
        .Q(\remden_reg[20]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[21] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[21]_1 ),
        .Q(\remden_reg[21]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[22] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[22]_1 ),
        .Q(\remden_reg[22]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[23] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[23]_1 ),
        .Q(\remden_reg[23]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[24] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[24]_1 ),
        .Q(\remden_reg[24]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[25] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[25]_1 ),
        .Q(\remden_reg[25]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\remden[26]_i_1_n_0 ),
        .Q(\remden_reg[26]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\remden[27]_i_1_n_0 ),
        .Q(\remden_reg[27]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\remden[28]_i_1_n_0 ),
        .Q(\remden_reg[28]_1 ),
        .R(\<const0> ));
  FDRE \remden_reg[29] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[29]_2 ),
        .Q(\remden_reg[29]_1 ),
        .R(\<const0> ));
  FDRE \remden_reg[2] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[2]_1 ),
        .Q(\remden_reg[2]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[30] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[30]_2 ),
        .Q(\remden_reg[30]_1 ),
        .R(\<const0> ));
  FDRE \remden_reg[31] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[31]_0 ),
        .Q(DI[0]),
        .R(\<const0> ));
  FDRE \remden_reg[32] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[32]_0 ),
        .Q(DI[1]),
        .R(\<const0> ));
  FDRE \remden_reg[33] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[33]_0 ),
        .Q(DI[2]),
        .R(\<const0> ));
  FDRE \remden_reg[34] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[34]_0 ),
        .Q(DI[3]),
        .R(\<const0> ));
  FDRE \remden_reg[35] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[35]_0 ),
        .Q(\remden_reg[38]_1 [0]),
        .R(\<const0> ));
  FDRE \remden_reg[36] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[36]_0 ),
        .Q(\remden_reg[38]_1 [1]),
        .R(\<const0> ));
  FDRE \remden_reg[37] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[37]_0 ),
        .Q(\remden_reg[38]_1 [2]),
        .R(\<const0> ));
  FDRE \remden_reg[38] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[38]_2 ),
        .Q(\remden_reg[38]_1 [3]),
        .R(\<const0> ));
  FDRE \remden_reg[39] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[39]_0 ),
        .Q(\remden_reg[42]_1 [0]),
        .R(\<const0> ));
  FDRE \remden_reg[3] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[3]_1 ),
        .Q(\remden_reg[3]_0 ),
        .R(\<const0> ));
  FDRE \remden_reg[40] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[40]_0 ),
        .Q(\remden_reg[42]_1 [1]),
        .R(\<const0> ));
  FDRE \remden_reg[41] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[41]_0 ),
        .Q(\remden_reg[42]_1 [2]),
        .R(\<const0> ));
  FDRE \remden_reg[42] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[42]_2 ),
        .Q(\remden_reg[42]_1 [3]),
        .R(\<const0> ));
  FDRE \remden_reg[43] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[43]_0 ),
        .Q(\remden_reg[46]_1 [0]),
        .R(\<const0> ));
  FDRE \remden_reg[44] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[44]_0 ),
        .Q(\remden_reg[46]_1 [1]),
        .R(\<const0> ));
  FDRE \remden_reg[45] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[45]_0 ),
        .Q(\remden_reg[46]_1 [2]),
        .R(\<const0> ));
  FDRE \remden_reg[46] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[46]_2 ),
        .Q(\remden_reg[46]_1 [3]),
        .R(\<const0> ));
  FDRE \remden_reg[47] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[47]_0 ),
        .Q(\remden_reg[50]_1 [0]),
        .R(\<const0> ));
  FDRE \remden_reg[48] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[48]_0 ),
        .Q(\remden_reg[50]_1 [1]),
        .R(\<const0> ));
  FDRE \remden_reg[49] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[49]_0 ),
        .Q(\remden_reg[50]_1 [2]),
        .R(\<const0> ));
  FDRE \remden_reg[4] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[4]_2 ),
        .Q(\remden_reg[4]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[50] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[50]_2 ),
        .Q(\remden_reg[50]_1 [3]),
        .R(\<const0> ));
  FDRE \remden_reg[51] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[51]_0 ),
        .Q(\remden_reg[54]_1 [0]),
        .R(\<const0> ));
  FDRE \remden_reg[52] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[52]_0 ),
        .Q(\remden_reg[54]_1 [1]),
        .R(\<const0> ));
  FDRE \remden_reg[53] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[53]_0 ),
        .Q(\remden_reg[54]_1 [2]),
        .R(\<const0> ));
  FDRE \remden_reg[54] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[54]_2 ),
        .Q(\remden_reg[54]_1 [3]),
        .R(\<const0> ));
  FDRE \remden_reg[55] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[55]_0 ),
        .Q(\remden_reg[58]_1 [0]),
        .R(\<const0> ));
  FDRE \remden_reg[56] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[56]_0 ),
        .Q(\remden_reg[58]_1 [1]),
        .R(\<const0> ));
  FDRE \remden_reg[57] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[57]_0 ),
        .Q(\remden_reg[58]_1 [2]),
        .R(\<const0> ));
  FDRE \remden_reg[58] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[58]_2 ),
        .Q(\remden_reg[58]_1 [3]),
        .R(\<const0> ));
  FDRE \remden_reg[59] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[59]_0 ),
        .Q(\remden_reg[62]_1 [0]),
        .R(\<const0> ));
  FDRE \remden_reg[5] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[5]_1 ),
        .Q(\remden_reg[5]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[60] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[60]_0 ),
        .Q(\remden_reg[62]_1 [1]),
        .R(\<const0> ));
  FDRE \remden_reg[61] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[61]_0 ),
        .Q(\remden_reg[62]_1 [2]),
        .R(\<const0> ));
  FDRE \remden_reg[62] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[62]_2 ),
        .Q(\remden_reg[62]_1 [3]),
        .R(\<const0> ));
  FDRE \remden_reg[63] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[63]_0 ),
        .Q(\remden_reg_n_0_[63] ),
        .R(\<const0> ));
  FDRE \remden_reg[64] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[64]_2 ),
        .Q(\remden_reg_n_0_[64] ),
        .R(\<const0> ));
  FDRE \remden_reg[6] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[6]_1 ),
        .Q(\remden_reg[6]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[7] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[7]_1 ),
        .Q(\remden_reg[7]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[8] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[8]_1 ),
        .Q(\remden_reg[8]_0 ),
        .R(\remden_reg[4]_1 ));
  FDRE \remden_reg[9] 
       (.C(clk),
        .CE(\remden_reg[64]_1 ),
        .D(\remden_reg[9]_1 ),
        .Q(\remden_reg[9]_0 ),
        .R(\remden_reg[4]_1 ));
endmodule

module niho_div_reg_dso
   (\remden_reg[31] ,
    \dso_reg[31]_0 ,
    Q,
    dctl_sign,
    DI,
    rgf_sr_nh,
    chg_quo_sgn_reg,
    dctl_long_f,
    p_0_in,
    E,
    D,
    clk);
  output \remden_reg[31] ;
  output \dso_reg[31]_0 ;
  output [31:0]Q;
  input dctl_sign;
  input [0:0]DI;
  input rgf_sr_nh;
  input chg_quo_sgn_reg;
  input dctl_long_f;
  input p_0_in;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]DI;
  wire [0:0]E;
  wire [31:0]Q;
  wire chg_quo_sgn_reg;
  wire clk;
  wire dctl_long_f;
  wire dctl_sign;
  wire \dso_reg[31]_0 ;
  wire p_0_in;
  wire \remden_reg[31] ;
  wire rgf_sr_nh;

  LUT5 #(
    .INIT(32'h4540757F)) 
    chg_quo_sgn_i_2
       (.I0(Q[31]),
        .I1(rgf_sr_nh),
        .I2(chg_quo_sgn_reg),
        .I3(dctl_long_f),
        .I4(Q[15]),
        .O(\dso_reg[31]_0 ));
  LUT3 #(
    .INIT(8'h3B)) 
    \dctl_stat[3]_i_2 
       (.I0(\dso_reg[31]_0 ),
        .I1(dctl_sign),
        .I2(DI),
        .O(\remden_reg[31] ));
  FDRE \dso_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in));
  FDRE \dso_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(p_0_in));
  FDRE \dso_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(p_0_in));
  FDRE \dso_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(p_0_in));
  FDRE \dso_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(p_0_in));
  FDRE \dso_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(p_0_in));
  FDRE \dso_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(p_0_in));
  FDRE \dso_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(Q[16]),
        .R(p_0_in));
  FDRE \dso_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(Q[17]),
        .R(p_0_in));
  FDRE \dso_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(Q[18]),
        .R(p_0_in));
  FDRE \dso_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(Q[19]),
        .R(p_0_in));
  FDRE \dso_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in));
  FDRE \dso_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(Q[20]),
        .R(p_0_in));
  FDRE \dso_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(Q[21]),
        .R(p_0_in));
  FDRE \dso_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(Q[22]),
        .R(p_0_in));
  FDRE \dso_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(Q[23]),
        .R(p_0_in));
  FDRE \dso_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(Q[24]),
        .R(p_0_in));
  FDRE \dso_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(Q[25]),
        .R(p_0_in));
  FDRE \dso_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(Q[26]),
        .R(p_0_in));
  FDRE \dso_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(Q[27]),
        .R(p_0_in));
  FDRE \dso_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(Q[28]),
        .R(p_0_in));
  FDRE \dso_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(Q[29]),
        .R(p_0_in));
  FDRE \dso_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in));
  FDRE \dso_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(Q[30]),
        .R(p_0_in));
  FDRE \dso_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(Q[31]),
        .R(p_0_in));
  FDRE \dso_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(p_0_in));
  FDRE \dso_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(p_0_in));
  FDRE \dso_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(p_0_in));
  FDRE \dso_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(p_0_in));
  FDRE \dso_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(p_0_in));
  FDRE \dso_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(p_0_in));
  FDRE \dso_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(p_0_in));
endmodule

module niho_div_reg_quo
   (\niho_dsp_c[31] ,
    Q,
    \tr[31]_i_5 ,
    niho_dsp_c,
    \tr[31]_i_5_0 ,
    \tr[31]_i_5_1 ,
    \tr[31]_i_5_2 ,
    p_0_in,
    E,
    D,
    clk);
  output \niho_dsp_c[31] ;
  output [31:0]Q;
  input \tr[31]_i_5 ;
  input [0:0]niho_dsp_c;
  input \tr[31]_i_5_0 ;
  input [0:0]\tr[31]_i_5_1 ;
  input \tr[31]_i_5_2 ;
  input p_0_in;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire [31:0]Q;
  wire clk;
  wire [0:0]niho_dsp_c;
  wire \niho_dsp_c[31] ;
  wire p_0_in;
  wire \tr[31]_i_5 ;
  wire \tr[31]_i_5_0 ;
  wire [0:0]\tr[31]_i_5_1 ;
  wire \tr[31]_i_5_2 ;

  FDRE \quo_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in));
  FDRE \quo_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(p_0_in));
  FDRE \quo_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(p_0_in));
  FDRE \quo_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(p_0_in));
  FDRE \quo_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(p_0_in));
  FDRE \quo_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(p_0_in));
  FDRE \quo_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(p_0_in));
  FDRE \quo_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(Q[16]),
        .R(p_0_in));
  FDRE \quo_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(Q[17]),
        .R(p_0_in));
  FDRE \quo_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(Q[18]),
        .R(p_0_in));
  FDRE \quo_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(Q[19]),
        .R(p_0_in));
  FDRE \quo_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in));
  FDRE \quo_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(Q[20]),
        .R(p_0_in));
  FDRE \quo_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(Q[21]),
        .R(p_0_in));
  FDRE \quo_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(Q[22]),
        .R(p_0_in));
  FDRE \quo_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(Q[23]),
        .R(p_0_in));
  FDRE \quo_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(Q[24]),
        .R(p_0_in));
  FDRE \quo_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(Q[25]),
        .R(p_0_in));
  FDRE \quo_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(Q[26]),
        .R(p_0_in));
  FDRE \quo_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(Q[27]),
        .R(p_0_in));
  FDRE \quo_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(Q[28]),
        .R(p_0_in));
  FDRE \quo_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(Q[29]),
        .R(p_0_in));
  FDRE \quo_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in));
  FDRE \quo_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(Q[30]),
        .R(p_0_in));
  FDRE \quo_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(Q[31]),
        .R(p_0_in));
  FDRE \quo_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(p_0_in));
  FDRE \quo_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(p_0_in));
  FDRE \quo_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(p_0_in));
  FDRE \quo_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(p_0_in));
  FDRE \quo_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(p_0_in));
  FDRE \quo_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(p_0_in));
  FDRE \quo_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(p_0_in));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[31]_i_14 
       (.I0(\tr[31]_i_5 ),
        .I1(niho_dsp_c),
        .I2(Q[31]),
        .I3(\tr[31]_i_5_0 ),
        .I4(\tr[31]_i_5_1 ),
        .I5(\tr[31]_i_5_2 ),
        .O(\niho_dsp_c[31] ));
endmodule

module niho_div_reg_rem
   (Q,
    p_0_in,
    E,
    D,
    clk);
  output [31:0]Q;
  input p_0_in;
  input [0:0]E;
  input [31:0]D;
  input clk;

  wire [31:0]D;
  wire [0:0]E;
  wire [31:0]Q;
  wire clk;
  wire p_0_in;

  FDRE \rem_reg[0] 
       (.C(clk),
        .CE(E),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in));
  FDRE \rem_reg[10] 
       (.C(clk),
        .CE(E),
        .D(D[10]),
        .Q(Q[10]),
        .R(p_0_in));
  FDRE \rem_reg[11] 
       (.C(clk),
        .CE(E),
        .D(D[11]),
        .Q(Q[11]),
        .R(p_0_in));
  FDRE \rem_reg[12] 
       (.C(clk),
        .CE(E),
        .D(D[12]),
        .Q(Q[12]),
        .R(p_0_in));
  FDRE \rem_reg[13] 
       (.C(clk),
        .CE(E),
        .D(D[13]),
        .Q(Q[13]),
        .R(p_0_in));
  FDRE \rem_reg[14] 
       (.C(clk),
        .CE(E),
        .D(D[14]),
        .Q(Q[14]),
        .R(p_0_in));
  FDRE \rem_reg[15] 
       (.C(clk),
        .CE(E),
        .D(D[15]),
        .Q(Q[15]),
        .R(p_0_in));
  FDRE \rem_reg[16] 
       (.C(clk),
        .CE(E),
        .D(D[16]),
        .Q(Q[16]),
        .R(p_0_in));
  FDRE \rem_reg[17] 
       (.C(clk),
        .CE(E),
        .D(D[17]),
        .Q(Q[17]),
        .R(p_0_in));
  FDRE \rem_reg[18] 
       (.C(clk),
        .CE(E),
        .D(D[18]),
        .Q(Q[18]),
        .R(p_0_in));
  FDRE \rem_reg[19] 
       (.C(clk),
        .CE(E),
        .D(D[19]),
        .Q(Q[19]),
        .R(p_0_in));
  FDRE \rem_reg[1] 
       (.C(clk),
        .CE(E),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in));
  FDRE \rem_reg[20] 
       (.C(clk),
        .CE(E),
        .D(D[20]),
        .Q(Q[20]),
        .R(p_0_in));
  FDRE \rem_reg[21] 
       (.C(clk),
        .CE(E),
        .D(D[21]),
        .Q(Q[21]),
        .R(p_0_in));
  FDRE \rem_reg[22] 
       (.C(clk),
        .CE(E),
        .D(D[22]),
        .Q(Q[22]),
        .R(p_0_in));
  FDRE \rem_reg[23] 
       (.C(clk),
        .CE(E),
        .D(D[23]),
        .Q(Q[23]),
        .R(p_0_in));
  FDRE \rem_reg[24] 
       (.C(clk),
        .CE(E),
        .D(D[24]),
        .Q(Q[24]),
        .R(p_0_in));
  FDRE \rem_reg[25] 
       (.C(clk),
        .CE(E),
        .D(D[25]),
        .Q(Q[25]),
        .R(p_0_in));
  FDRE \rem_reg[26] 
       (.C(clk),
        .CE(E),
        .D(D[26]),
        .Q(Q[26]),
        .R(p_0_in));
  FDRE \rem_reg[27] 
       (.C(clk),
        .CE(E),
        .D(D[27]),
        .Q(Q[27]),
        .R(p_0_in));
  FDRE \rem_reg[28] 
       (.C(clk),
        .CE(E),
        .D(D[28]),
        .Q(Q[28]),
        .R(p_0_in));
  FDRE \rem_reg[29] 
       (.C(clk),
        .CE(E),
        .D(D[29]),
        .Q(Q[29]),
        .R(p_0_in));
  FDRE \rem_reg[2] 
       (.C(clk),
        .CE(E),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in));
  FDRE \rem_reg[30] 
       (.C(clk),
        .CE(E),
        .D(D[30]),
        .Q(Q[30]),
        .R(p_0_in));
  FDRE \rem_reg[31] 
       (.C(clk),
        .CE(E),
        .D(D[31]),
        .Q(Q[31]),
        .R(p_0_in));
  FDRE \rem_reg[3] 
       (.C(clk),
        .CE(E),
        .D(D[3]),
        .Q(Q[3]),
        .R(p_0_in));
  FDRE \rem_reg[4] 
       (.C(clk),
        .CE(E),
        .D(D[4]),
        .Q(Q[4]),
        .R(p_0_in));
  FDRE \rem_reg[5] 
       (.C(clk),
        .CE(E),
        .D(D[5]),
        .Q(Q[5]),
        .R(p_0_in));
  FDRE \rem_reg[6] 
       (.C(clk),
        .CE(E),
        .D(D[6]),
        .Q(Q[6]),
        .R(p_0_in));
  FDRE \rem_reg[7] 
       (.C(clk),
        .CE(E),
        .D(D[7]),
        .Q(Q[7]),
        .R(p_0_in));
  FDRE \rem_reg[8] 
       (.C(clk),
        .CE(E),
        .D(D[8]),
        .Q(Q[8]),
        .R(p_0_in));
  FDRE \rem_reg[9] 
       (.C(clk),
        .CE(E),
        .D(D[9]),
        .Q(Q[9]),
        .R(p_0_in));
endmodule

module niho_fch
   (.out({ir[15],ir[14],ir[13],ir[12],ir[11],ir[10],ir[7],ir[6],ir[3],ir[0]}),
    \sr_reg[8] ,
    \sr_reg[4] ,
    \sr_reg[5] ,
    cbus,
    \sr_reg[11] ,
    \stat_reg[2] ,
    \sr_reg[10] ,
    \sr_reg[8]_0 ,
    \sr_reg[1] ,
    \sr_reg[2] ,
    \sr_reg[3] ,
    \sr_reg[0] ,
    bbus_sr,
    bbus_sel_cr,
    D,
    \cbus_i[30] ,
    \stat_reg[2]_0 ,
    ctl_sp_inc,
    \tr[31]_i_44_0 ,
    \sr[6]_i_25_0 ,
    \stat_reg[0] ,
    \stat_reg[0]_0 ,
    \stat_reg[0]_1 ,
    bbus_0,
    \tr[29]_i_14_0 ,
    \tr[28]_i_13_0 ,
    rst_n_fl_reg_0,
    \stat_reg[2]_1 ,
    \stat_reg[0]_2 ,
    \tr[21]_i_14_0 ,
    \tr[23]_i_15_0 ,
    \tr[27]_i_14 ,
    \niho_dsp_a[15]_INST_0_i_2_0 ,
    \tr[19]_i_14_0 ,
    \niho_dsp_a[32]_INST_0_i_5_0 ,
    \niho_dsp_a[32]_INST_0_i_5_1 ,
    \stat_reg[2]_2 ,
    \sr_reg[8]_1 ,
    \niho_dsp_a[32]_INST_0_i_7_0 ,
    \iv[3]_i_16 ,
    \iv[12]_i_10 ,
    \iv[15]_i_19_0 ,
    \sr[4]_i_40_0 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr[7]_i_21 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \iv[0]_i_27_0 ,
    \iv[8]_i_34_0 ,
    \sr[7]_i_20_0 ,
    \iv[9]_i_35 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \bdatw[12]_INST_0_i_1_0 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \iv[13]_i_23 ,
    \sr_reg[8]_20 ,
    \iv[12]_i_22_0 ,
    \sr_reg[8]_21 ,
    \iv[10]_i_21 ,
    \sr_reg[8]_22 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \sr_reg[8]_28 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \sr_reg[8]_33 ,
    \bdatw[12]_INST_0_i_1_1 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \bdatw[12]_INST_0_i_1_2 ,
    \sr_reg[8]_36 ,
    \sr_reg[6] ,
    \iv[10]_i_34 ,
    \iv[12]_i_34 ,
    \sr_reg[6]_0 ,
    \iv[15]_i_103 ,
    \bdatw[10]_INST_0_i_1_0 ,
    \bdatw[8]_INST_0_i_1 ,
    \badr[6]_INST_0_i_1 ,
    \badr[5]_INST_0_i_1 ,
    \badr[2]_INST_0_i_1 ,
    \badr[0]_INST_0_i_1 ,
    rst_n_fl_reg_1,
    rst_n_fl_reg_2,
    rst_n_fl_reg_3,
    rst_n_fl_reg_4,
    rst_n_fl_reg_5,
    rst_n_fl_reg_6,
    rst_n_fl_reg_7,
    rst_n_fl_reg_8,
    rst_n_fl_reg_9,
    rst_n_fl_reg_10,
    rst_n_fl_reg_11,
    rst_n_fl_reg_12,
    rst_n_fl_reg_13,
    rst_n_fl_reg_14,
    \niho_dsp_a[32]_INST_0_i_5_2 ,
    mul_b,
    dctl_sign,
    \niho_dsp_a[32]_INST_0_i_5_3 ,
    \sr_reg[6]_1 ,
    div_crdy_reg,
    div_crdy_reg_0,
    \stat_reg[2]_3 ,
    \niho_dsp_a[32]_INST_0_i_5_4 ,
    \sr_reg[4]_0 ,
    \iv[15]_i_19_1 ,
    \sr_reg[8]_37 ,
    \stat_reg[2]_4 ,
    \stat_reg[0]_3 ,
    \sr_reg[6]_2 ,
    rst_n_fl_reg_15,
    bdatw,
    \stat_reg[0]_4 ,
    rst_n_fl_reg_16,
    in0,
    ctl_sp_id4,
    rst_n_fl_reg_17,
    rst_n_fl_reg_18,
    \stat_reg[0]_5 ,
    ctl_selb_0,
    rst_n_fl_reg_19,
    rst_n_fl_reg_20,
    ccmd,
    ctl_sp_dec,
    \stat_reg[2]_5 ,
    rst_n_fl_reg_21,
    rst_n_fl_reg_22,
    rst_n_fl_reg_23,
    \stat_reg[2]_6 ,
    \stat_reg[0]_6 ,
    brdy_0,
    ctl_selb_rn,
    div_crdy_reg_1,
    \stat_reg[1] ,
    bbus_o,
    \sr_reg[6]_3 ,
    \sr_reg[8]_38 ,
    \sr_reg[8]_39 ,
    \sr_reg[8]_40 ,
    \sr_reg[8]_41 ,
    \sr_reg[8]_42 ,
    \sr_reg[6]_4 ,
    \sr_reg[8]_43 ,
    \sr_reg[8]_44 ,
    \sr_reg[8]_45 ,
    \sr_reg[8]_46 ,
    \sr_reg[8]_47 ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    \sr_reg[8]_50 ,
    \sr_reg[8]_51 ,
    \sr_reg[8]_52 ,
    rst_n_0,
    \stat_reg[2]_7 ,
    \stat_reg[0]_7 ,
    \stat_reg[2]_8 ,
    abus_sel_cr,
    \tr_reg[0] ,
    \tr_reg[1] ,
    \tr_reg[2] ,
    \tr_reg[3] ,
    \tr_reg[4] ,
    \tr_reg[5] ,
    \tr_reg[6] ,
    \tr_reg[7] ,
    \tr_reg[8] ,
    \tr_reg[9] ,
    \tr_reg[10] ,
    \tr_reg[11] ,
    \tr_reg[12] ,
    \tr_reg[13] ,
    \tr_reg[14] ,
    \tr_reg[15] ,
    \tr_reg[31] ,
    \tr_reg[30] ,
    \tr_reg[29] ,
    \tr_reg[28] ,
    \tr_reg[27] ,
    \tr_reg[26] ,
    \tr_reg[25] ,
    \tr_reg[24] ,
    \tr_reg[23] ,
    \tr_reg[22] ,
    \tr_reg[21] ,
    \tr_reg[20] ,
    \tr_reg[19] ,
    \tr_reg[18] ,
    \tr_reg[17] ,
    \tr_reg[16] ,
    E,
    \stat_reg[2]_9 ,
    \sr_reg[1]_0 ,
    \sr_reg[1]_1 ,
    \sr_reg[1]_2 ,
    \sr_reg[1]_3 ,
    \sr_reg[1]_4 ,
    \sr_reg[1]_5 ,
    \sr_reg[1]_6 ,
    \sr_reg[1]_7 ,
    \sr_reg[1]_8 ,
    \sr_reg[1]_9 ,
    \sr_reg[1]_10 ,
    \sr_reg[1]_11 ,
    \sr_reg[1]_12 ,
    \sr_reg[1]_13 ,
    \sr_reg[1]_14 ,
    \sr_reg[1]_15 ,
    \sr_reg[1]_16 ,
    \sr_reg[1]_17 ,
    \sr_reg[1]_18 ,
    \sr_reg[1]_19 ,
    \sr_reg[1]_20 ,
    \sr_reg[1]_21 ,
    \sr_reg[1]_22 ,
    \sr_reg[6]_5 ,
    \sr_reg[7] ,
    \pc_reg[15] ,
    niho_dsp_b,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    \sr_reg[8]_57 ,
    \sr_reg[8]_58 ,
    \sr_reg[8]_59 ,
    \sr_reg[8]_60 ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    \sr_reg[8]_63 ,
    \sr_reg[8]_64 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    rst_n_1,
    rst_n_2,
    brdy_1,
    badr,
    \sr_reg[8]_67 ,
    \sr_reg[8]_68 ,
    \sr_reg[8]_69 ,
    \sr_reg[8]_70 ,
    \sr_reg[8]_71 ,
    \iv[8]_i_35 ,
    S,
    \bdatw[11]_INST_0_i_2_0 ,
    \bdatw[15]_INST_0_i_1_0 ,
    \bdatw[11]_INST_0_i_1_0 ,
    \sr_reg[8]_72 ,
    abus_sel_0,
    bbus_sel_0,
    \stat_reg[0]_8 ,
    \stat_reg[2]_10 ,
    \stat_reg[0]_9 ,
    \stat_reg[2]_11 ,
    cbus_sel_0,
    fch_irq_req,
    clk,
    ctl_fetch_fl_reg_0,
    rst_n,
    \sr_reg[7]_0 ,
    \sr_reg[13] ,
    \sr_reg[4]_1 ,
    \sr_reg[4]_2 ,
    \sr_reg[5]_0 ,
    \tr_reg[4]_0 ,
    \tr_reg[4]_1 ,
    cpuid,
    \sp_reg[15] ,
    \sp_reg[30] ,
    \sp_reg[26] ,
    \sp_reg[22] ,
    \sp_reg[20] ,
    \sp_reg[18] ,
    \sp_reg[16] ,
    \sp_reg[17] ,
    \sp_reg[25] ,
    \sp_reg[24] ,
    \sp_reg[14] ,
    \sp_reg[13] ,
    \sp_reg[12] ,
    \sp_reg[11] ,
    \sp_reg[10] ,
    \sp_reg[9] ,
    \sp_reg[8] ,
    \sp_reg[7] ,
    \sp_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    O,
    \sp_reg[0] ,
    \sp_reg[4] ,
    \iv[15]_i_9_0 ,
    \sr[7]_i_4_0 ,
    mulh,
    niho_dsp_c,
    \sr_reg[4]_3 ,
    abus_0,
    \tr[23]_i_5_0 ,
    \iv[15]_i_28_0 ,
    \tr[23]_i_2 ,
    \tr[21]_i_5_0 ,
    \tr[21]_i_2 ,
    \tr[20]_i_5_0 ,
    \sr[4]_i_10_0 ,
    \tr_reg[30]_0 ,
    \tr_reg[30]_1 ,
    \tr[22]_i_5_0 ,
    \sr[4]_i_10_1 ,
    \tr_reg[26]_0 ,
    \tr[18]_i_5_0 ,
    \tr[18]_i_2_0 ,
    \tr_reg[22]_0 ,
    \tr_reg[20]_0 ,
    \tr_reg[18]_0 ,
    \tr[27]_i_5_0 ,
    \tr[24]_i_5_0 ,
    \tr_reg[17]_0 ,
    \tr[25]_i_5_0 ,
    \tr[19]_i_5_0 ,
    \tr_reg[25]_0 ,
    \tr_reg[24]_0 ,
    \tr[16]_i_7_0 ,
    \tr[27]_i_5_1 ,
    \tr[25]_i_5_1 ,
    \sr[4]_i_7_0 ,
    \iv[6]_i_2_0 ,
    \tr_reg[16]_0 ,
    \sr_reg[5]_1 ,
    \sr[4]_i_7_1 ,
    \sr[4]_i_7_2 ,
    \bdatw[5] ,
    \tr_reg[7]_0 ,
    \tr_reg[7]_1 ,
    \tr_reg[7]_2 ,
    \tr_reg[11]_0 ,
    \tr_reg[11]_1 ,
    \tr_reg[11]_2 ,
    \sr[4]_i_19 ,
    \sr[4]_i_19_0 ,
    \sr[4]_i_19_1 ,
    \tr_reg[3]_0 ,
    \tr_reg[3]_1 ,
    \tr_reg[13]_0 ,
    \tr_reg[13]_1 ,
    \tr_reg[12]_0 ,
    \sr[4]_i_5 ,
    \sr[4]_i_5_0 ,
    \tr_reg[0]_0 ,
    \tr_reg[0]_1 ,
    \tr_reg[0]_2 ,
    \tr_reg[10]_0 ,
    \tr_reg[10]_1 ,
    \tr_reg[5]_0 ,
    \tr_reg[5]_1 ,
    \tr_reg[5]_2 ,
    \tr_reg[4]_2 ,
    \tr_reg[4]_3 ,
    \tr_reg[4]_4 ,
    \sr[4]_i_5_1 ,
    \tr_reg[8]_0 ,
    \tr_reg[8]_1 ,
    \sr[4]_i_18_0 ,
    \sr[4]_i_18_1 ,
    \sr[4]_i_18_2 ,
    \tr_reg[14]_0 ,
    \tr_reg[14]_1 ,
    \sr[4]_i_18_3 ,
    \sr[4]_i_18_4 ,
    \sr[4]_i_18_5 ,
    \tr_reg[9]_0 ,
    \tr_reg[9]_1 ,
    \tr_reg[9]_2 ,
    \sr[4]_i_18_6 ,
    \sr[4]_i_18_7 ,
    \sr[4]_i_18_8 ,
    \tr_reg[6]_0 ,
    \tr_reg[15]_0 ,
    \tr_reg[15]_1 ,
    \tr_reg[15]_2 ,
    \sr[4]_i_66_0 ,
    \tr[20]_i_3 ,
    \tr[22]_i_3 ,
    \tr[21]_i_3 ,
    \tr[19]_i_9 ,
    \tr[24]_i_3 ,
    \tr[28]_i_3 ,
    \iv[7]_i_10 ,
    \sr[4]_i_91_0 ,
    \sr[4]_i_91_1 ,
    \sr[4]_i_21 ,
    \iv[6]_i_8_0 ,
    \iv[3]_i_8_0 ,
    \sr[4]_i_20 ,
    \iv[12]_i_4_0 ,
    \iv[12]_i_4_1 ,
    \iv[8]_i_2_0 ,
    \iv[8]_i_4_0 ,
    \sr[4]_i_69 ,
    \sr[4]_i_66_1 ,
    \sr[4]_i_18_9 ,
    \iv[6]_i_8_1 ,
    \tr[24]_i_7 ,
    \sr[7]_i_7 ,
    \sr[7]_i_7_0 ,
    \iv[15]_i_22 ,
    \iv[15]_i_22_0 ,
    \tr[23]_i_3 ,
    \iv[7]_i_11_0 ,
    \iv[11]_i_7_0 ,
    \sr[4]_i_43_0 ,
    \sr[4]_i_43_1 ,
    \iv[11]_i_7_1 ,
    \sr[4]_i_91_2 ,
    \iv[13]_i_2_0 ,
    \iv[12]_i_2_0 ,
    \iv[10]_i_2_0 ,
    \iv[10]_i_2_1 ,
    \sr[4]_i_39_0 ,
    \iv[8]_i_7_0 ,
    \iv[8]_i_7_1 ,
    \sr[4]_i_40_1 ,
    \iv[14]_i_7_0 ,
    \sr[4]_i_78_0 ,
    \sr[4]_i_37_0 ,
    \sr[4]_i_37_1 ,
    \iv[9]_i_7_0 ,
    \sr[4]_i_66_2 ,
    \iv[6]_i_3_0 ,
    \iv[6]_i_3_1 ,
    \iv[13]_i_5 ,
    \sr[4]_i_45 ,
    \sr[4]_i_45_0 ,
    \tr[21]_i_7 ,
    \sr[4]_i_44 ,
    \sr[4]_i_44_0 ,
    \tr[20]_i_7 ,
    \iv[14]_i_2_0 ,
    \iv[14]_i_2_1 ,
    \sr[4]_i_80 ,
    \tr[22]_i_7_0 ,
    \tr[19]_i_3 ,
    \tr[19]_i_3_0 ,
    \tr[18]_i_3 ,
    \tr[18]_i_3_0 ,
    \tr[17]_i_3 ,
    \tr[17]_i_3_0 ,
    \tr[23]_i_3_0 ,
    \iv[13]_i_6_0 ,
    \sr[4]_i_81 ,
    \iv[10]_i_5 ,
    \iv[0]_i_9 ,
    \sr[4]_i_46 ,
    \sr[4]_i_98 ,
    \iv[0]_i_21 ,
    \sr[4]_i_74_0 ,
    \sr[4]_i_74_1 ,
    \sr[4]_i_77 ,
    \iv[12]_i_6_0 ,
    \iv[13]_i_6_1 ,
    \sr[4]_i_85 ,
    \sr[4]_i_85_0 ,
    \iv[14]_i_7_1 ,
    \iv[14]_i_7_2 ,
    \tr[30]_i_8 ,
    \iv[6]_i_10_0 ,
    \sr[4]_i_78_1 ,
    \iv[10]_i_6_0 ,
    \sr[4]_i_85_1 ,
    \tr[29]_i_7 ,
    \iv[1]_i_21 ,
    \tr[28]_i_9_0 ,
    \iv[11]_i_7_2 ,
    \iv[7]_i_11_1 ,
    \iv[3]_i_21 ,
    \sr[4]_i_91_3 ,
    \iv[7]_i_10_0 ,
    \iv[6]_i_22 ,
    \sr[4]_i_24_0 ,
    \iv[3]_i_2_0 ,
    \sr[4]_i_24_1 ,
    \sr[4]_i_24_2 ,
    \sr[4]_i_7_3 ,
    \sr[4]_i_7_4 ,
    mul_rslt,
    div_crdy,
    dctl_sign_f,
    \iv[3]_i_2_1 ,
    \tr[30]_i_2_0 ,
    Q,
    \iv[7]_i_2_0 ,
    \iv[11]_i_3_0 ,
    \tr[16]_i_3_0 ,
    \tr[17]_i_2_0 ,
    \tr[18]_i_2_1 ,
    \tr[20]_i_2_0 ,
    \tr[22]_i_2_0 ,
    \tr[24]_i_2_0 ,
    \tr[25]_i_2_0 ,
    \tr[26]_i_2_0 ,
    \tr[30]_i_2_1 ,
    cbus_i,
    bdatr,
    \tr_reg[15]_3 ,
    read_cyc,
    \mul_b_reg[15] ,
    \mul_b_reg[15]_0 ,
    \mul_b_reg[14] ,
    \mul_b_reg[14]_0 ,
    \mul_b_reg[13] ,
    \mul_b_reg[13]_0 ,
    \mul_b_reg[12] ,
    \mul_b_reg[12]_0 ,
    \mul_b_reg[11] ,
    \mul_b_reg[11]_0 ,
    \mul_b_reg[10] ,
    \mul_b_reg[10]_0 ,
    \mul_b_reg[9] ,
    \mul_b_reg[9]_0 ,
    \mul_b_reg[8] ,
    \mul_b_reg[8]_0 ,
    \tr_reg[7]_3 ,
    \tr_reg[7]_4 ,
    \mul_b_reg[7] ,
    \mul_b_reg[7]_0 ,
    \tr_reg[6]_1 ,
    \tr_reg[6]_2 ,
    \mul_b_reg[6] ,
    \mul_b_reg[6]_0 ,
    \tr_reg[5]_3 ,
    \tr_reg[5]_4 ,
    \tr_reg[1]_0 ,
    \tr_reg[1]_1 ,
    \tr_reg[1]_2 ,
    \tr_reg[2]_0 ,
    \tr_reg[2]_1 ,
    \tr_reg[2]_2 ,
    \tr_reg[3]_2 ,
    \tr_reg[3]_3 ,
    \tr_reg[0]_3 ,
    \tr_reg[0]_4 ,
    \mul_b_reg[4] ,
    \mul_b_reg[4]_0 ,
    \mul_b_reg[4]_1 ,
    \mul_b_reg[3] ,
    \mul_b_reg[3]_0 ,
    \mul_b_reg[3]_1 ,
    \mul_b_reg[2] ,
    \mul_b_reg[2]_0 ,
    \mul_b_reg[2]_1 ,
    \mul_b_reg[1] ,
    \mul_b_reg[1]_0 ,
    \mul_b_reg[1]_1 ,
    \mul_b_reg[31] ,
    \mul_b_reg[31]_0 ,
    \bbus_o[30] ,
    \bbus_o[30]_0 ,
    .bbus_o_29_sp_1(bbus_o_29_sn_1),
    \bbus_o[29]_0 ,
    .bbus_o_28_sp_1(bbus_o_28_sn_1),
    \bbus_o[28]_0 ,
    .bbus_o_27_sp_1(bbus_o_27_sn_1),
    \bbus_o[27]_0 ,
    .bbus_o_26_sp_1(bbus_o_26_sn_1),
    \bbus_o[26]_0 ,
    .bbus_o_25_sp_1(bbus_o_25_sn_1),
    \bbus_o[25]_0 ,
    .bbus_o_24_sp_1(bbus_o_24_sn_1),
    \bbus_o[24]_0 ,
    .bbus_o_23_sp_1(bbus_o_23_sn_1),
    \bbus_o[23]_0 ,
    .bbus_o_22_sp_1(bbus_o_22_sn_1),
    \bbus_o[22]_0 ,
    .bbus_o_21_sp_1(bbus_o_21_sn_1),
    \bbus_o[21]_0 ,
    .bbus_o_20_sp_1(bbus_o_20_sn_1),
    \bbus_o[20]_0 ,
    .bbus_o_19_sp_1(bbus_o_19_sn_1),
    \bbus_o[19]_0 ,
    .bbus_o_18_sp_1(bbus_o_18_sn_1),
    \bbus_o[18]_0 ,
    .bbus_o_17_sp_1(bbus_o_17_sn_1),
    \bbus_o[17]_0 ,
    .bbus_o_16_sp_1(bbus_o_16_sn_1),
    \bbus_o[16]_0 ,
    ctl_fetch_fl_reg_1,
    \bcmd[3] ,
    \stat_reg[2]_12 ,
    brdy,
    \iv_reg[0] ,
    \iv[15]_i_13_0 ,
    \iv[15]_i_122_0 ,
    \ccmd[1]_INST_0_i_1_0 ,
    \iv_reg[0]_0 ,
    \stat_reg[1]_0 ,
    \ccmd[0]_INST_0_i_4_0 ,
    ctl_fetch_fl_reg_2,
    ctl_fetch_inferred_i_21_0,
    .ccmd_2_sp_1(ccmd_2_sn_1),
    \ccmd[2]_INST_0_i_2_0 ,
    \eir_fl_reg[31]_0 ,
    \iv_reg[0]_1 ,
    \stat_reg[1]_1 ,
    \stat[1]_i_10_0 ,
    \stat_reg[0]_10 ,
    ctl_fetch_inferred_i_5_0,
    ctl_fetch_inferred_i_6_0,
    \bcmd[2] ,
    irq_vec,
    \eir_fl_reg[31]_1 ,
    \stat[0]_i_2_0 ,
    \stat_reg[2]_13 ,
    \mul_b_reg[15]_1 ,
    \bcmd[0] ,
    crdy,
    \niho_dsp_a[32]_INST_0_i_9_0 ,
    \badr[31]_INST_0_i_36_0 ,
    \niho_dsp_a[32]_INST_0_i_6_0 ,
    \iv[15]_i_38_0 ,
    \tr[31]_i_12_0 ,
    \sp[0]_i_13_0 ,
    ctl_fetch_inferred_i_11_0,
    \bdatw[31]_INST_0_i_7_0 ,
    \bdatw[31]_INST_0_i_7_1 ,
    \mul_a_reg[15] ,
    ctl_fetch_inferred_i_29_0,
    irq,
    \fch_irq_lev[1]_i_2_0 ,
    \stat[1]_i_6_0 ,
    \stat_reg[0]_11 ,
    \ccmd[2]_INST_0_i_2_1 ,
    \sr[4]_i_41 ,
    \sr[4]_i_38 ,
    \sr[4]_i_46_0 ,
    \sr[4]_i_38_0 ,
    \iv[0]_i_21_0 ,
    \tr[22]_i_5_1 ,
    \tr[21]_i_5_1 ,
    \tr[20]_i_5_1 ,
    \tr[19]_i_5_1 ,
    \tr[18]_i_5_1 ,
    \tr[17]_i_5_0 ,
    \tr[16]_i_7_1 ,
    \stat_reg[2]_14 ,
    \badr[31]_INST_0_i_1 ,
    alu_sr_flag,
    fch_pc,
    rgf_pc,
    .niho_dsp_b_16_sp_1(niho_dsp_b_16_sn_1),
    .niho_dsp_b_17_sp_1(niho_dsp_b_17_sn_1),
    .niho_dsp_b_18_sp_1(niho_dsp_b_18_sn_1),
    .niho_dsp_b_19_sp_1(niho_dsp_b_19_sn_1),
    .niho_dsp_b_20_sp_1(niho_dsp_b_20_sn_1),
    .niho_dsp_b_21_sp_1(niho_dsp_b_21_sn_1),
    .niho_dsp_b_22_sp_1(niho_dsp_b_22_sn_1),
    .niho_dsp_b_23_sp_1(niho_dsp_b_23_sn_1),
    .niho_dsp_b_24_sp_1(niho_dsp_b_24_sn_1),
    .niho_dsp_b_25_sp_1(niho_dsp_b_25_sn_1),
    .niho_dsp_b_26_sp_1(niho_dsp_b_26_sn_1),
    .niho_dsp_b_27_sp_1(niho_dsp_b_27_sn_1),
    .niho_dsp_b_28_sp_1(niho_dsp_b_28_sn_1),
    .niho_dsp_b_29_sp_1(niho_dsp_b_29_sn_1),
    \niho_dsp_b[30] ,
    \niho_dsp_b[32] ,
    .niho_dsp_b_15_sp_1(niho_dsp_b_15_sn_1),
    .niho_dsp_b_1_sp_1(niho_dsp_b_1_sn_1),
    .niho_dsp_b_2_sp_1(niho_dsp_b_2_sn_1),
    .niho_dsp_b_3_sp_1(niho_dsp_b_3_sn_1),
    .niho_dsp_b_6_sp_1(niho_dsp_b_6_sn_1),
    .niho_dsp_b_7_sp_1(niho_dsp_b_7_sn_1),
    .niho_dsp_b_8_sp_1(niho_dsp_b_8_sn_1),
    .niho_dsp_b_9_sp_1(niho_dsp_b_9_sn_1),
    .niho_dsp_b_10_sp_1(niho_dsp_b_10_sn_1),
    .niho_dsp_b_11_sp_1(niho_dsp_b_11_sn_1),
    .niho_dsp_b_12_sp_1(niho_dsp_b_12_sn_1),
    .niho_dsp_b_13_sp_1(niho_dsp_b_13_sn_1),
    .niho_dsp_b_14_sp_1(niho_dsp_b_14_sn_1),
    \sr[4]_i_8_0 ,
    \iv[13]_i_8_0 ,
    \iv[4]_i_8 ,
    \iv[4]_i_8_0 ,
    \iv[1]_i_21_0 ,
    \iv[1]_i_21_1 ,
    \sr[4]_i_81_0 ,
    \sr[4]_i_81_1 ,
    \iv[5]_i_8 ,
    \iv[5]_i_8_0 ,
    irq_lev,
    p_0_in,
    fdat);
  output \sr_reg[8] ;
  output \sr_reg[4] ;
  output \sr_reg[5] ;
  output [24:0]cbus;
  output \sr_reg[11] ;
  output \stat_reg[2] ;
  output \sr_reg[10] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[1] ;
  output \sr_reg[2] ;
  output \sr_reg[3] ;
  output \sr_reg[0] ;
  output [1:0]bbus_sr;
  output [5:0]bbus_sel_cr;
  output [1:0]D;
  output [24:0]\cbus_i[30] ;
  output [2:0]\stat_reg[2]_0 ;
  output ctl_sp_inc;
  output \tr[31]_i_44_0 ;
  output \sr[6]_i_25_0 ;
  output \stat_reg[0] ;
  output \stat_reg[0]_0 ;
  output \stat_reg[0]_1 ;
  output [28:0]bbus_0;
  output \tr[29]_i_14_0 ;
  output \tr[28]_i_13_0 ;
  output rst_n_fl_reg_0;
  output \stat_reg[2]_1 ;
  output \stat_reg[0]_2 ;
  output \tr[21]_i_14_0 ;
  output \tr[23]_i_15_0 ;
  output \tr[27]_i_14 ;
  output \niho_dsp_a[15]_INST_0_i_2_0 ;
  output \tr[19]_i_14_0 ;
  output \niho_dsp_a[32]_INST_0_i_5_0 ;
  output \niho_dsp_a[32]_INST_0_i_5_1 ;
  output \stat_reg[2]_2 ;
  output \sr_reg[8]_1 ;
  output \niho_dsp_a[32]_INST_0_i_7_0 ;
  output \iv[3]_i_16 ;
  output \iv[12]_i_10 ;
  output \iv[15]_i_19_0 ;
  output \sr[4]_i_40_0 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr[7]_i_21 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \iv[0]_i_27_0 ;
  output \iv[8]_i_34_0 ;
  output \sr[7]_i_20_0 ;
  output \iv[9]_i_35 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \bdatw[12]_INST_0_i_1_0 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \iv[13]_i_23 ;
  output \sr_reg[8]_20 ;
  output \iv[12]_i_22_0 ;
  output \sr_reg[8]_21 ;
  output \iv[10]_i_21 ;
  output \sr_reg[8]_22 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \sr_reg[8]_28 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \sr_reg[8]_33 ;
  output \bdatw[12]_INST_0_i_1_1 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \bdatw[12]_INST_0_i_1_2 ;
  output \sr_reg[8]_36 ;
  output \sr_reg[6] ;
  output \iv[10]_i_34 ;
  output \iv[12]_i_34 ;
  output \sr_reg[6]_0 ;
  output \iv[15]_i_103 ;
  output \bdatw[10]_INST_0_i_1_0 ;
  output \bdatw[8]_INST_0_i_1 ;
  output \badr[6]_INST_0_i_1 ;
  output \badr[5]_INST_0_i_1 ;
  output \badr[2]_INST_0_i_1 ;
  output \badr[0]_INST_0_i_1 ;
  output rst_n_fl_reg_1;
  output rst_n_fl_reg_2;
  output rst_n_fl_reg_3;
  output rst_n_fl_reg_4;
  output rst_n_fl_reg_5;
  output rst_n_fl_reg_6;
  output rst_n_fl_reg_7;
  output rst_n_fl_reg_8;
  output rst_n_fl_reg_9;
  output rst_n_fl_reg_10;
  output rst_n_fl_reg_11;
  output rst_n_fl_reg_12;
  output rst_n_fl_reg_13;
  output rst_n_fl_reg_14;
  output \niho_dsp_a[32]_INST_0_i_5_2 ;
  output mul_b;
  output dctl_sign;
  output \niho_dsp_a[32]_INST_0_i_5_3 ;
  output \sr_reg[6]_1 ;
  output div_crdy_reg;
  output div_crdy_reg_0;
  output \stat_reg[2]_3 ;
  output \niho_dsp_a[32]_INST_0_i_5_4 ;
  output \sr_reg[4]_0 ;
  output \iv[15]_i_19_1 ;
  output \sr_reg[8]_37 ;
  output \stat_reg[2]_4 ;
  output \stat_reg[0]_3 ;
  output \sr_reg[6]_2 ;
  output rst_n_fl_reg_15;
  output [31:0]bdatw;
  output \stat_reg[0]_4 ;
  output rst_n_fl_reg_16;
  output in0;
  output ctl_sp_id4;
  output rst_n_fl_reg_17;
  output rst_n_fl_reg_18;
  output \stat_reg[0]_5 ;
  output [0:0]ctl_selb_0;
  output rst_n_fl_reg_19;
  output rst_n_fl_reg_20;
  output [3:0]ccmd;
  output ctl_sp_dec;
  output [2:0]\stat_reg[2]_5 ;
  output rst_n_fl_reg_21;
  output rst_n_fl_reg_22;
  output rst_n_fl_reg_23;
  output \stat_reg[2]_6 ;
  output \stat_reg[0]_6 ;
  output brdy_0;
  output [1:0]ctl_selb_rn;
  output div_crdy_reg_1;
  output \stat_reg[1] ;
  output [29:0]bbus_o;
  output \sr_reg[6]_3 ;
  output \sr_reg[8]_38 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[8]_40 ;
  output \sr_reg[8]_41 ;
  output \sr_reg[8]_42 ;
  output \sr_reg[6]_4 ;
  output \sr_reg[8]_43 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[8]_45 ;
  output \sr_reg[8]_46 ;
  output \sr_reg[8]_47 ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output \sr_reg[8]_50 ;
  output \sr_reg[8]_51 ;
  output \sr_reg[8]_52 ;
  output [1:0]rst_n_0;
  output \stat_reg[2]_7 ;
  output \stat_reg[0]_7 ;
  output \stat_reg[2]_8 ;
  output [3:0]abus_sel_cr;
  output \tr_reg[0] ;
  output \tr_reg[1] ;
  output \tr_reg[2] ;
  output \tr_reg[3] ;
  output \tr_reg[4] ;
  output \tr_reg[5] ;
  output \tr_reg[6] ;
  output \tr_reg[7] ;
  output \tr_reg[8] ;
  output \tr_reg[9] ;
  output \tr_reg[10] ;
  output \tr_reg[11] ;
  output \tr_reg[12] ;
  output \tr_reg[13] ;
  output \tr_reg[14] ;
  output \tr_reg[15] ;
  output \tr_reg[31] ;
  output \tr_reg[30] ;
  output \tr_reg[29] ;
  output \tr_reg[28] ;
  output \tr_reg[27] ;
  output \tr_reg[26] ;
  output \tr_reg[25] ;
  output \tr_reg[24] ;
  output \tr_reg[23] ;
  output \tr_reg[22] ;
  output \tr_reg[21] ;
  output \tr_reg[20] ;
  output \tr_reg[19] ;
  output \tr_reg[18] ;
  output \tr_reg[17] ;
  output \tr_reg[16] ;
  output [0:0]E;
  output \stat_reg[2]_9 ;
  output [0:0]\sr_reg[1]_0 ;
  output [0:0]\sr_reg[1]_1 ;
  output [0:0]\sr_reg[1]_2 ;
  output [0:0]\sr_reg[1]_3 ;
  output [0:0]\sr_reg[1]_4 ;
  output [0:0]\sr_reg[1]_5 ;
  output [0:0]\sr_reg[1]_6 ;
  output [0:0]\sr_reg[1]_7 ;
  output [0:0]\sr_reg[1]_8 ;
  output [0:0]\sr_reg[1]_9 ;
  output [0:0]\sr_reg[1]_10 ;
  output [0:0]\sr_reg[1]_11 ;
  output [0:0]\sr_reg[1]_12 ;
  output [0:0]\sr_reg[1]_13 ;
  output [0:0]\sr_reg[1]_14 ;
  output [0:0]\sr_reg[1]_15 ;
  output [0:0]\sr_reg[1]_16 ;
  output [0:0]\sr_reg[1]_17 ;
  output [0:0]\sr_reg[1]_18 ;
  output [0:0]\sr_reg[1]_19 ;
  output [0:0]\sr_reg[1]_20 ;
  output [0:0]\sr_reg[1]_21 ;
  output [0:0]\sr_reg[1]_22 ;
  output \sr_reg[6]_5 ;
  output \sr_reg[7] ;
  output [15:0]\pc_reg[15] ;
  output [29:0]niho_dsp_b;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output \sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output \sr_reg[8]_57 ;
  output \sr_reg[8]_58 ;
  output \sr_reg[8]_59 ;
  output \sr_reg[8]_60 ;
  output \sr_reg[8]_61 ;
  output \sr_reg[8]_62 ;
  output \sr_reg[8]_63 ;
  output \sr_reg[8]_64 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output rst_n_1;
  output rst_n_2;
  output brdy_1;
  output [31:0]badr;
  output \sr_reg[8]_67 ;
  output \sr_reg[8]_68 ;
  output \sr_reg[8]_69 ;
  output \sr_reg[8]_70 ;
  output \sr_reg[8]_71 ;
  output \iv[8]_i_35 ;
  output [3:0]S;
  output [3:0]\bdatw[11]_INST_0_i_2_0 ;
  output [2:0]\bdatw[15]_INST_0_i_1_0 ;
  output [2:0]\bdatw[11]_INST_0_i_1_0 ;
  output [8:0]\sr_reg[8]_72 ;
  output [7:0]abus_sel_0;
  output [7:0]bbus_sel_0;
  output \stat_reg[0]_8 ;
  output \stat_reg[2]_10 ;
  output \stat_reg[0]_9 ;
  output \stat_reg[2]_11 ;
  output [0:0]cbus_sel_0;
  input fch_irq_req;
  input clk;
  input ctl_fetch_fl_reg_0;
  input rst_n;
  input \sr_reg[7]_0 ;
  input [12:0]\sr_reg[13] ;
  input \sr_reg[4]_1 ;
  input \sr_reg[4]_2 ;
  input \sr_reg[5]_0 ;
  input \tr_reg[4]_0 ;
  input \tr_reg[4]_1 ;
  input [1:0]cpuid;
  input \sp_reg[15] ;
  input \sp_reg[30] ;
  input \sp_reg[26] ;
  input \sp_reg[22] ;
  input \sp_reg[20] ;
  input \sp_reg[18] ;
  input \sp_reg[16] ;
  input \sp_reg[17] ;
  input \sp_reg[25] ;
  input \sp_reg[24] ;
  input \sp_reg[14] ;
  input \sp_reg[13] ;
  input \sp_reg[12] ;
  input \sp_reg[11] ;
  input \sp_reg[10] ;
  input \sp_reg[9] ;
  input \sp_reg[8] ;
  input \sp_reg[7] ;
  input \sp_reg[6] ;
  input \sp_reg[5] ;
  input \sp_reg[1] ;
  input \sp_reg[2] ;
  input \sp_reg[3] ;
  input [0:0]O;
  input [0:0]\sp_reg[0] ;
  input \sp_reg[4] ;
  input [3:0]\iv[15]_i_9_0 ;
  input [0:0]\sr[7]_i_4_0 ;
  input [15:0]mulh;
  input [24:0]niho_dsp_c;
  input \sr_reg[4]_3 ;
  input [31:0]abus_0;
  input \tr[23]_i_5_0 ;
  input \iv[15]_i_28_0 ;
  input \tr[23]_i_2 ;
  input \tr[21]_i_5_0 ;
  input \tr[21]_i_2 ;
  input \tr[20]_i_5_0 ;
  input \sr[4]_i_10_0 ;
  input \tr_reg[30]_0 ;
  input \tr_reg[30]_1 ;
  input \tr[22]_i_5_0 ;
  input \sr[4]_i_10_1 ;
  input \tr_reg[26]_0 ;
  input \tr[18]_i_5_0 ;
  input \tr[18]_i_2_0 ;
  input \tr_reg[22]_0 ;
  input \tr_reg[20]_0 ;
  input \tr_reg[18]_0 ;
  input \tr[27]_i_5_0 ;
  input \tr[24]_i_5_0 ;
  input \tr_reg[17]_0 ;
  input \tr[25]_i_5_0 ;
  input \tr[19]_i_5_0 ;
  input \tr_reg[25]_0 ;
  input \tr_reg[24]_0 ;
  input \tr[16]_i_7_0 ;
  input \tr[27]_i_5_1 ;
  input \tr[25]_i_5_1 ;
  input \sr[4]_i_7_0 ;
  input \iv[6]_i_2_0 ;
  input \tr_reg[16]_0 ;
  input \sr_reg[5]_1 ;
  input \sr[4]_i_7_1 ;
  input \sr[4]_i_7_2 ;
  input [1:0]\bdatw[5] ;
  input \tr_reg[7]_0 ;
  input \tr_reg[7]_1 ;
  input \tr_reg[7]_2 ;
  input \tr_reg[11]_0 ;
  input \tr_reg[11]_1 ;
  input \tr_reg[11]_2 ;
  input \sr[4]_i_19 ;
  input \sr[4]_i_19_0 ;
  input \sr[4]_i_19_1 ;
  input \tr_reg[3]_0 ;
  input \tr_reg[3]_1 ;
  input \tr_reg[13]_0 ;
  input \tr_reg[13]_1 ;
  input \tr_reg[12]_0 ;
  input \sr[4]_i_5 ;
  input \sr[4]_i_5_0 ;
  input \tr_reg[0]_0 ;
  input \tr_reg[0]_1 ;
  input \tr_reg[0]_2 ;
  input \tr_reg[10]_0 ;
  input \tr_reg[10]_1 ;
  input \tr_reg[5]_0 ;
  input \tr_reg[5]_1 ;
  input \tr_reg[5]_2 ;
  input \tr_reg[4]_2 ;
  input \tr_reg[4]_3 ;
  input \tr_reg[4]_4 ;
  input \sr[4]_i_5_1 ;
  input \tr_reg[8]_0 ;
  input \tr_reg[8]_1 ;
  input \sr[4]_i_18_0 ;
  input \sr[4]_i_18_1 ;
  input \sr[4]_i_18_2 ;
  input \tr_reg[14]_0 ;
  input \tr_reg[14]_1 ;
  input \sr[4]_i_18_3 ;
  input \sr[4]_i_18_4 ;
  input \sr[4]_i_18_5 ;
  input \tr_reg[9]_0 ;
  input \tr_reg[9]_1 ;
  input \tr_reg[9]_2 ;
  input \sr[4]_i_18_6 ;
  input \sr[4]_i_18_7 ;
  input \sr[4]_i_18_8 ;
  input \tr_reg[6]_0 ;
  input \tr_reg[15]_0 ;
  input \tr_reg[15]_1 ;
  input \tr_reg[15]_2 ;
  input \sr[4]_i_66_0 ;
  input \tr[20]_i_3 ;
  input \tr[22]_i_3 ;
  input \tr[21]_i_3 ;
  input \tr[19]_i_9 ;
  input \tr[24]_i_3 ;
  input \tr[28]_i_3 ;
  input \iv[7]_i_10 ;
  input \sr[4]_i_91_0 ;
  input \sr[4]_i_91_1 ;
  input \sr[4]_i_21 ;
  input \iv[6]_i_8_0 ;
  input \iv[3]_i_8_0 ;
  input \sr[4]_i_20 ;
  input \iv[12]_i_4_0 ;
  input \iv[12]_i_4_1 ;
  input \iv[8]_i_2_0 ;
  input \iv[8]_i_4_0 ;
  input \sr[4]_i_69 ;
  input \sr[4]_i_66_1 ;
  input \sr[4]_i_18_9 ;
  input \iv[6]_i_8_1 ;
  input \tr[24]_i_7 ;
  input \sr[7]_i_7 ;
  input \sr[7]_i_7_0 ;
  input \iv[15]_i_22 ;
  input \iv[15]_i_22_0 ;
  input \tr[23]_i_3 ;
  input \iv[7]_i_11_0 ;
  input \iv[11]_i_7_0 ;
  input \sr[4]_i_43_0 ;
  input \sr[4]_i_43_1 ;
  input \iv[11]_i_7_1 ;
  input \sr[4]_i_91_2 ;
  input \iv[13]_i_2_0 ;
  input \iv[12]_i_2_0 ;
  input \iv[10]_i_2_0 ;
  input \iv[10]_i_2_1 ;
  input \sr[4]_i_39_0 ;
  input \iv[8]_i_7_0 ;
  input \iv[8]_i_7_1 ;
  input \sr[4]_i_40_1 ;
  input \iv[14]_i_7_0 ;
  input \sr[4]_i_78_0 ;
  input \sr[4]_i_37_0 ;
  input \sr[4]_i_37_1 ;
  input \iv[9]_i_7_0 ;
  input \sr[4]_i_66_2 ;
  input \iv[6]_i_3_0 ;
  input \iv[6]_i_3_1 ;
  input \iv[13]_i_5 ;
  input \sr[4]_i_45 ;
  input \sr[4]_i_45_0 ;
  input \tr[21]_i_7 ;
  input \sr[4]_i_44 ;
  input \sr[4]_i_44_0 ;
  input \tr[20]_i_7 ;
  input \iv[14]_i_2_0 ;
  input \iv[14]_i_2_1 ;
  input \sr[4]_i_80 ;
  input \tr[22]_i_7_0 ;
  input \tr[19]_i_3 ;
  input \tr[19]_i_3_0 ;
  input \tr[18]_i_3 ;
  input \tr[18]_i_3_0 ;
  input \tr[17]_i_3 ;
  input \tr[17]_i_3_0 ;
  input \tr[23]_i_3_0 ;
  input \iv[13]_i_6_0 ;
  input \sr[4]_i_81 ;
  input \iv[10]_i_5 ;
  input \iv[0]_i_9 ;
  input \sr[4]_i_46 ;
  input \sr[4]_i_98 ;
  input \iv[0]_i_21 ;
  input \sr[4]_i_74_0 ;
  input \sr[4]_i_74_1 ;
  input \sr[4]_i_77 ;
  input \iv[12]_i_6_0 ;
  input \iv[13]_i_6_1 ;
  input \sr[4]_i_85 ;
  input \sr[4]_i_85_0 ;
  input \iv[14]_i_7_1 ;
  input \iv[14]_i_7_2 ;
  input \tr[30]_i_8 ;
  input \iv[6]_i_10_0 ;
  input \sr[4]_i_78_1 ;
  input \iv[10]_i_6_0 ;
  input \sr[4]_i_85_1 ;
  input \tr[29]_i_7 ;
  input \iv[1]_i_21 ;
  input \tr[28]_i_9_0 ;
  input \iv[11]_i_7_2 ;
  input \iv[7]_i_11_1 ;
  input \iv[3]_i_21 ;
  input \sr[4]_i_91_3 ;
  input \iv[7]_i_10_0 ;
  input \iv[6]_i_22 ;
  input \sr[4]_i_24_0 ;
  input \iv[3]_i_2_0 ;
  input \sr[4]_i_24_1 ;
  input \sr[4]_i_24_2 ;
  input \sr[4]_i_7_3 ;
  input \sr[4]_i_7_4 ;
  input mul_rslt;
  input div_crdy;
  input dctl_sign_f;
  input [3:0]\iv[3]_i_2_1 ;
  input [24:0]\tr[30]_i_2_0 ;
  input [24:0]Q;
  input [3:0]\iv[7]_i_2_0 ;
  input [3:0]\iv[11]_i_3_0 ;
  input \tr[16]_i_3_0 ;
  input \tr[17]_i_2_0 ;
  input \tr[18]_i_2_1 ;
  input \tr[20]_i_2_0 ;
  input \tr[22]_i_2_0 ;
  input \tr[24]_i_2_0 ;
  input \tr[25]_i_2_0 ;
  input \tr[26]_i_2_0 ;
  input \tr[30]_i_2_1 ;
  input [24:0]cbus_i;
  input [16:0]bdatr;
  input \tr_reg[15]_3 ;
  input [2:0]read_cyc;
  input \mul_b_reg[15] ;
  input \mul_b_reg[15]_0 ;
  input \mul_b_reg[14] ;
  input \mul_b_reg[14]_0 ;
  input \mul_b_reg[13] ;
  input \mul_b_reg[13]_0 ;
  input \mul_b_reg[12] ;
  input \mul_b_reg[12]_0 ;
  input \mul_b_reg[11] ;
  input \mul_b_reg[11]_0 ;
  input \mul_b_reg[10] ;
  input \mul_b_reg[10]_0 ;
  input \mul_b_reg[9] ;
  input \mul_b_reg[9]_0 ;
  input \mul_b_reg[8] ;
  input \mul_b_reg[8]_0 ;
  input \tr_reg[7]_3 ;
  input \tr_reg[7]_4 ;
  input \mul_b_reg[7] ;
  input \mul_b_reg[7]_0 ;
  input \tr_reg[6]_1 ;
  input \tr_reg[6]_2 ;
  input \mul_b_reg[6] ;
  input \mul_b_reg[6]_0 ;
  input \tr_reg[5]_3 ;
  input \tr_reg[5]_4 ;
  input \tr_reg[1]_0 ;
  input \tr_reg[1]_1 ;
  input \tr_reg[1]_2 ;
  input \tr_reg[2]_0 ;
  input \tr_reg[2]_1 ;
  input \tr_reg[2]_2 ;
  input \tr_reg[3]_2 ;
  input \tr_reg[3]_3 ;
  input \tr_reg[0]_3 ;
  input \tr_reg[0]_4 ;
  input \mul_b_reg[4] ;
  input \mul_b_reg[4]_0 ;
  input \mul_b_reg[4]_1 ;
  input \mul_b_reg[3] ;
  input \mul_b_reg[3]_0 ;
  input \mul_b_reg[3]_1 ;
  input \mul_b_reg[2] ;
  input \mul_b_reg[2]_0 ;
  input \mul_b_reg[2]_1 ;
  input \mul_b_reg[1] ;
  input \mul_b_reg[1]_0 ;
  input \mul_b_reg[1]_1 ;
  input \mul_b_reg[31] ;
  input \mul_b_reg[31]_0 ;
  input \bbus_o[30] ;
  input \bbus_o[30]_0 ;
  input \bbus_o[29]_0 ;
  input \bbus_o[28]_0 ;
  input \bbus_o[27]_0 ;
  input \bbus_o[26]_0 ;
  input \bbus_o[25]_0 ;
  input \bbus_o[24]_0 ;
  input \bbus_o[23]_0 ;
  input \bbus_o[22]_0 ;
  input \bbus_o[21]_0 ;
  input \bbus_o[20]_0 ;
  input \bbus_o[19]_0 ;
  input \bbus_o[18]_0 ;
  input \bbus_o[17]_0 ;
  input \bbus_o[16]_0 ;
  input ctl_fetch_fl_reg_1;
  input \bcmd[3] ;
  input [2:0]\stat_reg[2]_12 ;
  input brdy;
  input \iv_reg[0] ;
  input \iv[15]_i_13_0 ;
  input \iv[15]_i_122_0 ;
  input \ccmd[1]_INST_0_i_1_0 ;
  input \iv_reg[0]_0 ;
  input \stat_reg[1]_0 ;
  input \ccmd[0]_INST_0_i_4_0 ;
  input ctl_fetch_fl_reg_2;
  input ctl_fetch_inferred_i_21_0;
  input \ccmd[2]_INST_0_i_2_0 ;
  input \eir_fl_reg[31]_0 ;
  input \iv_reg[0]_1 ;
  input \stat_reg[1]_1 ;
  input \stat[1]_i_10_0 ;
  input \stat_reg[0]_10 ;
  input ctl_fetch_inferred_i_5_0;
  input ctl_fetch_inferred_i_6_0;
  input \bcmd[2] ;
  input [5:0]irq_vec;
  input \eir_fl_reg[31]_1 ;
  input \stat[0]_i_2_0 ;
  input \stat_reg[2]_13 ;
  input \mul_b_reg[15]_1 ;
  input \bcmd[0] ;
  input crdy;
  input \niho_dsp_a[32]_INST_0_i_9_0 ;
  input \badr[31]_INST_0_i_36_0 ;
  input \niho_dsp_a[32]_INST_0_i_6_0 ;
  input \iv[15]_i_38_0 ;
  input \tr[31]_i_12_0 ;
  input \sp[0]_i_13_0 ;
  input ctl_fetch_inferred_i_11_0;
  input \bdatw[31]_INST_0_i_7_0 ;
  input \bdatw[31]_INST_0_i_7_1 ;
  input [15:0]\mul_a_reg[15] ;
  input ctl_fetch_inferred_i_29_0;
  input irq;
  input \fch_irq_lev[1]_i_2_0 ;
  input \stat[1]_i_6_0 ;
  input \stat_reg[0]_11 ;
  input \ccmd[2]_INST_0_i_2_1 ;
  input \sr[4]_i_41 ;
  input \sr[4]_i_38 ;
  input \sr[4]_i_46_0 ;
  input \sr[4]_i_38_0 ;
  input \iv[0]_i_21_0 ;
  input \tr[22]_i_5_1 ;
  input \tr[21]_i_5_1 ;
  input \tr[20]_i_5_1 ;
  input \tr[19]_i_5_1 ;
  input \tr[18]_i_5_1 ;
  input \tr[17]_i_5_0 ;
  input \tr[16]_i_7_1 ;
  input \stat_reg[2]_14 ;
  input [31:0]\badr[31]_INST_0_i_1 ;
  input [0:0]alu_sr_flag;
  input [15:0]fch_pc;
  input [15:0]rgf_pc;
  input \niho_dsp_b[30] ;
  input [1:0]\niho_dsp_b[32] ;
  input \sr[4]_i_8_0 ;
  input \iv[13]_i_8_0 ;
  input \iv[4]_i_8 ;
  input \iv[4]_i_8_0 ;
  input \iv[1]_i_21_0 ;
  input \iv[1]_i_21_1 ;
  input \sr[4]_i_81_0 ;
  input \sr[4]_i_81_1 ;
  input \iv[5]_i_8 ;
  input \iv[5]_i_8_0 ;
  input [1:0]irq_lev;
  input p_0_in;
  input [15:0]fdat;
     output [15:0]ir;
  input bbus_o_29_sn_1;
  input bbus_o_28_sn_1;
  input bbus_o_27_sn_1;
  input bbus_o_26_sn_1;
  input bbus_o_25_sn_1;
  input bbus_o_24_sn_1;
  input bbus_o_23_sn_1;
  input bbus_o_22_sn_1;
  input bbus_o_21_sn_1;
  input bbus_o_20_sn_1;
  input bbus_o_19_sn_1;
  input bbus_o_18_sn_1;
  input bbus_o_17_sn_1;
  input bbus_o_16_sn_1;
  input ccmd_2_sn_1;
  input niho_dsp_b_16_sn_1;
  input niho_dsp_b_17_sn_1;
  input niho_dsp_b_18_sn_1;
  input niho_dsp_b_19_sn_1;
  input niho_dsp_b_20_sn_1;
  input niho_dsp_b_21_sn_1;
  input niho_dsp_b_22_sn_1;
  input niho_dsp_b_23_sn_1;
  input niho_dsp_b_24_sn_1;
  input niho_dsp_b_25_sn_1;
  input niho_dsp_b_26_sn_1;
  input niho_dsp_b_27_sn_1;
  input niho_dsp_b_28_sn_1;
  input niho_dsp_b_29_sn_1;
  input niho_dsp_b_15_sn_1;
  input niho_dsp_b_1_sn_1;
  input niho_dsp_b_2_sn_1;
  input niho_dsp_b_3_sn_1;
  input niho_dsp_b_6_sn_1;
  input niho_dsp_b_7_sn_1;
  input niho_dsp_b_8_sn_1;
  input niho_dsp_b_9_sn_1;
  input niho_dsp_b_10_sn_1;
  input niho_dsp_b_11_sn_1;
  input niho_dsp_b_12_sn_1;
  input niho_dsp_b_13_sn_1;
  input niho_dsp_b_14_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [1:0]D;
  wire [0:0]E;
  wire [0:0]O;
  wire [24:0]Q;
  wire [3:0]S;
  wire [31:0]abus_0;
  wire [7:0]abus_sel_0;
  wire [3:0]abus_sel_cr;
  wire [4:4]acmd;
  wire [0:0]alu_sr_flag;
  wire [31:0]badr;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[15]_INST_0_i_7_n_0 ;
  wire \badr[2]_INST_0_i_1 ;
  wire [31:0]\badr[31]_INST_0_i_1 ;
  wire \badr[31]_INST_0_i_100_n_0 ;
  wire \badr[31]_INST_0_i_101_n_0 ;
  wire \badr[31]_INST_0_i_102_n_0 ;
  wire \badr[31]_INST_0_i_103_n_0 ;
  wire \badr[31]_INST_0_i_104_n_0 ;
  wire \badr[31]_INST_0_i_105_n_0 ;
  wire \badr[31]_INST_0_i_106_n_0 ;
  wire \badr[31]_INST_0_i_107_n_0 ;
  wire \badr[31]_INST_0_i_108_n_0 ;
  wire \badr[31]_INST_0_i_109_n_0 ;
  wire \badr[31]_INST_0_i_110_n_0 ;
  wire \badr[31]_INST_0_i_111_n_0 ;
  wire \badr[31]_INST_0_i_113_n_0 ;
  wire \badr[31]_INST_0_i_114_n_0 ;
  wire \badr[31]_INST_0_i_115_n_0 ;
  wire \badr[31]_INST_0_i_116_n_0 ;
  wire \badr[31]_INST_0_i_117_n_0 ;
  wire \badr[31]_INST_0_i_118_n_0 ;
  wire \badr[31]_INST_0_i_119_n_0 ;
  wire \badr[31]_INST_0_i_11_n_0 ;
  wire \badr[31]_INST_0_i_120_n_0 ;
  wire \badr[31]_INST_0_i_121_n_0 ;
  wire \badr[31]_INST_0_i_122_n_0 ;
  wire \badr[31]_INST_0_i_123_n_0 ;
  wire \badr[31]_INST_0_i_124_n_0 ;
  wire \badr[31]_INST_0_i_125_n_0 ;
  wire \badr[31]_INST_0_i_126_n_0 ;
  wire \badr[31]_INST_0_i_127_n_0 ;
  wire \badr[31]_INST_0_i_128_n_0 ;
  wire \badr[31]_INST_0_i_129_n_0 ;
  wire \badr[31]_INST_0_i_12_n_0 ;
  wire \badr[31]_INST_0_i_130_n_0 ;
  wire \badr[31]_INST_0_i_131_n_0 ;
  wire \badr[31]_INST_0_i_132_n_0 ;
  wire \badr[31]_INST_0_i_133_n_0 ;
  wire \badr[31]_INST_0_i_134_n_0 ;
  wire \badr[31]_INST_0_i_135_n_0 ;
  wire \badr[31]_INST_0_i_136_n_0 ;
  wire \badr[31]_INST_0_i_137_n_0 ;
  wire \badr[31]_INST_0_i_138_n_0 ;
  wire \badr[31]_INST_0_i_139_n_0 ;
  wire \badr[31]_INST_0_i_13_n_0 ;
  wire \badr[31]_INST_0_i_140_n_0 ;
  wire \badr[31]_INST_0_i_141_n_0 ;
  wire \badr[31]_INST_0_i_142_n_0 ;
  wire \badr[31]_INST_0_i_143_n_0 ;
  wire \badr[31]_INST_0_i_144_n_0 ;
  wire \badr[31]_INST_0_i_145_n_0 ;
  wire \badr[31]_INST_0_i_146_n_0 ;
  wire \badr[31]_INST_0_i_147_n_0 ;
  wire \badr[31]_INST_0_i_148_n_0 ;
  wire \badr[31]_INST_0_i_149_n_0 ;
  wire \badr[31]_INST_0_i_150_n_0 ;
  wire \badr[31]_INST_0_i_151_n_0 ;
  wire \badr[31]_INST_0_i_152_n_0 ;
  wire \badr[31]_INST_0_i_153_n_0 ;
  wire \badr[31]_INST_0_i_154_n_0 ;
  wire \badr[31]_INST_0_i_155_n_0 ;
  wire \badr[31]_INST_0_i_156_n_0 ;
  wire \badr[31]_INST_0_i_157_n_0 ;
  wire \badr[31]_INST_0_i_158_n_0 ;
  wire \badr[31]_INST_0_i_159_n_0 ;
  wire \badr[31]_INST_0_i_29_n_0 ;
  wire \badr[31]_INST_0_i_2_n_0 ;
  wire \badr[31]_INST_0_i_31_n_0 ;
  wire \badr[31]_INST_0_i_32_n_0 ;
  wire \badr[31]_INST_0_i_33_n_0 ;
  wire \badr[31]_INST_0_i_34_n_0 ;
  wire \badr[31]_INST_0_i_36_0 ;
  wire \badr[31]_INST_0_i_36_n_0 ;
  wire \badr[31]_INST_0_i_48_n_0 ;
  wire \badr[31]_INST_0_i_49_n_0 ;
  wire \badr[31]_INST_0_i_50_n_0 ;
  wire \badr[31]_INST_0_i_51_n_0 ;
  wire \badr[31]_INST_0_i_52_n_0 ;
  wire \badr[31]_INST_0_i_53_n_0 ;
  wire \badr[31]_INST_0_i_54_n_0 ;
  wire \badr[31]_INST_0_i_55_n_0 ;
  wire \badr[31]_INST_0_i_56_n_0 ;
  wire \badr[31]_INST_0_i_57_n_0 ;
  wire \badr[31]_INST_0_i_58_n_0 ;
  wire \badr[31]_INST_0_i_59_n_0 ;
  wire \badr[31]_INST_0_i_60_n_0 ;
  wire \badr[31]_INST_0_i_61_n_0 ;
  wire \badr[31]_INST_0_i_62_n_0 ;
  wire \badr[31]_INST_0_i_63_n_0 ;
  wire \badr[31]_INST_0_i_64_n_0 ;
  wire \badr[31]_INST_0_i_65_n_0 ;
  wire \badr[31]_INST_0_i_66_n_0 ;
  wire \badr[31]_INST_0_i_67_n_0 ;
  wire \badr[31]_INST_0_i_68_n_0 ;
  wire \badr[31]_INST_0_i_69_n_0 ;
  wire \badr[31]_INST_0_i_70_n_0 ;
  wire \badr[31]_INST_0_i_71_n_0 ;
  wire \badr[31]_INST_0_i_72_n_0 ;
  wire \badr[31]_INST_0_i_73_n_0 ;
  wire \badr[31]_INST_0_i_74_n_0 ;
  wire \badr[31]_INST_0_i_75_n_0 ;
  wire \badr[31]_INST_0_i_76_n_0 ;
  wire \badr[31]_INST_0_i_77_n_0 ;
  wire \badr[31]_INST_0_i_78_n_0 ;
  wire \badr[31]_INST_0_i_79_n_0 ;
  wire \badr[31]_INST_0_i_80_n_0 ;
  wire \badr[31]_INST_0_i_81_n_0 ;
  wire \badr[31]_INST_0_i_82_n_0 ;
  wire \badr[31]_INST_0_i_83_n_0 ;
  wire \badr[31]_INST_0_i_84_n_0 ;
  wire \badr[31]_INST_0_i_85_n_0 ;
  wire \badr[31]_INST_0_i_86_n_0 ;
  wire \badr[31]_INST_0_i_87_n_0 ;
  wire \badr[31]_INST_0_i_88_n_0 ;
  wire \badr[31]_INST_0_i_89_n_0 ;
  wire \badr[31]_INST_0_i_90_n_0 ;
  wire \badr[31]_INST_0_i_91_n_0 ;
  wire \badr[31]_INST_0_i_92_n_0 ;
  wire \badr[31]_INST_0_i_93_n_0 ;
  wire \badr[31]_INST_0_i_94_n_0 ;
  wire \badr[31]_INST_0_i_95_n_0 ;
  wire \badr[31]_INST_0_i_96_n_0 ;
  wire \badr[31]_INST_0_i_97_n_0 ;
  wire \badr[31]_INST_0_i_98_n_0 ;
  wire \badr[31]_INST_0_i_99_n_0 ;
  wire \badr[31]_INST_0_i_9_n_0 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1 ;
  wire [28:0]bbus_0;
  wire [29:0]bbus_o;
  wire \bbus_o[16]_0 ;
  wire \bbus_o[17]_0 ;
  wire \bbus_o[18]_0 ;
  wire \bbus_o[19]_0 ;
  wire \bbus_o[20]_0 ;
  wire \bbus_o[21]_0 ;
  wire \bbus_o[22]_0 ;
  wire \bbus_o[23]_0 ;
  wire \bbus_o[24]_0 ;
  wire \bbus_o[25]_0 ;
  wire \bbus_o[26]_0 ;
  wire \bbus_o[27]_0 ;
  wire \bbus_o[28]_0 ;
  wire \bbus_o[29]_0 ;
  wire \bbus_o[30] ;
  wire \bbus_o[30]_0 ;
  wire bbus_o_16_sn_1;
  wire bbus_o_17_sn_1;
  wire bbus_o_18_sn_1;
  wire bbus_o_19_sn_1;
  wire bbus_o_20_sn_1;
  wire bbus_o_21_sn_1;
  wire bbus_o_22_sn_1;
  wire bbus_o_23_sn_1;
  wire bbus_o_24_sn_1;
  wire bbus_o_25_sn_1;
  wire bbus_o_26_sn_1;
  wire bbus_o_27_sn_1;
  wire bbus_o_28_sn_1;
  wire bbus_o_29_sn_1;
  wire [7:0]bbus_sel_0;
  wire [5:0]bbus_sel_cr;
  wire [1:0]bbus_sr;
  wire \bcmd[0] ;
  wire \bcmd[0]_INST_0_i_11_n_0 ;
  wire \bcmd[0]_INST_0_i_12_n_0 ;
  wire \bcmd[0]_INST_0_i_1_n_0 ;
  wire \bcmd[0]_INST_0_i_2_n_0 ;
  wire \bcmd[0]_INST_0_i_3_n_0 ;
  wire \bcmd[0]_INST_0_i_4_n_0 ;
  wire \bcmd[0]_INST_0_i_5_n_0 ;
  wire \bcmd[0]_INST_0_i_6_n_0 ;
  wire \bcmd[0]_INST_0_i_7_n_0 ;
  wire \bcmd[0]_INST_0_i_8_n_0 ;
  wire \bcmd[0]_INST_0_i_9_n_0 ;
  wire \bcmd[1]_INST_0_i_10_n_0 ;
  wire \bcmd[1]_INST_0_i_11_n_0 ;
  wire \bcmd[1]_INST_0_i_12_n_0 ;
  wire \bcmd[1]_INST_0_i_13_n_0 ;
  wire \bcmd[1]_INST_0_i_15_n_0 ;
  wire \bcmd[1]_INST_0_i_16_n_0 ;
  wire \bcmd[1]_INST_0_i_1_n_0 ;
  wire \bcmd[1]_INST_0_i_2_n_0 ;
  wire \bcmd[1]_INST_0_i_3_n_0 ;
  wire \bcmd[1]_INST_0_i_4_n_0 ;
  wire \bcmd[1]_INST_0_i_5_n_0 ;
  wire \bcmd[1]_INST_0_i_7_n_0 ;
  wire \bcmd[1]_INST_0_i_8_n_0 ;
  wire \bcmd[1]_INST_0_i_9_n_0 ;
  wire \bcmd[2] ;
  wire \bcmd[3] ;
  wire \bcmd[3]_INST_0_i_10_n_0 ;
  wire \bcmd[3]_INST_0_i_11_n_0 ;
  wire \bcmd[3]_INST_0_i_12_n_0 ;
  wire \bcmd[3]_INST_0_i_13_n_0 ;
  wire \bcmd[3]_INST_0_i_14_n_0 ;
  wire \bcmd[3]_INST_0_i_15_n_0 ;
  wire \bcmd[3]_INST_0_i_16_n_0 ;
  wire \bcmd[3]_INST_0_i_1_n_0 ;
  wire \bcmd[3]_INST_0_i_2_n_0 ;
  wire \bcmd[3]_INST_0_i_4_n_0 ;
  wire \bcmd[3]_INST_0_i_5_n_0 ;
  wire \bcmd[3]_INST_0_i_6_n_0 ;
  wire \bcmd[3]_INST_0_i_8_n_0 ;
  wire \bcmd[3]_INST_0_i_9_n_0 ;
  wire [16:0]bdatr;
  wire [31:0]bdatw;
  wire \bdatw[10]_INST_0_i_10_n_0 ;
  wire \bdatw[10]_INST_0_i_1_0 ;
  wire \bdatw[10]_INST_0_i_3_n_0 ;
  wire \bdatw[10]_INST_0_i_7_n_0 ;
  wire \bdatw[11]_INST_0_i_19_n_0 ;
  wire [2:0]\bdatw[11]_INST_0_i_1_0 ;
  wire [3:0]\bdatw[11]_INST_0_i_2_0 ;
  wire \bdatw[11]_INST_0_i_6_n_0 ;
  wire \bdatw[11]_INST_0_i_7_n_0 ;
  wire \bdatw[12]_INST_0_i_1_0 ;
  wire \bdatw[12]_INST_0_i_1_1 ;
  wire \bdatw[12]_INST_0_i_1_2 ;
  wire \bdatw[12]_INST_0_i_22_n_0 ;
  wire \bdatw[12]_INST_0_i_23_n_0 ;
  wire \bdatw[12]_INST_0_i_3_n_0 ;
  wire \bdatw[12]_INST_0_i_4_n_0 ;
  wire \bdatw[12]_INST_0_i_9_n_0 ;
  wire \bdatw[13]_INST_0_i_12_n_0 ;
  wire \bdatw[13]_INST_0_i_27_n_0 ;
  wire \bdatw[13]_INST_0_i_9_n_0 ;
  wire \bdatw[14]_INST_0_i_3_n_0 ;
  wire \bdatw[14]_INST_0_i_6_n_0 ;
  wire \bdatw[14]_INST_0_i_9_n_0 ;
  wire \bdatw[15]_INST_0_i_10_n_0 ;
  wire \bdatw[15]_INST_0_i_11_n_0 ;
  wire \bdatw[15]_INST_0_i_12_n_0 ;
  wire \bdatw[15]_INST_0_i_13_n_0 ;
  wire \bdatw[15]_INST_0_i_14_n_0 ;
  wire [2:0]\bdatw[15]_INST_0_i_1_0 ;
  wire \bdatw[15]_INST_0_i_28_n_0 ;
  wire \bdatw[15]_INST_0_i_29_n_0 ;
  wire \bdatw[15]_INST_0_i_3_n_0 ;
  wire \bdatw[15]_INST_0_i_70_n_0 ;
  wire \bdatw[15]_INST_0_i_71_n_0 ;
  wire \bdatw[15]_INST_0_i_72_n_0 ;
  wire \bdatw[15]_INST_0_i_73_n_0 ;
  wire \bdatw[15]_INST_0_i_74_n_0 ;
  wire \bdatw[15]_INST_0_i_75_n_0 ;
  wire \bdatw[15]_INST_0_i_76_n_0 ;
  wire \bdatw[15]_INST_0_i_77_n_0 ;
  wire \bdatw[15]_INST_0_i_78_n_0 ;
  wire \bdatw[15]_INST_0_i_79_n_0 ;
  wire \bdatw[15]_INST_0_i_7_n_0 ;
  wire \bdatw[31]_INST_0_i_100_n_0 ;
  wire \bdatw[31]_INST_0_i_101_n_0 ;
  wire \bdatw[31]_INST_0_i_102_n_0 ;
  wire \bdatw[31]_INST_0_i_103_n_0 ;
  wire \bdatw[31]_INST_0_i_18_n_0 ;
  wire \bdatw[31]_INST_0_i_19_n_0 ;
  wire \bdatw[31]_INST_0_i_20_n_0 ;
  wire \bdatw[31]_INST_0_i_21_n_0 ;
  wire \bdatw[31]_INST_0_i_22_n_0 ;
  wire \bdatw[31]_INST_0_i_23_n_0 ;
  wire \bdatw[31]_INST_0_i_24_n_0 ;
  wire \bdatw[31]_INST_0_i_25_n_0 ;
  wire \bdatw[31]_INST_0_i_26_n_0 ;
  wire \bdatw[31]_INST_0_i_27_n_0 ;
  wire \bdatw[31]_INST_0_i_28_n_0 ;
  wire \bdatw[31]_INST_0_i_2_n_0 ;
  wire \bdatw[31]_INST_0_i_3_n_0 ;
  wire \bdatw[31]_INST_0_i_46_n_0 ;
  wire \bdatw[31]_INST_0_i_47_n_0 ;
  wire \bdatw[31]_INST_0_i_48_n_0 ;
  wire \bdatw[31]_INST_0_i_49_n_0 ;
  wire \bdatw[31]_INST_0_i_50_n_0 ;
  wire \bdatw[31]_INST_0_i_51_n_0 ;
  wire \bdatw[31]_INST_0_i_52_n_0 ;
  wire \bdatw[31]_INST_0_i_53_n_0 ;
  wire \bdatw[31]_INST_0_i_54_n_0 ;
  wire \bdatw[31]_INST_0_i_55_n_0 ;
  wire \bdatw[31]_INST_0_i_56_n_0 ;
  wire \bdatw[31]_INST_0_i_57_n_0 ;
  wire \bdatw[31]_INST_0_i_58_n_0 ;
  wire \bdatw[31]_INST_0_i_59_n_0 ;
  wire \bdatw[31]_INST_0_i_60_n_0 ;
  wire \bdatw[31]_INST_0_i_63_n_0 ;
  wire \bdatw[31]_INST_0_i_64_n_0 ;
  wire \bdatw[31]_INST_0_i_65_n_0 ;
  wire \bdatw[31]_INST_0_i_66_n_0 ;
  wire \bdatw[31]_INST_0_i_67_n_0 ;
  wire \bdatw[31]_INST_0_i_68_n_0 ;
  wire \bdatw[31]_INST_0_i_69_n_0 ;
  wire \bdatw[31]_INST_0_i_70_n_0 ;
  wire \bdatw[31]_INST_0_i_71_n_0 ;
  wire \bdatw[31]_INST_0_i_72_n_0 ;
  wire \bdatw[31]_INST_0_i_73_n_0 ;
  wire \bdatw[31]_INST_0_i_74_n_0 ;
  wire \bdatw[31]_INST_0_i_75_n_0 ;
  wire \bdatw[31]_INST_0_i_76_n_0 ;
  wire \bdatw[31]_INST_0_i_77_n_0 ;
  wire \bdatw[31]_INST_0_i_78_n_0 ;
  wire \bdatw[31]_INST_0_i_79_n_0 ;
  wire \bdatw[31]_INST_0_i_7_0 ;
  wire \bdatw[31]_INST_0_i_7_1 ;
  wire \bdatw[31]_INST_0_i_80_n_0 ;
  wire \bdatw[31]_INST_0_i_81_n_0 ;
  wire \bdatw[31]_INST_0_i_82_n_0 ;
  wire \bdatw[31]_INST_0_i_83_n_0 ;
  wire \bdatw[31]_INST_0_i_84_n_0 ;
  wire \bdatw[31]_INST_0_i_85_n_0 ;
  wire \bdatw[31]_INST_0_i_86_n_0 ;
  wire \bdatw[31]_INST_0_i_87_n_0 ;
  wire \bdatw[31]_INST_0_i_88_n_0 ;
  wire \bdatw[31]_INST_0_i_89_n_0 ;
  wire \bdatw[31]_INST_0_i_8_n_0 ;
  wire \bdatw[31]_INST_0_i_90_n_0 ;
  wire \bdatw[31]_INST_0_i_91_n_0 ;
  wire \bdatw[31]_INST_0_i_92_n_0 ;
  wire \bdatw[31]_INST_0_i_93_n_0 ;
  wire \bdatw[31]_INST_0_i_94_n_0 ;
  wire \bdatw[31]_INST_0_i_95_n_0 ;
  wire \bdatw[31]_INST_0_i_96_n_0 ;
  wire \bdatw[31]_INST_0_i_97_n_0 ;
  wire \bdatw[31]_INST_0_i_98_n_0 ;
  wire \bdatw[31]_INST_0_i_99_n_0 ;
  wire [1:0]\bdatw[5] ;
  wire \bdatw[8]_INST_0_i_1 ;
  wire \bdatw[8]_INST_0_i_9_n_0 ;
  wire \bdatw[9]_INST_0_i_10_n_0 ;
  wire \bdatw[9]_INST_0_i_20_n_0 ;
  wire \bdatw[9]_INST_0_i_3_n_0 ;
  wire \bdatw[9]_INST_0_i_7_n_0 ;
  wire brdy;
  wire brdy_0;
  wire brdy_1;
  wire [24:0]cbus;
  wire [24:0]cbus_i;
  wire [24:0]\cbus_i[30] ;
  wire [0:0]cbus_sel_0;
  wire [3:0]ccmd;
  wire \ccmd[0]_INST_0_i_10_n_0 ;
  wire \ccmd[0]_INST_0_i_11_n_0 ;
  wire \ccmd[0]_INST_0_i_12_n_0 ;
  wire \ccmd[0]_INST_0_i_13_n_0 ;
  wire \ccmd[0]_INST_0_i_15_n_0 ;
  wire \ccmd[0]_INST_0_i_17_n_0 ;
  wire \ccmd[0]_INST_0_i_18_n_0 ;
  wire \ccmd[0]_INST_0_i_19_n_0 ;
  wire \ccmd[0]_INST_0_i_1_n_0 ;
  wire \ccmd[0]_INST_0_i_20_n_0 ;
  wire \ccmd[0]_INST_0_i_21_n_0 ;
  wire \ccmd[0]_INST_0_i_22_n_0 ;
  wire \ccmd[0]_INST_0_i_2_n_0 ;
  wire \ccmd[0]_INST_0_i_3_n_0 ;
  wire \ccmd[0]_INST_0_i_4_0 ;
  wire \ccmd[0]_INST_0_i_4_n_0 ;
  wire \ccmd[0]_INST_0_i_5_n_0 ;
  wire \ccmd[0]_INST_0_i_7_n_0 ;
  wire \ccmd[0]_INST_0_i_8_n_0 ;
  wire \ccmd[0]_INST_0_i_9_n_0 ;
  wire \ccmd[1]_INST_0_i_11_n_0 ;
  wire \ccmd[1]_INST_0_i_13_n_0 ;
  wire \ccmd[1]_INST_0_i_14_n_0 ;
  wire \ccmd[1]_INST_0_i_15_n_0 ;
  wire \ccmd[1]_INST_0_i_16_n_0 ;
  wire \ccmd[1]_INST_0_i_17_n_0 ;
  wire \ccmd[1]_INST_0_i_18_n_0 ;
  wire \ccmd[1]_INST_0_i_1_0 ;
  wire \ccmd[1]_INST_0_i_1_n_0 ;
  wire \ccmd[1]_INST_0_i_2_n_0 ;
  wire \ccmd[1]_INST_0_i_3_n_0 ;
  wire \ccmd[1]_INST_0_i_4_n_0 ;
  wire \ccmd[1]_INST_0_i_5_n_0 ;
  wire \ccmd[1]_INST_0_i_6_n_0 ;
  wire \ccmd[1]_INST_0_i_7_n_0 ;
  wire \ccmd[1]_INST_0_i_8_n_0 ;
  wire \ccmd[1]_INST_0_i_9_n_0 ;
  wire \ccmd[2]_INST_0_i_10_n_0 ;
  wire \ccmd[2]_INST_0_i_11_n_0 ;
  wire \ccmd[2]_INST_0_i_12_n_0 ;
  wire \ccmd[2]_INST_0_i_15_n_0 ;
  wire \ccmd[2]_INST_0_i_16_n_0 ;
  wire \ccmd[2]_INST_0_i_17_n_0 ;
  wire \ccmd[2]_INST_0_i_1_n_0 ;
  wire \ccmd[2]_INST_0_i_2_0 ;
  wire \ccmd[2]_INST_0_i_2_1 ;
  wire \ccmd[2]_INST_0_i_2_n_0 ;
  wire \ccmd[2]_INST_0_i_4_n_0 ;
  wire \ccmd[2]_INST_0_i_5_n_0 ;
  wire \ccmd[2]_INST_0_i_6_n_0 ;
  wire \ccmd[2]_INST_0_i_7_n_0 ;
  wire \ccmd[2]_INST_0_i_8_n_0 ;
  wire \ccmd[2]_INST_0_i_9_n_0 ;
  wire \ccmd[3]_INST_0_i_10_n_0 ;
  wire \ccmd[3]_INST_0_i_11_n_0 ;
  wire \ccmd[3]_INST_0_i_12_n_0 ;
  wire \ccmd[3]_INST_0_i_13_n_0 ;
  wire \ccmd[3]_INST_0_i_15_n_0 ;
  wire \ccmd[3]_INST_0_i_16_n_0 ;
  wire \ccmd[3]_INST_0_i_17_n_0 ;
  wire \ccmd[3]_INST_0_i_18_n_0 ;
  wire \ccmd[3]_INST_0_i_19_n_0 ;
  wire \ccmd[3]_INST_0_i_1_n_0 ;
  wire \ccmd[3]_INST_0_i_20_n_0 ;
  wire \ccmd[3]_INST_0_i_21_n_0 ;
  wire \ccmd[3]_INST_0_i_22_n_0 ;
  wire \ccmd[3]_INST_0_i_23_n_0 ;
  wire \ccmd[3]_INST_0_i_24_n_0 ;
  wire \ccmd[3]_INST_0_i_25_n_0 ;
  wire \ccmd[3]_INST_0_i_2_n_0 ;
  wire \ccmd[3]_INST_0_i_3_n_0 ;
  wire \ccmd[3]_INST_0_i_4_n_0 ;
  wire \ccmd[3]_INST_0_i_5_n_0 ;
  wire \ccmd[3]_INST_0_i_6_n_0 ;
  wire \ccmd[3]_INST_0_i_7_n_0 ;
  wire \ccmd[3]_INST_0_i_8_n_0 ;
  wire \ccmd[3]_INST_0_i_9_n_0 ;
  wire \ccmd[4]_INST_0_i_1_n_0 ;
  wire \ccmd[4]_INST_0_i_2_n_0 ;
  wire \ccmd[4]_INST_0_i_3_n_0 ;
  wire \ccmd[4]_INST_0_i_4_n_0 ;
  wire ccmd_2_sn_1;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  wire ctl_fetch_ext;
  wire ctl_fetch_ext_fl;
  wire ctl_fetch_ext_fl_i_2_n_0;
  wire ctl_fetch_ext_fl_i_3_n_0;
  wire ctl_fetch_ext_fl_i_4_n_0;
  wire ctl_fetch_ext_fl_i_5_n_0;
  wire ctl_fetch_fl;
  wire ctl_fetch_fl_reg_0;
  wire ctl_fetch_fl_reg_1;
  wire ctl_fetch_fl_reg_2;
  wire ctl_fetch_inferred_i_11_0;
  wire ctl_fetch_inferred_i_11_n_0;
  wire ctl_fetch_inferred_i_12_n_0;
  wire ctl_fetch_inferred_i_13_n_0;
  wire ctl_fetch_inferred_i_14_n_0;
  wire ctl_fetch_inferred_i_15_n_0;
  wire ctl_fetch_inferred_i_16_n_0;
  wire ctl_fetch_inferred_i_17_n_0;
  wire ctl_fetch_inferred_i_18_n_0;
  wire ctl_fetch_inferred_i_19_n_0;
  wire ctl_fetch_inferred_i_20_n_0;
  wire ctl_fetch_inferred_i_21_0;
  wire ctl_fetch_inferred_i_21_n_0;
  wire ctl_fetch_inferred_i_22_n_0;
  wire ctl_fetch_inferred_i_23_n_0;
  wire ctl_fetch_inferred_i_24_n_0;
  wire ctl_fetch_inferred_i_26_n_0;
  wire ctl_fetch_inferred_i_27_n_0;
  wire ctl_fetch_inferred_i_28_n_0;
  wire ctl_fetch_inferred_i_29_0;
  wire ctl_fetch_inferred_i_29_n_0;
  wire ctl_fetch_inferred_i_2_n_0;
  wire ctl_fetch_inferred_i_31_n_0;
  wire ctl_fetch_inferred_i_32_n_0;
  wire ctl_fetch_inferred_i_33_n_0;
  wire ctl_fetch_inferred_i_34_n_0;
  wire ctl_fetch_inferred_i_35_n_0;
  wire ctl_fetch_inferred_i_36_n_0;
  wire ctl_fetch_inferred_i_37_n_0;
  wire ctl_fetch_inferred_i_38_n_0;
  wire ctl_fetch_inferred_i_39_n_0;
  wire ctl_fetch_inferred_i_41_n_0;
  wire ctl_fetch_inferred_i_42_n_0;
  wire ctl_fetch_inferred_i_44_n_0;
  wire ctl_fetch_inferred_i_45_n_0;
  wire ctl_fetch_inferred_i_46_n_0;
  wire ctl_fetch_inferred_i_47_n_0;
  wire ctl_fetch_inferred_i_48_n_0;
  wire ctl_fetch_inferred_i_49_n_0;
  wire ctl_fetch_inferred_i_4_n_0;
  wire ctl_fetch_inferred_i_51_n_0;
  wire ctl_fetch_inferred_i_53_n_0;
  wire ctl_fetch_inferred_i_5_0;
  wire ctl_fetch_inferred_i_5_n_0;
  wire ctl_fetch_inferred_i_6_0;
  wire ctl_fetch_inferred_i_6_n_0;
  wire ctl_fetch_inferred_i_7_n_0;
  wire ctl_fetch_inferred_i_8_n_0;
  wire [0:0]ctl_sela;
  wire [0:0]ctl_sela_rn;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire [1:0]ctl_selc;
  wire [1:0]ctl_selc_rn;
  wire ctl_sp_dec;
  wire ctl_sp_id4;
  wire ctl_sp_inc;
  wire ctl_sr_ldie;
  wire ctl_sr_upd;
  wire dctl_sign;
  wire dctl_sign_f;
  wire div_crdy;
  wire div_crdy_reg;
  wire div_crdy_reg_0;
  wire div_crdy_reg_1;
  (* DONT_TOUCH *) wire [31:0]eir;
  wire eir_fl0;
  wire \eir_fl[1]_i_1_n_0 ;
  wire \eir_fl[2]_i_1_n_0 ;
  wire \eir_fl[31]_i_1_n_0 ;
  wire \eir_fl[31]_i_2_n_0 ;
  wire \eir_fl[31]_i_4_n_0 ;
  wire \eir_fl[31]_i_5_n_0 ;
  wire \eir_fl[3]_i_1_n_0 ;
  wire \eir_fl[4]_i_1_n_0 ;
  wire \eir_fl[5]_i_1_n_0 ;
  wire \eir_fl[6]_i_2_n_0 ;
  wire \eir_fl_reg[31]_0 ;
  wire \eir_fl_reg[31]_1 ;
  wire \eir_fl_reg_n_0_[0] ;
  wire \eir_fl_reg_n_0_[10] ;
  wire \eir_fl_reg_n_0_[11] ;
  wire \eir_fl_reg_n_0_[12] ;
  wire \eir_fl_reg_n_0_[13] ;
  wire \eir_fl_reg_n_0_[14] ;
  wire \eir_fl_reg_n_0_[15] ;
  wire \eir_fl_reg_n_0_[16] ;
  wire \eir_fl_reg_n_0_[17] ;
  wire \eir_fl_reg_n_0_[18] ;
  wire \eir_fl_reg_n_0_[19] ;
  wire \eir_fl_reg_n_0_[1] ;
  wire \eir_fl_reg_n_0_[20] ;
  wire \eir_fl_reg_n_0_[21] ;
  wire \eir_fl_reg_n_0_[22] ;
  wire \eir_fl_reg_n_0_[23] ;
  wire \eir_fl_reg_n_0_[24] ;
  wire \eir_fl_reg_n_0_[25] ;
  wire \eir_fl_reg_n_0_[26] ;
  wire \eir_fl_reg_n_0_[27] ;
  wire \eir_fl_reg_n_0_[28] ;
  wire \eir_fl_reg_n_0_[29] ;
  wire \eir_fl_reg_n_0_[2] ;
  wire \eir_fl_reg_n_0_[30] ;
  wire \eir_fl_reg_n_0_[31] ;
  wire \eir_fl_reg_n_0_[3] ;
  wire \eir_fl_reg_n_0_[4] ;
  wire \eir_fl_reg_n_0_[5] ;
  wire \eir_fl_reg_n_0_[6] ;
  wire \eir_fl_reg_n_0_[7] ;
  wire \eir_fl_reg_n_0_[8] ;
  wire \eir_fl_reg_n_0_[9] ;
  wire [1:0]fch_irq_lev;
  wire fch_irq_lev0;
  wire \fch_irq_lev[0]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_1_n_0 ;
  wire \fch_irq_lev[1]_i_2_0 ;
  wire \fch_irq_lev[1]_i_3_n_0 ;
  wire \fch_irq_lev[1]_i_4_n_0 ;
  wire \fch_irq_lev[1]_i_5_n_0 ;
  wire fch_irq_req;
  wire fch_irq_req_fl;
  wire [15:0]fch_pc;
  wire [15:0]fdat;
  wire \grn[15]_i_2__0_n_0 ;
  wire \grn[15]_i_2__2_n_0 ;
  wire in0;
  (* DONT_TOUCH *) wire [15:0]ir;
  wire [15:0]ir_fl;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire \iv[0]_i_13_n_0 ;
  wire \iv[0]_i_21 ;
  wire \iv[0]_i_21_0 ;
  wire \iv[0]_i_27_0 ;
  wire \iv[0]_i_2_n_0 ;
  wire \iv[0]_i_3_n_0 ;
  wire \iv[0]_i_6_n_0 ;
  wire \iv[0]_i_7_n_0 ;
  wire \iv[0]_i_9 ;
  wire \iv[10]_i_15_n_0 ;
  wire \iv[10]_i_17_n_0 ;
  wire \iv[10]_i_18_n_0 ;
  wire \iv[10]_i_19_n_0 ;
  wire \iv[10]_i_20_n_0 ;
  wire \iv[10]_i_21 ;
  wire \iv[10]_i_2_0 ;
  wire \iv[10]_i_2_1 ;
  wire \iv[10]_i_2_n_0 ;
  wire \iv[10]_i_34 ;
  wire \iv[10]_i_37_n_0 ;
  wire \iv[10]_i_3_n_0 ;
  wire \iv[10]_i_5 ;
  wire \iv[10]_i_6_0 ;
  wire \iv[10]_i_6_n_0 ;
  wire \iv[10]_i_7_n_0 ;
  wire \iv[10]_i_8_n_0 ;
  wire \iv[11]_i_17_n_0 ;
  wire \iv[11]_i_18_n_0 ;
  wire \iv[11]_i_19_n_0 ;
  wire \iv[11]_i_20_n_0 ;
  wire \iv[11]_i_21_n_0 ;
  wire \iv[11]_i_2_n_0 ;
  wire \iv[11]_i_39_n_0 ;
  wire [3:0]\iv[11]_i_3_0 ;
  wire \iv[11]_i_3_n_0 ;
  wire \iv[11]_i_40_n_0 ;
  wire \iv[11]_i_7_0 ;
  wire \iv[11]_i_7_1 ;
  wire \iv[11]_i_7_2 ;
  wire \iv[11]_i_7_n_0 ;
  wire \iv[11]_i_8_n_0 ;
  wire \iv[11]_i_9_n_0 ;
  wire \iv[12]_i_10 ;
  wire \iv[12]_i_15_n_0 ;
  wire \iv[12]_i_17_n_0 ;
  wire \iv[12]_i_18_n_0 ;
  wire \iv[12]_i_19_n_0 ;
  wire \iv[12]_i_20_n_0 ;
  wire \iv[12]_i_22_0 ;
  wire \iv[12]_i_26_n_0 ;
  wire \iv[12]_i_2_0 ;
  wire \iv[12]_i_2_n_0 ;
  wire \iv[12]_i_34 ;
  wire \iv[12]_i_37_n_0 ;
  wire \iv[12]_i_3_n_0 ;
  wire \iv[12]_i_4_0 ;
  wire \iv[12]_i_4_1 ;
  wire \iv[12]_i_6_0 ;
  wire \iv[12]_i_6_n_0 ;
  wire \iv[12]_i_7_n_0 ;
  wire \iv[12]_i_8_n_0 ;
  wire \iv[12]_i_9_n_0 ;
  wire \iv[13]_i_15_n_0 ;
  wire \iv[13]_i_17_n_0 ;
  wire \iv[13]_i_18_n_0 ;
  wire \iv[13]_i_19_n_0 ;
  wire \iv[13]_i_20_n_0 ;
  wire \iv[13]_i_23 ;
  wire \iv[13]_i_28_n_0 ;
  wire \iv[13]_i_2_0 ;
  wire \iv[13]_i_2_n_0 ;
  wire \iv[13]_i_3_n_0 ;
  wire \iv[13]_i_5 ;
  wire \iv[13]_i_6_0 ;
  wire \iv[13]_i_6_1 ;
  wire \iv[13]_i_6_n_0 ;
  wire \iv[13]_i_7_n_0 ;
  wire \iv[13]_i_8_0 ;
  wire \iv[13]_i_8_n_0 ;
  wire \iv[14]_i_17_n_0 ;
  wire \iv[14]_i_18_n_0 ;
  wire \iv[14]_i_19_n_0 ;
  wire \iv[14]_i_20_n_0 ;
  wire \iv[14]_i_21_n_0 ;
  wire \iv[14]_i_22_n_0 ;
  wire \iv[14]_i_28_n_0 ;
  wire \iv[14]_i_2_0 ;
  wire \iv[14]_i_2_1 ;
  wire \iv[14]_i_2_n_0 ;
  wire \iv[14]_i_3_n_0 ;
  wire \iv[14]_i_40_n_0 ;
  wire \iv[14]_i_41_n_0 ;
  wire \iv[14]_i_6_n_0 ;
  wire \iv[14]_i_7_0 ;
  wire \iv[14]_i_7_1 ;
  wire \iv[14]_i_7_2 ;
  wire \iv[14]_i_7_n_0 ;
  wire \iv[14]_i_8_n_0 ;
  wire \iv[14]_i_9_n_0 ;
  wire \iv[15]_i_100_n_0 ;
  wire \iv[15]_i_103 ;
  wire \iv[15]_i_107_n_0 ;
  wire \iv[15]_i_109_n_0 ;
  wire \iv[15]_i_10_n_0 ;
  wire \iv[15]_i_111_n_0 ;
  wire \iv[15]_i_112_n_0 ;
  wire \iv[15]_i_113_n_0 ;
  wire \iv[15]_i_114_n_0 ;
  wire \iv[15]_i_115_n_0 ;
  wire \iv[15]_i_116_n_0 ;
  wire \iv[15]_i_117_n_0 ;
  wire \iv[15]_i_118_n_0 ;
  wire \iv[15]_i_11_n_0 ;
  wire \iv[15]_i_120_n_0 ;
  wire \iv[15]_i_121_n_0 ;
  wire \iv[15]_i_122_0 ;
  wire \iv[15]_i_122_n_0 ;
  wire \iv[15]_i_123_n_0 ;
  wire \iv[15]_i_124_n_0 ;
  wire \iv[15]_i_125_n_0 ;
  wire \iv[15]_i_126_n_0 ;
  wire \iv[15]_i_12_n_0 ;
  wire \iv[15]_i_13_0 ;
  wire \iv[15]_i_13_n_0 ;
  wire \iv[15]_i_14_n_0 ;
  wire \iv[15]_i_158_n_0 ;
  wire \iv[15]_i_159_n_0 ;
  wire \iv[15]_i_15_n_0 ;
  wire \iv[15]_i_160_n_0 ;
  wire \iv[15]_i_161_n_0 ;
  wire \iv[15]_i_162_n_0 ;
  wire \iv[15]_i_16_n_0 ;
  wire \iv[15]_i_173_n_0 ;
  wire \iv[15]_i_174_n_0 ;
  wire \iv[15]_i_175_n_0 ;
  wire \iv[15]_i_176_n_0 ;
  wire \iv[15]_i_177_n_0 ;
  wire \iv[15]_i_17_n_0 ;
  wire \iv[15]_i_18_n_0 ;
  wire \iv[15]_i_19_0 ;
  wire \iv[15]_i_19_1 ;
  wire \iv[15]_i_22 ;
  wire \iv[15]_i_22_0 ;
  wire \iv[15]_i_25_n_0 ;
  wire \iv[15]_i_26_n_0 ;
  wire \iv[15]_i_27_n_0 ;
  wire \iv[15]_i_28_0 ;
  wire \iv[15]_i_28_n_0 ;
  wire \iv[15]_i_29_n_0 ;
  wire \iv[15]_i_30_n_0 ;
  wire \iv[15]_i_31_n_0 ;
  wire \iv[15]_i_32_n_0 ;
  wire \iv[15]_i_33_n_0 ;
  wire \iv[15]_i_34_n_0 ;
  wire \iv[15]_i_35_n_0 ;
  wire \iv[15]_i_36_n_0 ;
  wire \iv[15]_i_37_n_0 ;
  wire \iv[15]_i_38_0 ;
  wire \iv[15]_i_38_n_0 ;
  wire \iv[15]_i_39_n_0 ;
  wire \iv[15]_i_40_n_0 ;
  wire \iv[15]_i_41_n_0 ;
  wire \iv[15]_i_42_n_0 ;
  wire \iv[15]_i_43_n_0 ;
  wire \iv[15]_i_44_n_0 ;
  wire \iv[15]_i_45_n_0 ;
  wire \iv[15]_i_46_n_0 ;
  wire \iv[15]_i_47_n_0 ;
  wire \iv[15]_i_48_n_0 ;
  wire \iv[15]_i_49_n_0 ;
  wire \iv[15]_i_67_n_0 ;
  wire \iv[15]_i_68_n_0 ;
  wire \iv[15]_i_69_n_0 ;
  wire \iv[15]_i_6_n_0 ;
  wire \iv[15]_i_70_n_0 ;
  wire \iv[15]_i_71_n_0 ;
  wire \iv[15]_i_72_n_0 ;
  wire \iv[15]_i_73_n_0 ;
  wire \iv[15]_i_74_n_0 ;
  wire \iv[15]_i_75_n_0 ;
  wire \iv[15]_i_76_n_0 ;
  wire \iv[15]_i_77_n_0 ;
  wire \iv[15]_i_78_n_0 ;
  wire \iv[15]_i_79_n_0 ;
  wire \iv[15]_i_80_n_0 ;
  wire \iv[15]_i_81_n_0 ;
  wire \iv[15]_i_82_n_0 ;
  wire \iv[15]_i_83_n_0 ;
  wire \iv[15]_i_84_n_0 ;
  wire \iv[15]_i_85_n_0 ;
  wire \iv[15]_i_86_n_0 ;
  wire \iv[15]_i_87_n_0 ;
  wire \iv[15]_i_88_n_0 ;
  wire \iv[15]_i_89_n_0 ;
  wire \iv[15]_i_90_n_0 ;
  wire \iv[15]_i_91_n_0 ;
  wire \iv[15]_i_92_n_0 ;
  wire \iv[15]_i_93_n_0 ;
  wire [3:0]\iv[15]_i_9_0 ;
  wire \iv[15]_i_9_n_0 ;
  wire \iv[1]_i_12_n_0 ;
  wire \iv[1]_i_13_n_0 ;
  wire \iv[1]_i_21 ;
  wire \iv[1]_i_21_0 ;
  wire \iv[1]_i_21_1 ;
  wire \iv[1]_i_2_n_0 ;
  wire \iv[1]_i_6_n_0 ;
  wire \iv[1]_i_7_n_0 ;
  wire \iv[2]_i_12_n_0 ;
  wire \iv[2]_i_13_n_0 ;
  wire \iv[2]_i_2_n_0 ;
  wire \iv[2]_i_6_n_0 ;
  wire \iv[2]_i_7_n_0 ;
  wire \iv[3]_i_13_n_0 ;
  wire \iv[3]_i_14_n_0 ;
  wire \iv[3]_i_15_n_0 ;
  wire \iv[3]_i_16 ;
  wire \iv[3]_i_21 ;
  wire \iv[3]_i_2_0 ;
  wire [3:0]\iv[3]_i_2_1 ;
  wire \iv[3]_i_2_n_0 ;
  wire \iv[3]_i_37_n_0 ;
  wire \iv[3]_i_3_n_0 ;
  wire \iv[3]_i_6_n_0 ;
  wire \iv[3]_i_7_n_0 ;
  wire \iv[3]_i_8_0 ;
  wire \iv[4]_i_12_n_0 ;
  wire \iv[4]_i_13_n_0 ;
  wire \iv[4]_i_2_n_0 ;
  wire \iv[4]_i_3_n_0 ;
  wire \iv[4]_i_6_n_0 ;
  wire \iv[4]_i_7_n_0 ;
  wire \iv[4]_i_8 ;
  wire \iv[4]_i_8_0 ;
  wire \iv[5]_i_13_n_0 ;
  wire \iv[5]_i_2_n_0 ;
  wire \iv[5]_i_3_n_0 ;
  wire \iv[5]_i_6_n_0 ;
  wire \iv[5]_i_7_n_0 ;
  wire \iv[5]_i_8 ;
  wire \iv[5]_i_8_0 ;
  wire \iv[6]_i_10_0 ;
  wire \iv[6]_i_10_n_0 ;
  wire \iv[6]_i_13_n_0 ;
  wire \iv[6]_i_14_n_0 ;
  wire \iv[6]_i_15_n_0 ;
  wire \iv[6]_i_20_n_0 ;
  wire \iv[6]_i_21_n_0 ;
  wire \iv[6]_i_22 ;
  wire \iv[6]_i_2_0 ;
  wire \iv[6]_i_2_n_0 ;
  wire \iv[6]_i_3_0 ;
  wire \iv[6]_i_3_1 ;
  wire \iv[6]_i_3_n_0 ;
  wire \iv[6]_i_6_n_0 ;
  wire \iv[6]_i_7_n_0 ;
  wire \iv[6]_i_8_0 ;
  wire \iv[6]_i_8_1 ;
  wire \iv[6]_i_8_n_0 ;
  wire \iv[7]_i_10 ;
  wire \iv[7]_i_10_0 ;
  wire \iv[7]_i_11_0 ;
  wire \iv[7]_i_11_1 ;
  wire \iv[7]_i_11_n_0 ;
  wire \iv[7]_i_14_n_0 ;
  wire \iv[7]_i_15_n_0 ;
  wire \iv[7]_i_27_n_0 ;
  wire \iv[7]_i_28_n_0 ;
  wire [3:0]\iv[7]_i_2_0 ;
  wire \iv[7]_i_2_n_0 ;
  wire \iv[7]_i_34_n_0 ;
  wire \iv[7]_i_3_n_0 ;
  wire \iv[7]_i_6_n_0 ;
  wire \iv[7]_i_7_n_0 ;
  wire \iv[8]_i_10_n_0 ;
  wire \iv[8]_i_17_n_0 ;
  wire \iv[8]_i_18_n_0 ;
  wire \iv[8]_i_19_n_0 ;
  wire \iv[8]_i_22_n_0 ;
  wire \iv[8]_i_2_0 ;
  wire \iv[8]_i_2_n_0 ;
  wire \iv[8]_i_34_0 ;
  wire \iv[8]_i_35 ;
  wire \iv[8]_i_39_n_0 ;
  wire \iv[8]_i_3_n_0 ;
  wire \iv[8]_i_40_n_0 ;
  wire \iv[8]_i_4_0 ;
  wire \iv[8]_i_4_n_0 ;
  wire \iv[8]_i_7_0 ;
  wire \iv[8]_i_7_1 ;
  wire \iv[8]_i_7_n_0 ;
  wire \iv[8]_i_8_n_0 ;
  wire \iv[8]_i_9_n_0 ;
  wire \iv[9]_i_18_n_0 ;
  wire \iv[9]_i_19_n_0 ;
  wire \iv[9]_i_20_n_0 ;
  wire \iv[9]_i_21_n_0 ;
  wire \iv[9]_i_22_n_0 ;
  wire \iv[9]_i_23_n_0 ;
  wire \iv[9]_i_24_n_0 ;
  wire \iv[9]_i_2_n_0 ;
  wire \iv[9]_i_35 ;
  wire \iv[9]_i_3_n_0 ;
  wire \iv[9]_i_42_n_0 ;
  wire \iv[9]_i_7_0 ;
  wire \iv[9]_i_7_n_0 ;
  wire \iv[9]_i_8_n_0 ;
  wire \iv[9]_i_9_n_0 ;
  wire \iv_reg[0] ;
  wire \iv_reg[0]_0 ;
  wire \iv_reg[0]_1 ;
  wire \iv_reg[11]_i_22_n_0 ;
  wire \iv_reg[14]_i_23_n_0 ;
  wire \iv_reg[8]_i_23_n_0 ;
  wire [15:0]\mul_a_reg[15] ;
  wire mul_b;
  wire \mul_b_reg[10] ;
  wire \mul_b_reg[10]_0 ;
  wire \mul_b_reg[11] ;
  wire \mul_b_reg[11]_0 ;
  wire \mul_b_reg[12] ;
  wire \mul_b_reg[12]_0 ;
  wire \mul_b_reg[13] ;
  wire \mul_b_reg[13]_0 ;
  wire \mul_b_reg[14] ;
  wire \mul_b_reg[14]_0 ;
  wire \mul_b_reg[15] ;
  wire \mul_b_reg[15]_0 ;
  wire \mul_b_reg[15]_1 ;
  wire \mul_b_reg[1] ;
  wire \mul_b_reg[1]_0 ;
  wire \mul_b_reg[1]_1 ;
  wire \mul_b_reg[2] ;
  wire \mul_b_reg[2]_0 ;
  wire \mul_b_reg[2]_1 ;
  wire \mul_b_reg[31] ;
  wire \mul_b_reg[31]_0 ;
  wire \mul_b_reg[3] ;
  wire \mul_b_reg[3]_0 ;
  wire \mul_b_reg[3]_1 ;
  wire \mul_b_reg[4] ;
  wire \mul_b_reg[4]_0 ;
  wire \mul_b_reg[4]_1 ;
  wire \mul_b_reg[6] ;
  wire \mul_b_reg[6]_0 ;
  wire \mul_b_reg[7] ;
  wire \mul_b_reg[7]_0 ;
  wire \mul_b_reg[8] ;
  wire \mul_b_reg[8]_0 ;
  wire \mul_b_reg[9] ;
  wire \mul_b_reg[9]_0 ;
  wire mul_rslt;
  wire [15:0]mulh;
  wire \niho_dsp_a[15]_INST_0_i_2_0 ;
  wire \niho_dsp_a[32]_INST_0_i_10_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_11_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_12_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_13_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_14_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_15_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_17_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_18_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_3_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_4_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_5_0 ;
  wire \niho_dsp_a[32]_INST_0_i_5_1 ;
  wire \niho_dsp_a[32]_INST_0_i_5_2 ;
  wire \niho_dsp_a[32]_INST_0_i_5_3 ;
  wire \niho_dsp_a[32]_INST_0_i_5_4 ;
  wire \niho_dsp_a[32]_INST_0_i_6_0 ;
  wire \niho_dsp_a[32]_INST_0_i_7_0 ;
  wire \niho_dsp_a[32]_INST_0_i_8_n_0 ;
  wire \niho_dsp_a[32]_INST_0_i_9_0 ;
  wire \niho_dsp_a[32]_INST_0_i_9_n_0 ;
  wire [29:0]niho_dsp_b;
  wire \niho_dsp_b[30] ;
  wire [1:0]\niho_dsp_b[32] ;
  wire niho_dsp_b_10_sn_1;
  wire niho_dsp_b_11_sn_1;
  wire niho_dsp_b_12_sn_1;
  wire niho_dsp_b_13_sn_1;
  wire niho_dsp_b_14_sn_1;
  wire niho_dsp_b_15_sn_1;
  wire niho_dsp_b_16_sn_1;
  wire niho_dsp_b_17_sn_1;
  wire niho_dsp_b_18_sn_1;
  wire niho_dsp_b_19_sn_1;
  wire niho_dsp_b_1_sn_1;
  wire niho_dsp_b_20_sn_1;
  wire niho_dsp_b_21_sn_1;
  wire niho_dsp_b_22_sn_1;
  wire niho_dsp_b_23_sn_1;
  wire niho_dsp_b_24_sn_1;
  wire niho_dsp_b_25_sn_1;
  wire niho_dsp_b_26_sn_1;
  wire niho_dsp_b_27_sn_1;
  wire niho_dsp_b_28_sn_1;
  wire niho_dsp_b_29_sn_1;
  wire niho_dsp_b_2_sn_1;
  wire niho_dsp_b_3_sn_1;
  wire niho_dsp_b_6_sn_1;
  wire niho_dsp_b_7_sn_1;
  wire niho_dsp_b_8_sn_1;
  wire niho_dsp_b_9_sn_1;
  wire [24:0]niho_dsp_c;
  wire p_0_in;
  wire [30:17]p_2_in;
  wire [15:0]\pc_reg[15] ;
  wire [2:0]read_cyc;
  wire [1:1]\rgf/cbus_sel_cr ;
  wire [15:0]rgf_pc;
  wire rst_n;
  wire [1:0]rst_n_0;
  wire rst_n_1;
  wire rst_n_2;
  wire rst_n_fl;
  wire rst_n_fl_reg_0;
  wire rst_n_fl_reg_1;
  wire rst_n_fl_reg_10;
  wire rst_n_fl_reg_11;
  wire rst_n_fl_reg_12;
  wire rst_n_fl_reg_13;
  wire rst_n_fl_reg_14;
  wire rst_n_fl_reg_15;
  wire rst_n_fl_reg_16;
  wire rst_n_fl_reg_17;
  wire rst_n_fl_reg_18;
  wire rst_n_fl_reg_19;
  wire rst_n_fl_reg_2;
  wire rst_n_fl_reg_20;
  wire rst_n_fl_reg_21;
  wire rst_n_fl_reg_22;
  wire rst_n_fl_reg_23;
  wire rst_n_fl_reg_3;
  wire rst_n_fl_reg_4;
  wire rst_n_fl_reg_5;
  wire rst_n_fl_reg_6;
  wire rst_n_fl_reg_7;
  wire rst_n_fl_reg_8;
  wire rst_n_fl_reg_9;
  wire \sp[0]_i_10_n_0 ;
  wire \sp[0]_i_11_n_0 ;
  wire \sp[0]_i_12_n_0 ;
  wire \sp[0]_i_13_0 ;
  wire \sp[0]_i_13_n_0 ;
  wire \sp[0]_i_14_n_0 ;
  wire \sp[0]_i_15_n_0 ;
  wire \sp[0]_i_16_n_0 ;
  wire \sp[0]_i_6_n_0 ;
  wire \sp[0]_i_7_n_0 ;
  wire \sp[0]_i_8_n_0 ;
  wire \sp[31]_i_10_n_0 ;
  wire \sp[31]_i_11_n_0 ;
  wire \sp[31]_i_6_n_0 ;
  wire \sp[31]_i_7_n_0 ;
  wire \sp[31]_i_8_n_0 ;
  wire \sp[31]_i_9_n_0 ;
  wire [0:0]\sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[16] ;
  wire \sp_reg[17] ;
  wire \sp_reg[18] ;
  wire \sp_reg[1] ;
  wire \sp_reg[20] ;
  wire \sp_reg[22] ;
  wire \sp_reg[24] ;
  wire \sp_reg[25] ;
  wire \sp_reg[26] ;
  wire \sp_reg[2] ;
  wire \sp_reg[30] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[12]_i_2_n_0 ;
  wire \sr[13]_i_2_n_0 ;
  wire \sr[13]_i_3_n_0 ;
  wire \sr[13]_i_4_n_0 ;
  wire \sr[13]_i_6_n_0 ;
  wire \sr[13]_i_7_n_0 ;
  wire \sr[13]_i_8_n_0 ;
  wire \sr[2]_i_2_n_0 ;
  wire \sr[3]_i_2_n_0 ;
  wire \sr[4]_i_10_0 ;
  wire \sr[4]_i_10_1 ;
  wire \sr[4]_i_10_n_0 ;
  wire \sr[4]_i_115_n_0 ;
  wire \sr[4]_i_117_n_0 ;
  wire \sr[4]_i_124_n_0 ;
  wire \sr[4]_i_126_n_0 ;
  wire \sr[4]_i_131_n_0 ;
  wire \sr[4]_i_133_n_0 ;
  wire \sr[4]_i_146_n_0 ;
  wire \sr[4]_i_148_n_0 ;
  wire \sr[4]_i_157_n_0 ;
  wire \sr[4]_i_161_n_0 ;
  wire \sr[4]_i_166_n_0 ;
  wire \sr[4]_i_18_0 ;
  wire \sr[4]_i_18_1 ;
  wire \sr[4]_i_18_2 ;
  wire \sr[4]_i_18_3 ;
  wire \sr[4]_i_18_4 ;
  wire \sr[4]_i_18_5 ;
  wire \sr[4]_i_18_6 ;
  wire \sr[4]_i_18_7 ;
  wire \sr[4]_i_18_8 ;
  wire \sr[4]_i_18_9 ;
  wire \sr[4]_i_19 ;
  wire \sr[4]_i_19_0 ;
  wire \sr[4]_i_19_1 ;
  wire \sr[4]_i_20 ;
  wire \sr[4]_i_21 ;
  wire \sr[4]_i_22_n_0 ;
  wire \sr[4]_i_23_n_0 ;
  wire \sr[4]_i_24_0 ;
  wire \sr[4]_i_24_1 ;
  wire \sr[4]_i_24_2 ;
  wire \sr[4]_i_24_n_0 ;
  wire \sr[4]_i_25_n_0 ;
  wire \sr[4]_i_26_n_0 ;
  wire \sr[4]_i_27_n_0 ;
  wire \sr[4]_i_2_n_0 ;
  wire \sr[4]_i_37_0 ;
  wire \sr[4]_i_37_1 ;
  wire \sr[4]_i_37_n_0 ;
  wire \sr[4]_i_38 ;
  wire \sr[4]_i_38_0 ;
  wire \sr[4]_i_39_0 ;
  wire \sr[4]_i_39_n_0 ;
  wire \sr[4]_i_3_n_0 ;
  wire \sr[4]_i_40_0 ;
  wire \sr[4]_i_40_1 ;
  wire \sr[4]_i_40_n_0 ;
  wire \sr[4]_i_41 ;
  wire \sr[4]_i_43_0 ;
  wire \sr[4]_i_43_1 ;
  wire \sr[4]_i_44 ;
  wire \sr[4]_i_44_0 ;
  wire \sr[4]_i_45 ;
  wire \sr[4]_i_45_0 ;
  wire \sr[4]_i_46 ;
  wire \sr[4]_i_46_0 ;
  wire \sr[4]_i_5 ;
  wire \sr[4]_i_5_0 ;
  wire \sr[4]_i_5_1 ;
  wire \sr[4]_i_66_0 ;
  wire \sr[4]_i_66_1 ;
  wire \sr[4]_i_66_2 ;
  wire \sr[4]_i_66_n_0 ;
  wire \sr[4]_i_69 ;
  wire \sr[4]_i_6_n_0 ;
  wire \sr[4]_i_74_0 ;
  wire \sr[4]_i_74_1 ;
  wire \sr[4]_i_74_n_0 ;
  wire \sr[4]_i_77 ;
  wire \sr[4]_i_78_0 ;
  wire \sr[4]_i_78_1 ;
  wire \sr[4]_i_78_n_0 ;
  wire \sr[4]_i_7_0 ;
  wire \sr[4]_i_7_1 ;
  wire \sr[4]_i_7_2 ;
  wire \sr[4]_i_7_3 ;
  wire \sr[4]_i_7_4 ;
  wire \sr[4]_i_7_n_0 ;
  wire \sr[4]_i_80 ;
  wire \sr[4]_i_81 ;
  wire \sr[4]_i_81_0 ;
  wire \sr[4]_i_81_1 ;
  wire \sr[4]_i_85 ;
  wire \sr[4]_i_85_0 ;
  wire \sr[4]_i_85_1 ;
  wire \sr[4]_i_8_0 ;
  wire \sr[4]_i_8_n_0 ;
  wire \sr[4]_i_91_0 ;
  wire \sr[4]_i_91_1 ;
  wire \sr[4]_i_91_2 ;
  wire \sr[4]_i_91_3 ;
  wire \sr[4]_i_91_n_0 ;
  wire \sr[4]_i_98 ;
  wire \sr[4]_i_9_n_0 ;
  wire \sr[5]_i_3_n_0 ;
  wire \sr[5]_i_8_n_0 ;
  wire \sr[5]_i_9_n_0 ;
  wire \sr[6]_i_14_n_0 ;
  wire \sr[6]_i_25_0 ;
  wire \sr[6]_i_25_n_0 ;
  wire \sr[6]_i_2_n_0 ;
  wire \sr[6]_i_32_n_0 ;
  wire \sr[7]_i_15_n_0 ;
  wire \sr[7]_i_20_0 ;
  wire \sr[7]_i_21 ;
  wire \sr[7]_i_23_n_0 ;
  wire \sr[7]_i_31_n_0 ;
  wire \sr[7]_i_32_n_0 ;
  wire \sr[7]_i_3_n_0 ;
  wire \sr[7]_i_44_n_0 ;
  wire [0:0]\sr[7]_i_4_0 ;
  wire \sr[7]_i_4_n_0 ;
  wire \sr[7]_i_5_n_0 ;
  wire \sr[7]_i_6_n_0 ;
  wire \sr[7]_i_7 ;
  wire \sr[7]_i_7_0 ;
  wire \sr[7]_i_8_n_0 ;
  wire \sr_reg[0] ;
  wire \sr_reg[10] ;
  wire \sr_reg[11] ;
  wire [12:0]\sr_reg[13] ;
  wire \sr_reg[1] ;
  wire [0:0]\sr_reg[1]_0 ;
  wire [0:0]\sr_reg[1]_1 ;
  wire [0:0]\sr_reg[1]_10 ;
  wire [0:0]\sr_reg[1]_11 ;
  wire [0:0]\sr_reg[1]_12 ;
  wire [0:0]\sr_reg[1]_13 ;
  wire [0:0]\sr_reg[1]_14 ;
  wire [0:0]\sr_reg[1]_15 ;
  wire [0:0]\sr_reg[1]_16 ;
  wire [0:0]\sr_reg[1]_17 ;
  wire [0:0]\sr_reg[1]_18 ;
  wire [0:0]\sr_reg[1]_19 ;
  wire [0:0]\sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_20 ;
  wire [0:0]\sr_reg[1]_21 ;
  wire [0:0]\sr_reg[1]_22 ;
  wire [0:0]\sr_reg[1]_3 ;
  wire [0:0]\sr_reg[1]_4 ;
  wire [0:0]\sr_reg[1]_5 ;
  wire [0:0]\sr_reg[1]_6 ;
  wire [0:0]\sr_reg[1]_7 ;
  wire [0:0]\sr_reg[1]_8 ;
  wire [0:0]\sr_reg[1]_9 ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_51 ;
  wire \sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire \sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire \sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_60 ;
  wire \sr_reg[8]_61 ;
  wire \sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire \sr_reg[8]_71 ;
  wire [8:0]\sr_reg[8]_72 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;
  wire \stat[0]_i_10_n_0 ;
  wire \stat[0]_i_11_n_0 ;
  wire \stat[0]_i_12_n_0 ;
  wire \stat[0]_i_13_n_0 ;
  wire \stat[0]_i_14_n_0 ;
  wire \stat[0]_i_15_n_0 ;
  wire \stat[0]_i_16_n_0 ;
  wire \stat[0]_i_18_n_0 ;
  wire \stat[0]_i_20_n_0 ;
  wire \stat[0]_i_21_n_0 ;
  wire \stat[0]_i_22_n_0 ;
  wire \stat[0]_i_23_n_0 ;
  wire \stat[0]_i_24_n_0 ;
  wire \stat[0]_i_25_n_0 ;
  wire \stat[0]_i_26_n_0 ;
  wire \stat[0]_i_27_n_0 ;
  wire \stat[0]_i_28_n_0 ;
  wire \stat[0]_i_29_n_0 ;
  wire \stat[0]_i_2_0 ;
  wire \stat[0]_i_2_n_0 ;
  wire \stat[0]_i_30_n_0 ;
  wire \stat[0]_i_31_n_0 ;
  wire \stat[0]_i_32_n_0 ;
  wire \stat[0]_i_33_n_0 ;
  wire \stat[0]_i_34_n_0 ;
  wire \stat[0]_i_35_n_0 ;
  wire \stat[0]_i_36_n_0 ;
  wire \stat[0]_i_4_n_0 ;
  wire \stat[0]_i_5_n_0 ;
  wire \stat[0]_i_6_n_0 ;
  wire \stat[0]_i_7_n_0 ;
  wire \stat[0]_i_8_n_0 ;
  wire \stat[0]_i_9_n_0 ;
  wire \stat[1]_i_10_0 ;
  wire \stat[1]_i_10_n_0 ;
  wire \stat[1]_i_11_n_0 ;
  wire \stat[1]_i_13_n_0 ;
  wire \stat[1]_i_14_n_0 ;
  wire \stat[1]_i_15_n_0 ;
  wire \stat[1]_i_16_n_0 ;
  wire \stat[1]_i_17_n_0 ;
  wire \stat[1]_i_18_n_0 ;
  wire \stat[1]_i_19_n_0 ;
  wire \stat[1]_i_20_n_0 ;
  wire \stat[1]_i_21_n_0 ;
  wire \stat[1]_i_22_n_0 ;
  wire \stat[1]_i_23_n_0 ;
  wire \stat[1]_i_24_n_0 ;
  wire \stat[1]_i_25_n_0 ;
  wire \stat[1]_i_26_n_0 ;
  wire \stat[1]_i_2_n_0 ;
  wire \stat[1]_i_3_n_0 ;
  wire \stat[1]_i_5_n_0 ;
  wire \stat[1]_i_6_0 ;
  wire \stat[1]_i_6_n_0 ;
  wire \stat[1]_i_7_n_0 ;
  wire \stat[1]_i_8_n_0 ;
  wire \stat[1]_i_9_n_0 ;
  wire \stat[2]_i_11_n_0 ;
  wire \stat[2]_i_3_n_0 ;
  wire \stat[2]_i_6_n_0 ;
  wire \stat[2]_i_9_n_0 ;
  wire \stat_reg[0] ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_10 ;
  wire \stat_reg[0]_11 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[0]_7 ;
  wire \stat_reg[0]_8 ;
  wire \stat_reg[0]_9 ;
  wire \stat_reg[1] ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[2] ;
  wire [2:0]\stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_10 ;
  wire \stat_reg[2]_11 ;
  wire [2:0]\stat_reg[2]_12 ;
  wire \stat_reg[2]_13 ;
  wire \stat_reg[2]_14 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;
  wire [2:0]\stat_reg[2]_5 ;
  wire \stat_reg[2]_6 ;
  wire \stat_reg[2]_7 ;
  wire \stat_reg[2]_8 ;
  wire \stat_reg[2]_9 ;
  wire \tr[16]_i_18_n_0 ;
  wire \tr[16]_i_19_n_0 ;
  wire \tr[16]_i_21_n_0 ;
  wire \tr[16]_i_22_n_0 ;
  wire \tr[16]_i_3_0 ;
  wire \tr[16]_i_3_n_0 ;
  wire \tr[16]_i_7_0 ;
  wire \tr[16]_i_7_1 ;
  wire \tr[16]_i_7_n_0 ;
  wire \tr[16]_i_8_n_0 ;
  wire \tr[17]_i_11_n_0 ;
  wire \tr[17]_i_12_n_0 ;
  wire \tr[17]_i_13_n_0 ;
  wire \tr[17]_i_15_n_0 ;
  wire \tr[17]_i_2_0 ;
  wire \tr[17]_i_3 ;
  wire \tr[17]_i_3_0 ;
  wire \tr[17]_i_4_n_0 ;
  wire \tr[17]_i_5_0 ;
  wire \tr[17]_i_5_n_0 ;
  wire \tr[18]_i_11_n_0 ;
  wire \tr[18]_i_12_n_0 ;
  wire \tr[18]_i_13_n_0 ;
  wire \tr[18]_i_15_n_0 ;
  wire \tr[18]_i_2_0 ;
  wire \tr[18]_i_2_1 ;
  wire \tr[18]_i_3 ;
  wire \tr[18]_i_3_0 ;
  wire \tr[18]_i_4_n_0 ;
  wire \tr[18]_i_5_0 ;
  wire \tr[18]_i_5_1 ;
  wire \tr[18]_i_5_n_0 ;
  wire \tr[19]_i_10_n_0 ;
  wire \tr[19]_i_11_n_0 ;
  wire \tr[19]_i_12_n_0 ;
  wire \tr[19]_i_14_0 ;
  wire \tr[19]_i_14_n_0 ;
  wire \tr[19]_i_3 ;
  wire \tr[19]_i_3_0 ;
  wire \tr[19]_i_5_0 ;
  wire \tr[19]_i_5_1 ;
  wire \tr[19]_i_9 ;
  wire \tr[20]_i_11_n_0 ;
  wire \tr[20]_i_12_n_0 ;
  wire \tr[20]_i_14_n_0 ;
  wire \tr[20]_i_15_n_0 ;
  wire \tr[20]_i_2_0 ;
  wire \tr[20]_i_3 ;
  wire \tr[20]_i_4_n_0 ;
  wire \tr[20]_i_5_0 ;
  wire \tr[20]_i_5_1 ;
  wire \tr[20]_i_5_n_0 ;
  wire \tr[20]_i_7 ;
  wire \tr[21]_i_10_n_0 ;
  wire \tr[21]_i_11_n_0 ;
  wire \tr[21]_i_13_n_0 ;
  wire \tr[21]_i_14_0 ;
  wire \tr[21]_i_14_n_0 ;
  wire \tr[21]_i_2 ;
  wire \tr[21]_i_3 ;
  wire \tr[21]_i_5_0 ;
  wire \tr[21]_i_5_1 ;
  wire \tr[21]_i_7 ;
  wire \tr[22]_i_11_n_0 ;
  wire \tr[22]_i_12_n_0 ;
  wire \tr[22]_i_13_n_0 ;
  wire \tr[22]_i_14_n_0 ;
  wire \tr[22]_i_16_n_0 ;
  wire \tr[22]_i_2_0 ;
  wire \tr[22]_i_3 ;
  wire \tr[22]_i_4_n_0 ;
  wire \tr[22]_i_5_0 ;
  wire \tr[22]_i_5_1 ;
  wire \tr[22]_i_5_n_0 ;
  wire \tr[22]_i_7_0 ;
  wire \tr[23]_i_12_n_0 ;
  wire \tr[23]_i_14_n_0 ;
  wire \tr[23]_i_15_0 ;
  wire \tr[23]_i_15_n_0 ;
  wire \tr[23]_i_2 ;
  wire \tr[23]_i_24_n_0 ;
  wire \tr[23]_i_25_n_0 ;
  wire \tr[23]_i_3 ;
  wire \tr[23]_i_3_0 ;
  wire \tr[23]_i_5_0 ;
  wire \tr[24]_i_12_n_0 ;
  wire \tr[24]_i_14_n_0 ;
  wire \tr[24]_i_15_n_0 ;
  wire \tr[24]_i_17_n_0 ;
  wire \tr[24]_i_18_n_0 ;
  wire \tr[24]_i_2_0 ;
  wire \tr[24]_i_3 ;
  wire \tr[24]_i_4_n_0 ;
  wire \tr[24]_i_5_0 ;
  wire \tr[24]_i_5_n_0 ;
  wire \tr[24]_i_7 ;
  wire \tr[25]_i_12_n_0 ;
  wire \tr[25]_i_13_n_0 ;
  wire \tr[25]_i_14_n_0 ;
  wire \tr[25]_i_15_n_0 ;
  wire \tr[25]_i_16_n_0 ;
  wire \tr[25]_i_2_0 ;
  wire \tr[25]_i_4_n_0 ;
  wire \tr[25]_i_5_0 ;
  wire \tr[25]_i_5_1 ;
  wire \tr[25]_i_5_n_0 ;
  wire \tr[26]_i_11_n_0 ;
  wire \tr[26]_i_12_n_0 ;
  wire \tr[26]_i_14_n_0 ;
  wire \tr[26]_i_16_n_0 ;
  wire \tr[26]_i_17_n_0 ;
  wire \tr[26]_i_2_0 ;
  wire \tr[26]_i_4_n_0 ;
  wire \tr[26]_i_5_n_0 ;
  wire \tr[27]_i_10_n_0 ;
  wire \tr[27]_i_11_n_0 ;
  wire \tr[27]_i_12_n_0 ;
  wire \tr[27]_i_13_n_0 ;
  wire \tr[27]_i_14 ;
  wire \tr[27]_i_5_0 ;
  wire \tr[27]_i_5_1 ;
  wire \tr[28]_i_10_n_0 ;
  wire \tr[28]_i_12_n_0 ;
  wire \tr[28]_i_13_0 ;
  wire \tr[28]_i_13_n_0 ;
  wire \tr[28]_i_14_n_0 ;
  wire \tr[28]_i_15_n_0 ;
  wire \tr[28]_i_16_n_0 ;
  wire \tr[28]_i_3 ;
  wire \tr[28]_i_9_0 ;
  wire \tr[29]_i_11_n_0 ;
  wire \tr[29]_i_13_n_0 ;
  wire \tr[29]_i_14_0 ;
  wire \tr[29]_i_14_n_0 ;
  wire \tr[29]_i_16_n_0 ;
  wire \tr[29]_i_17_n_0 ;
  wire \tr[29]_i_7 ;
  wire \tr[30]_i_12_n_0 ;
  wire \tr[30]_i_13_n_0 ;
  wire \tr[30]_i_15_n_0 ;
  wire \tr[30]_i_19_n_0 ;
  wire \tr[30]_i_20_n_0 ;
  wire \tr[30]_i_21_n_0 ;
  wire [24:0]\tr[30]_i_2_0 ;
  wire \tr[30]_i_2_1 ;
  wire \tr[30]_i_5_n_0 ;
  wire \tr[30]_i_6_n_0 ;
  wire \tr[30]_i_8 ;
  wire \tr[31]_i_10_n_0 ;
  wire \tr[31]_i_11_n_0 ;
  wire \tr[31]_i_12_0 ;
  wire \tr[31]_i_12_n_0 ;
  wire \tr[31]_i_16_n_0 ;
  wire \tr[31]_i_17_n_0 ;
  wire \tr[31]_i_18_n_0 ;
  wire \tr[31]_i_19_n_0 ;
  wire \tr[31]_i_20_n_0 ;
  wire \tr[31]_i_21_n_0 ;
  wire \tr[31]_i_22_n_0 ;
  wire \tr[31]_i_23_n_0 ;
  wire \tr[31]_i_24_n_0 ;
  wire \tr[31]_i_25_n_0 ;
  wire \tr[31]_i_26_n_0 ;
  wire \tr[31]_i_27_n_0 ;
  wire \tr[31]_i_28_n_0 ;
  wire \tr[31]_i_29_n_0 ;
  wire \tr[31]_i_30_n_0 ;
  wire \tr[31]_i_31_n_0 ;
  wire \tr[31]_i_41_n_0 ;
  wire \tr[31]_i_42_n_0 ;
  wire \tr[31]_i_44_0 ;
  wire \tr[31]_i_44_n_0 ;
  wire \tr[31]_i_45_n_0 ;
  wire \tr[31]_i_46_n_0 ;
  wire \tr[31]_i_47_n_0 ;
  wire \tr[31]_i_48_n_0 ;
  wire \tr[31]_i_49_n_0 ;
  wire \tr[31]_i_50_n_0 ;
  wire \tr[31]_i_51_n_0 ;
  wire \tr[31]_i_52_n_0 ;
  wire \tr[31]_i_53_n_0 ;
  wire \tr[31]_i_54_n_0 ;
  wire \tr[31]_i_55_n_0 ;
  wire \tr[31]_i_56_n_0 ;
  wire \tr[31]_i_58_n_0 ;
  wire \tr[31]_i_59_n_0 ;
  wire \tr[31]_i_60_n_0 ;
  wire \tr[31]_i_61_n_0 ;
  wire \tr[31]_i_6_n_0 ;
  wire \tr[31]_i_70_n_0 ;
  wire \tr[31]_i_71_n_0 ;
  wire \tr[31]_i_72_n_0 ;
  wire \tr[31]_i_73_n_0 ;
  wire \tr[31]_i_74_n_0 ;
  wire \tr[31]_i_75_n_0 ;
  wire \tr[31]_i_76_n_0 ;
  wire \tr[31]_i_77_n_0 ;
  wire \tr[31]_i_7_n_0 ;
  wire \tr[31]_i_8_n_0 ;
  wire \tr[31]_i_9_n_0 ;
  wire \tr_reg[0] ;
  wire \tr_reg[0]_0 ;
  wire \tr_reg[0]_1 ;
  wire \tr_reg[0]_2 ;
  wire \tr_reg[0]_3 ;
  wire \tr_reg[0]_4 ;
  wire \tr_reg[10] ;
  wire \tr_reg[10]_0 ;
  wire \tr_reg[10]_1 ;
  wire \tr_reg[11] ;
  wire \tr_reg[11]_0 ;
  wire \tr_reg[11]_1 ;
  wire \tr_reg[11]_2 ;
  wire \tr_reg[12] ;
  wire \tr_reg[12]_0 ;
  wire \tr_reg[13] ;
  wire \tr_reg[13]_0 ;
  wire \tr_reg[13]_1 ;
  wire \tr_reg[14] ;
  wire \tr_reg[14]_0 ;
  wire \tr_reg[14]_1 ;
  wire \tr_reg[15] ;
  wire \tr_reg[15]_0 ;
  wire \tr_reg[15]_1 ;
  wire \tr_reg[15]_2 ;
  wire \tr_reg[15]_3 ;
  wire \tr_reg[16] ;
  wire \tr_reg[16]_0 ;
  wire \tr_reg[17] ;
  wire \tr_reg[17]_0 ;
  wire \tr_reg[18] ;
  wire \tr_reg[18]_0 ;
  wire \tr_reg[19] ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[1]_1 ;
  wire \tr_reg[1]_2 ;
  wire \tr_reg[20] ;
  wire \tr_reg[20]_0 ;
  wire \tr_reg[21] ;
  wire \tr_reg[22] ;
  wire \tr_reg[22]_0 ;
  wire \tr_reg[23] ;
  wire \tr_reg[24] ;
  wire \tr_reg[24]_0 ;
  wire \tr_reg[25] ;
  wire \tr_reg[25]_0 ;
  wire \tr_reg[26] ;
  wire \tr_reg[26]_0 ;
  wire \tr_reg[27] ;
  wire \tr_reg[28] ;
  wire \tr_reg[29] ;
  wire \tr_reg[2] ;
  wire \tr_reg[2]_0 ;
  wire \tr_reg[2]_1 ;
  wire \tr_reg[2]_2 ;
  wire \tr_reg[30] ;
  wire \tr_reg[30]_0 ;
  wire \tr_reg[30]_1 ;
  wire \tr_reg[31] ;
  wire \tr_reg[3] ;
  wire \tr_reg[3]_0 ;
  wire \tr_reg[3]_1 ;
  wire \tr_reg[3]_2 ;
  wire \tr_reg[3]_3 ;
  wire \tr_reg[4] ;
  wire \tr_reg[4]_0 ;
  wire \tr_reg[4]_1 ;
  wire \tr_reg[4]_2 ;
  wire \tr_reg[4]_3 ;
  wire \tr_reg[4]_4 ;
  wire \tr_reg[5] ;
  wire \tr_reg[5]_0 ;
  wire \tr_reg[5]_1 ;
  wire \tr_reg[5]_2 ;
  wire \tr_reg[5]_3 ;
  wire \tr_reg[5]_4 ;
  wire \tr_reg[6] ;
  wire \tr_reg[6]_0 ;
  wire \tr_reg[6]_1 ;
  wire \tr_reg[6]_2 ;
  wire \tr_reg[7] ;
  wire \tr_reg[7]_0 ;
  wire \tr_reg[7]_1 ;
  wire \tr_reg[7]_2 ;
  wire \tr_reg[7]_3 ;
  wire \tr_reg[7]_4 ;
  wire \tr_reg[8] ;
  wire \tr_reg[8]_0 ;
  wire \tr_reg[8]_1 ;
  wire \tr_reg[9] ;
  wire \tr_reg[9]_0 ;
  wire \tr_reg[9]_1 ;
  wire \tr_reg[9]_2 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_23 
       (.I0(abus_0[3]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[2]),
        .O(\bdatw[11]_INST_0_i_1_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_24 
       (.I0(abus_0[2]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[1]),
        .O(\bdatw[11]_INST_0_i_1_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_25 
       (.I0(abus_0[1]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[0]),
        .O(\bdatw[11]_INST_0_i_1_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_29 
       (.I0(abus_0[7]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[5]),
        .O(\bdatw[15]_INST_0_i_1_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_30 
       (.I0(abus_0[6]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[4]),
        .O(\bdatw[15]_INST_0_i_1_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_32 
       (.I0(abus_0[4]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[3]),
        .O(\bdatw[15]_INST_0_i_1_0 [0]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_11 
       (.I0(abus_0[15]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[13]),
        .O(S[3]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_12 
       (.I0(abus_0[14]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[12]),
        .O(S[2]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_13 
       (.I0(abus_0[13]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[11]),
        .O(S[1]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_14 
       (.I0(abus_0[12]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[10]),
        .O(S[0]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_15 
       (.I0(abus_0[11]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[9]),
        .O(\bdatw[11]_INST_0_i_2_0 [3]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_16 
       (.I0(abus_0[10]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[8]),
        .O(\bdatw[11]_INST_0_i_2_0 [2]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_17 
       (.I0(abus_0[9]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[7]),
        .O(\bdatw[11]_INST_0_i_2_0 [1]));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/sr[5]_i_18 
       (.I0(abus_0[8]),
        .I1(\stat_reg[2]_3 ),
        .I2(bbus_0[6]),
        .O(\bdatw[11]_INST_0_i_2_0 [0]));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[0]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[0]),
        .O(badr[0]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[0]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [0]),
        .I5(\mul_a_reg[15] [0]),
        .O(\tr_reg[0] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[10]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[10]),
        .O(badr[10]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[10]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [10]),
        .I5(\mul_a_reg[15] [10]),
        .O(\tr_reg[10] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[11]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[11]),
        .O(badr[11]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[11]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [11]),
        .I5(\mul_a_reg[15] [11]),
        .O(\tr_reg[11] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[12]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[12]),
        .O(badr[12]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[12]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [12]),
        .I5(\mul_a_reg[15] [12]),
        .O(\tr_reg[12] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[13]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[13]),
        .O(badr[13]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[13]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [13]),
        .I5(\mul_a_reg[15] [13]),
        .O(\tr_reg[13] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[14]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[14]),
        .O(badr[14]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[14]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [14]),
        .I5(\mul_a_reg[15] [14]),
        .O(\tr_reg[14] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[15]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[15]),
        .O(badr[15]));
  LUT4 #(
    .INIT(16'h0001)) 
    \badr[15]_INST_0_i_16 
       (.I0(\badr[31]_INST_0_i_12_n_0 ),
        .I1(ctl_sela_rn),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(abus_sel_cr[0]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[15]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [15]),
        .I5(\mul_a_reg[15] [15]),
        .O(\tr_reg[15] ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[15]_INST_0_i_21 
       (.I0(\badr[31]_INST_0_i_29_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(ctl_sela_rn),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(abus_sel_cr[1]));
  LUT2 #(
    .INIT(4'h7)) 
    \badr[15]_INST_0_i_7 
       (.I0(\badr[31]_INST_0_i_29_n_0 ),
        .I1(ctl_sela_rn),
        .O(\badr[15]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[16]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(\badr[31]_INST_0_i_1 [0]),
        .I3(abus_0[16]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[16]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[16]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [16]),
        .O(\tr_reg[16] ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[17]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(\badr[31]_INST_0_i_1 [1]),
        .I3(abus_0[17]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[17]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[17]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [17]),
        .O(\tr_reg[17] ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[18]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(\badr[31]_INST_0_i_1 [2]),
        .I3(abus_0[18]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[18]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[18]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [18]),
        .O(\tr_reg[18] ));
  LUT5 #(
    .INIT(32'hF0F0EE00)) 
    \badr[19]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(\badr[31]_INST_0_i_1 [3]),
        .I3(abus_0[19]),
        .I4(\badr[31]_INST_0_i_2_n_0 ),
        .O(badr[19]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[19]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [19]),
        .O(\tr_reg[19] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[1]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[1]),
        .O(badr[1]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[1]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [1]),
        .I5(\mul_a_reg[15] [1]),
        .O(\tr_reg[1] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[20]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[20]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [4]),
        .O(badr[20]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[20]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [20]),
        .O(\tr_reg[20] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[21]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[21]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [5]),
        .O(badr[21]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[21]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [21]),
        .O(\tr_reg[21] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[22]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[22]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [6]),
        .O(badr[22]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[22]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [22]),
        .O(\tr_reg[22] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[23]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[23]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [7]),
        .O(badr[23]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[23]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [23]),
        .O(\tr_reg[23] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[24]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[24]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [8]),
        .O(badr[24]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[24]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [24]),
        .O(\tr_reg[24] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[25]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[25]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [9]),
        .O(badr[25]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[25]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [25]),
        .O(\tr_reg[25] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[26]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[26]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [10]),
        .O(badr[26]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[26]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [26]),
        .O(\tr_reg[26] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[27]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[27]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [11]),
        .O(badr[27]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[27]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [27]),
        .O(\tr_reg[27] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[28]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[28]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [12]),
        .O(badr[28]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[28]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [28]),
        .O(\tr_reg[28] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[29]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[29]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [13]),
        .O(badr[29]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[29]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [29]),
        .O(\tr_reg[29] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[2]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[2]),
        .O(badr[2]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[2]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [2]),
        .I5(\mul_a_reg[15] [2]),
        .O(\tr_reg[2] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[30]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[30]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [14]),
        .O(badr[30]));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[30]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [30]),
        .O(\tr_reg[30] ));
  LUT5 #(
    .INIT(32'hEEE000E0)) 
    \badr[31]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[31]),
        .I3(\badr[31]_INST_0_i_2_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [15]),
        .O(badr[31]));
  LUT6 #(
    .INIT(64'h0F70FFFFFF70FFFF)) 
    \badr[31]_INST_0_i_100 
       (.I0(div_crdy),
        .I1(crdy),
        .I2(ir[7]),
        .I3(ir[8]),
        .I4(ir[10]),
        .I5(ir[6]),
        .O(\badr[31]_INST_0_i_100_n_0 ));
  LUT6 #(
    .INIT(64'h00008A0000000000)) 
    \badr[31]_INST_0_i_101 
       (.I0(ir[9]),
        .I1(ir[8]),
        .I2(ir[7]),
        .I3(ir[2]),
        .I4(ir[6]),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_101_n_0 ));
  LUT6 #(
    .INIT(64'h1340137013701370)) 
    \badr[31]_INST_0_i_102 
       (.I0(ir[6]),
        .I1(ir[9]),
        .I2(ir[7]),
        .I3(ir[8]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\badr[31]_INST_0_i_102_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000007)) 
    \badr[31]_INST_0_i_103 
       (.I0(ir[8]),
        .I1(ir[9]),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(\stat[1]_i_10_0 ),
        .I4(ir[11]),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'h00E000E0EEEE00E0)) 
    \badr[31]_INST_0_i_104 
       (.I0(\badr[31]_INST_0_i_142_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\badr[31]_INST_0_i_143_n_0 ),
        .I3(\badr[31]_INST_0_i_144_n_0 ),
        .I4(ir[11]),
        .I5(\bcmd[3]_INST_0_i_16_n_0 ),
        .O(\badr[31]_INST_0_i_104_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_105 
       (.I0(ir[7]),
        .I1(ir[6]),
        .O(\badr[31]_INST_0_i_105_n_0 ));
  LUT6 #(
    .INIT(64'hEFEFFFFFEF00FFFF)) 
    \badr[31]_INST_0_i_106 
       (.I0(\iv[15]_i_78_n_0 ),
        .I1(\ccmd[3]_INST_0_i_18_n_0 ),
        .I2(\ccmd[1]_INST_0_i_11_n_0 ),
        .I3(\iv[15]_i_84_n_0 ),
        .I4(rst_n_fl_reg_20),
        .I5(\badr[31]_INST_0_i_145_n_0 ),
        .O(\badr[31]_INST_0_i_106_n_0 ));
  LUT6 #(
    .INIT(64'h5400545454005400)) 
    \badr[31]_INST_0_i_107 
       (.I0(\badr[31]_INST_0_i_146_n_0 ),
        .I1(\badr[31]_INST_0_i_147_n_0 ),
        .I2(\sr[13]_i_7_n_0 ),
        .I3(\badr[31]_INST_0_i_148_n_0 ),
        .I4(ir[7]),
        .I5(\ccmd[3]_INST_0_i_10_n_0 ),
        .O(\badr[31]_INST_0_i_107_n_0 ));
  LUT6 #(
    .INIT(64'h00000000CFCC7BCB)) 
    \badr[31]_INST_0_i_108 
       (.I0(ir[3]),
        .I1(ir[6]),
        .I2(ir[4]),
        .I3(ir[7]),
        .I4(ir[5]),
        .I5(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\badr[31]_INST_0_i_108_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00002A000000)) 
    \badr[31]_INST_0_i_109 
       (.I0(ir[7]),
        .I1(div_crdy),
        .I2(crdy),
        .I3(ir[8]),
        .I4(ir[10]),
        .I5(ir[9]),
        .O(\badr[31]_INST_0_i_109_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[31]_INST_0_i_11 
       (.I0(\badr[31]_INST_0_i_29_n_0 ),
        .I1(ctl_sela_rn),
        .O(\badr[31]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFD00FD)) 
    \badr[31]_INST_0_i_110 
       (.I0(\ccmd[4]_INST_0_i_2_n_0 ),
        .I1(\badr[31]_INST_0_i_149_n_0 ),
        .I2(ir[11]),
        .I3(ir[10]),
        .I4(\badr[31]_INST_0_i_150_n_0 ),
        .I5(\badr[31]_INST_0_i_9_n_0 ),
        .O(\badr[31]_INST_0_i_110_n_0 ));
  LUT5 #(
    .INIT(32'h0101F0F5)) 
    \badr[31]_INST_0_i_111 
       (.I0(ir[14]),
        .I1(\sr_reg[13] [7]),
        .I2(ir[15]),
        .I3(\sr_reg[13] [6]),
        .I4(ir[12]),
        .O(\badr[31]_INST_0_i_111_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000AB)) 
    \badr[31]_INST_0_i_113 
       (.I0(\badr[31]_INST_0_i_151_n_0 ),
        .I1(\eir_fl_reg[31]_0 ),
        .I2(\stat[0]_i_8_n_0 ),
        .I3(\badr[31]_INST_0_i_152_n_0 ),
        .I4(\stat[1]_i_16_n_0 ),
        .I5(\tr[31]_i_74_n_0 ),
        .O(\badr[31]_INST_0_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hB0BB0000FFFFFFFF)) 
    \badr[31]_INST_0_i_114 
       (.I0(\badr[31]_INST_0_i_153_n_0 ),
        .I1(\ccmd[3]_INST_0_i_24_n_0 ),
        .I2(\badr[31]_INST_0_i_154_n_0 ),
        .I3(\badr[31]_INST_0_i_99_n_0 ),
        .I4(\badr[31]_INST_0_i_62_n_0 ),
        .I5(\badr[31]_INST_0_i_85_n_0 ),
        .O(\badr[31]_INST_0_i_114_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8AAA8AAAAAAAA)) 
    \badr[31]_INST_0_i_115 
       (.I0(\bdatw[31]_INST_0_i_90_n_0 ),
        .I1(\badr[31]_INST_0_i_98_n_0 ),
        .I2(\badr[31]_INST_0_i_93_n_0 ),
        .I3(ir[5]),
        .I4(\badr[31]_INST_0_i_155_n_0 ),
        .I5(\badr[31]_INST_0_i_156_n_0 ),
        .O(\badr[31]_INST_0_i_115_n_0 ));
  LUT4 #(
    .INIT(16'hAABA)) 
    \badr[31]_INST_0_i_116 
       (.I0(ir[15]),
        .I1(\eir_fl_reg[31]_0 ),
        .I2(\badr[31]_INST_0_i_157_n_0 ),
        .I3(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\badr[31]_INST_0_i_116_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \badr[31]_INST_0_i_117 
       (.I0(ir[5]),
        .I1(ir[7]),
        .I2(ir[4]),
        .O(\badr[31]_INST_0_i_117_n_0 ));
  LUT5 #(
    .INIT(32'hAAAAA2AA)) 
    \badr[31]_INST_0_i_118 
       (.I0(ir[10]),
        .I1(ir[7]),
        .I2(ir[5]),
        .I3(ir[3]),
        .I4(ir[4]),
        .O(\badr[31]_INST_0_i_118_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \badr[31]_INST_0_i_119 
       (.I0(ir[2]),
        .I1(ir[3]),
        .I2(ir[0]),
        .I3(ir[1]),
        .O(\badr[31]_INST_0_i_119_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555555)) 
    \badr[31]_INST_0_i_12 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\badr[31]_INST_0_i_31_n_0 ),
        .I2(ir[15]),
        .I3(\badr[31]_INST_0_i_32_n_0 ),
        .I4(\badr[31]_INST_0_i_33_n_0 ),
        .I5(\badr[31]_INST_0_i_34_n_0 ),
        .O(\badr[31]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h000BFFFF)) 
    \badr[31]_INST_0_i_120 
       (.I0(ir[8]),
        .I1(ir[7]),
        .I2(ir[6]),
        .I3(ir[1]),
        .I4(ir[10]),
        .O(\badr[31]_INST_0_i_120_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \badr[31]_INST_0_i_121 
       (.I0(ir[4]),
        .I1(ir[6]),
        .I2(ir[9]),
        .O(\badr[31]_INST_0_i_121_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_122 
       (.I0(ir[4]),
        .I1(ir[1]),
        .I2(ir[8]),
        .O(\badr[31]_INST_0_i_122_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \badr[31]_INST_0_i_123 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(ir[9]),
        .O(\badr[31]_INST_0_i_123_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_124 
       (.I0(ir[4]),
        .I1(ir[6]),
        .O(\badr[31]_INST_0_i_124_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \badr[31]_INST_0_i_125 
       (.I0(ir[6]),
        .I1(ir[1]),
        .O(\badr[31]_INST_0_i_125_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \badr[31]_INST_0_i_126 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(ir[10]),
        .I3(ir[9]),
        .I4(ir[8]),
        .O(\badr[31]_INST_0_i_126_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_127 
       (.I0(ir[4]),
        .I1(ir[9]),
        .O(\badr[31]_INST_0_i_127_n_0 ));
  LUT5 #(
    .INIT(32'h89EF7FEF)) 
    \badr[31]_INST_0_i_128 
       (.I0(ir[4]),
        .I1(ir[5]),
        .I2(ir[1]),
        .I3(ir[6]),
        .I4(ir[3]),
        .O(\badr[31]_INST_0_i_128_n_0 ));
  LUT5 #(
    .INIT(32'h6F3E7F7F)) 
    \badr[31]_INST_0_i_129 
       (.I0(ir[5]),
        .I1(ir[3]),
        .I2(ir[6]),
        .I3(ir[4]),
        .I4(ir[1]),
        .O(\badr[31]_INST_0_i_129_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_13 
       (.I0(ctl_sela),
        .I1(\badr[31]_INST_0_i_36_n_0 ),
        .O(\badr[31]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[31]_INST_0_i_130 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[8]),
        .O(\badr[31]_INST_0_i_130_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \badr[31]_INST_0_i_131 
       (.I0(ir[9]),
        .I1(ir[8]),
        .I2(ir[1]),
        .I3(ir[7]),
        .I4(ir[4]),
        .O(\badr[31]_INST_0_i_131_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0F470000)) 
    \badr[31]_INST_0_i_132 
       (.I0(ir[1]),
        .I1(ir[8]),
        .I2(ir[4]),
        .I3(ir[6]),
        .I4(ir[9]),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_132_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFBF80)) 
    \badr[31]_INST_0_i_133 
       (.I0(ir[1]),
        .I1(ir[7]),
        .I2(ir[6]),
        .I3(ir[4]),
        .I4(ir[9]),
        .I5(ir[8]),
        .O(\badr[31]_INST_0_i_133_n_0 ));
  LUT6 #(
    .INIT(64'h31233B7320337F33)) 
    \badr[31]_INST_0_i_134 
       (.I0(ir[9]),
        .I1(ir[3]),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(ir[0]),
        .I5(ir[7]),
        .O(\badr[31]_INST_0_i_134_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \badr[31]_INST_0_i_135 
       (.I0(ir[9]),
        .I1(ir[3]),
        .O(\badr[31]_INST_0_i_135_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[31]_INST_0_i_136 
       (.I0(ir[11]),
        .I1(ir[10]),
        .O(\badr[31]_INST_0_i_136_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF7FF)) 
    \badr[31]_INST_0_i_137 
       (.I0(ir[0]),
        .I1(ir[8]),
        .I2(ir[6]),
        .I3(ir[9]),
        .I4(ir[10]),
        .O(\badr[31]_INST_0_i_137_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFBFFF)) 
    \badr[31]_INST_0_i_138 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[3]),
        .I3(ir[0]),
        .I4(ir[5]),
        .I5(ir[4]),
        .O(\badr[31]_INST_0_i_138_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \badr[31]_INST_0_i_139 
       (.I0(ir[10]),
        .I1(ir[8]),
        .I2(ir[9]),
        .O(\badr[31]_INST_0_i_139_n_0 ));
  LUT4 #(
    .INIT(16'h008A)) 
    \badr[31]_INST_0_i_140 
       (.I0(ir[0]),
        .I1(ir[8]),
        .I2(ir[7]),
        .I3(ir[6]),
        .O(\badr[31]_INST_0_i_140_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_141 
       (.I0(ir[9]),
        .I1(ir[10]),
        .O(\badr[31]_INST_0_i_141_n_0 ));
  LUT5 #(
    .INIT(32'hFBF6BFF4)) 
    \badr[31]_INST_0_i_142 
       (.I0(ir[3]),
        .I1(ir[6]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[7]),
        .O(\badr[31]_INST_0_i_142_n_0 ));
  LUT6 #(
    .INIT(64'h2300230000002300)) 
    \badr[31]_INST_0_i_143 
       (.I0(ir[8]),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[11]),
        .I4(ir[10]),
        .I5(ir[7]),
        .O(\badr[31]_INST_0_i_143_n_0 ));
  LUT5 #(
    .INIT(32'h8F000000)) 
    \badr[31]_INST_0_i_144 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(ir[7]),
        .I3(ir[8]),
        .I4(ir[10]),
        .O(\badr[31]_INST_0_i_144_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \badr[31]_INST_0_i_145 
       (.I0(ir[7]),
        .I1(ir[8]),
        .I2(ir[10]),
        .O(\badr[31]_INST_0_i_145_n_0 ));
  LUT5 #(
    .INIT(32'hD7D7FFEB)) 
    \badr[31]_INST_0_i_146 
       (.I0(ir[4]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(ir[3]),
        .I3(ir[6]),
        .I4(ir[5]),
        .O(\badr[31]_INST_0_i_146_n_0 ));
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \badr[31]_INST_0_i_147 
       (.I0(ir[12]),
        .I1(ir[13]),
        .I2(ir[14]),
        .I3(ir[9]),
        .I4(ir[8]),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_147_n_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    \badr[31]_INST_0_i_148 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[11]),
        .O(\badr[31]_INST_0_i_148_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \badr[31]_INST_0_i_149 
       (.I0(ir[13]),
        .I1(ir[12]),
        .I2(ir[15]),
        .I3(ir[14]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\badr[31]_INST_0_i_149_n_0 ));
  LUT6 #(
    .INIT(64'h000F0F0F07070000)) 
    \badr[31]_INST_0_i_150 
       (.I0(div_crdy),
        .I1(crdy),
        .I2(ir[9]),
        .I3(ir[6]),
        .I4(ir[7]),
        .I5(ir[8]),
        .O(\badr[31]_INST_0_i_150_n_0 ));
  LUT4 #(
    .INIT(16'h9DEA)) 
    \badr[31]_INST_0_i_151 
       (.I0(ir[1]),
        .I1(ir[0]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(ir[3]),
        .O(\badr[31]_INST_0_i_151_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \badr[31]_INST_0_i_152 
       (.I0(ir[2]),
        .I1(ir[14]),
        .I2(ir[12]),
        .I3(ir[15]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(ir[1]),
        .O(\badr[31]_INST_0_i_152_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_153 
       (.I0(ir[5]),
        .I1(ir[2]),
        .I2(ir[6]),
        .O(\badr[31]_INST_0_i_153_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_154 
       (.I0(ir[5]),
        .I1(ir[2]),
        .I2(ir[8]),
        .O(\badr[31]_INST_0_i_154_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF808A00F0FFFF)) 
    \badr[31]_INST_0_i_155 
       (.I0(ir[7]),
        .I1(\stat[1]_i_10_0 ),
        .I2(ir[8]),
        .I3(ir[6]),
        .I4(ir[9]),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_155_n_0 ));
  LUT6 #(
    .INIT(64'hFF7F7F7FFFFF7FFF)) 
    \badr[31]_INST_0_i_156 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[8]),
        .I3(ir[7]),
        .I4(\badr[31]_INST_0_i_158_n_0 ),
        .I5(\badr[31]_INST_0_i_159_n_0 ),
        .O(\badr[31]_INST_0_i_156_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \badr[31]_INST_0_i_157 
       (.I0(ir[10]),
        .I1(\tr[31]_i_23_n_0 ),
        .I2(\stat[1]_i_16_n_0 ),
        .I3(ir[9]),
        .I4(ir[8]),
        .I5(ir[7]),
        .O(\badr[31]_INST_0_i_157_n_0 ));
  LUT5 #(
    .INIT(32'hA9BBFCFD)) 
    \badr[31]_INST_0_i_158 
       (.I0(ir[3]),
        .I1(ir[5]),
        .I2(ir[4]),
        .I3(ir[2]),
        .I4(ir[6]),
        .O(\badr[31]_INST_0_i_158_n_0 ));
  LUT5 #(
    .INIT(32'hC00A8CC2)) 
    \badr[31]_INST_0_i_159 
       (.I0(ir[2]),
        .I1(ir[6]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[3]),
        .O(\badr[31]_INST_0_i_159_n_0 ));
  LUT6 #(
    .INIT(64'h0000040000000000)) 
    \badr[31]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_9_n_0 ),
        .I1(ir[13]),
        .I2(ir[11]),
        .I3(ir[10]),
        .I4(\ccmd[4]_INST_0_i_2_n_0 ),
        .I5(\iv_reg[0] ),
        .O(\badr[31]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \badr[31]_INST_0_i_26 
       (.I0(\badr[31]_INST_0_i_12_n_0 ),
        .I1(ctl_sela_rn),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(abus_sel_cr[2]));
  LUT4 #(
    .INIT(16'h0008)) 
    \badr[31]_INST_0_i_28 
       (.I0(\badr[31]_INST_0_i_12_n_0 ),
        .I1(ctl_sela_rn),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(\badr[31]_INST_0_i_13_n_0 ),
        .O(abus_sel_cr[3]));
  LUT6 #(
    .INIT(64'h4444444454555454)) 
    \badr[31]_INST_0_i_29 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\badr[31]_INST_0_i_48_n_0 ),
        .I2(\badr[31]_INST_0_i_49_n_0 ),
        .I3(\badr[31]_INST_0_i_50_n_0 ),
        .I4(\stat[0]_i_12_n_0 ),
        .I5(\badr[31]_INST_0_i_51_n_0 ),
        .O(\badr[31]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'h0400)) 
    \badr[31]_INST_0_i_3 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[31]_INST_0_i_1 [31]),
        .O(\tr_reg[31] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFB00000)) 
    \badr[31]_INST_0_i_30 
       (.I0(\badr[31]_INST_0_i_52_n_0 ),
        .I1(\badr[31]_INST_0_i_53_n_0 ),
        .I2(\badr[31]_INST_0_i_54_n_0 ),
        .I3(\badr[31]_INST_0_i_55_n_0 ),
        .I4(\iv_reg[0] ),
        .I5(\badr[31]_INST_0_i_56_n_0 ),
        .O(ctl_sela_rn));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF100)) 
    \badr[31]_INST_0_i_31 
       (.I0(\badr[31]_INST_0_i_57_n_0 ),
        .I1(\ccmd[1]_INST_0_i_11_n_0 ),
        .I2(\badr[31]_INST_0_i_58_n_0 ),
        .I3(\iv[15]_i_43_n_0 ),
        .I4(\tr[31]_i_9_n_0 ),
        .I5(\badr[31]_INST_0_i_59_n_0 ),
        .O(\badr[31]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \badr[31]_INST_0_i_32 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(ir[10]),
        .I2(\tr[31]_i_23_n_0 ),
        .I3(\tr[31]_i_22_n_0 ),
        .I4(\eir_fl_reg[31]_0 ),
        .O(\badr[31]_INST_0_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hB3F7B3B3FFFFFFFF)) 
    \badr[31]_INST_0_i_33 
       (.I0(ir[11]),
        .I1(ir[12]),
        .I2(\badr[31]_INST_0_i_60_n_0 ),
        .I3(\badr[31]_INST_0_i_61_n_0 ),
        .I4(\badr[31]_INST_0_i_62_n_0 ),
        .I5(\stat[0]_i_12_n_0 ),
        .O(\badr[31]_INST_0_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h55F70000FFFFFFFF)) 
    \badr[31]_INST_0_i_34 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(ir[14]),
        .I3(ctl_fetch_inferred_i_17_n_0),
        .I4(ir[15]),
        .I5(\iv[15]_i_122_0 ),
        .O(\badr[31]_INST_0_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA80808088)) 
    \badr[31]_INST_0_i_35 
       (.I0(\badr[31]_INST_0_i_63_n_0 ),
        .I1(rst_n_fl_reg_20),
        .I2(\badr[31]_INST_0_i_64_n_0 ),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\badr[31]_INST_0_i_65_n_0 ),
        .I5(ir[15]),
        .O(ctl_sela));
  LUT6 #(
    .INIT(64'h4540454045404545)) 
    \badr[31]_INST_0_i_36 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\badr[31]_INST_0_i_66_n_0 ),
        .I2(\badr[31]_INST_0_i_67_n_0 ),
        .I3(\badr[31]_INST_0_i_68_n_0 ),
        .I4(\badr[31]_INST_0_i_69_n_0 ),
        .I5(ir[11]),
        .O(\badr[31]_INST_0_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \badr[31]_INST_0_i_37 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\badr[31]_INST_0_i_70_n_0 ),
        .I2(\badr[31]_INST_0_i_36_n_0 ),
        .I3(ctl_sela),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(abus_sel_0[7]));
  LUT6 #(
    .INIT(64'h0000000000008880)) 
    \badr[31]_INST_0_i_38 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(\stat_reg[2]_12 [2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(abus_sel_0[0]));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \badr[31]_INST_0_i_39 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(ctl_sela_rn),
        .I3(\badr[31]_INST_0_i_29_n_0 ),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\badr[31]_INST_0_i_70_n_0 ),
        .O(abus_sel_0[6]));
  LUT6 #(
    .INIT(64'h0000000000000800)) 
    \badr[31]_INST_0_i_40 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(\badr[31]_INST_0_i_29_n_0 ),
        .I3(ctl_sela_rn),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\badr[31]_INST_0_i_70_n_0 ),
        .O(abus_sel_0[5]));
  LUT6 #(
    .INIT(64'h8880000000000000)) 
    \badr[31]_INST_0_i_41 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(\stat_reg[2]_12 [2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(abus_sel_0[3]));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \badr[31]_INST_0_i_42 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(ctl_sela_rn),
        .I3(\stat_reg[2]_12 [2]),
        .I4(\badr[31]_INST_0_i_70_n_0 ),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(abus_sel_0[4]));
  LUT6 #(
    .INIT(64'h0000000088800000)) 
    \badr[31]_INST_0_i_43 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(\stat_reg[2]_12 [2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(\badr[31]_INST_0_i_29_n_0 ),
        .I5(ctl_sela_rn),
        .O(abus_sel_0[2]));
  LUT6 #(
    .INIT(64'h0000000088800000)) 
    \badr[31]_INST_0_i_44 
       (.I0(\badr[31]_INST_0_i_36_n_0 ),
        .I1(ctl_sela),
        .I2(\stat_reg[2]_12 [2]),
        .I3(\badr[31]_INST_0_i_70_n_0 ),
        .I4(ctl_sela_rn),
        .I5(\badr[31]_INST_0_i_29_n_0 ),
        .O(abus_sel_0[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFF100FFFF)) 
    \badr[31]_INST_0_i_48 
       (.I0(\badr[31]_INST_0_i_71_n_0 ),
        .I1(\stat[0]_i_23_n_0 ),
        .I2(\badr[31]_INST_0_i_72_n_0 ),
        .I3(\iv[15]_i_43_n_0 ),
        .I4(\tr[31]_i_26_n_0 ),
        .I5(\badr[31]_INST_0_i_73_n_0 ),
        .O(\badr[31]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hBABAAABABAAABAAA)) 
    \badr[31]_INST_0_i_49 
       (.I0(ir[15]),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .I2(\stat[0]_i_10_n_0 ),
        .I3(ir[1]),
        .I4(ir[0]),
        .I5(ir[3]),
        .O(\badr[31]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h00F0FFFF2222FFFF)) 
    \badr[31]_INST_0_i_50 
       (.I0(\badr[31]_INST_0_i_74_n_0 ),
        .I1(\badr[31]_INST_0_i_75_n_0 ),
        .I2(\badr[31]_INST_0_i_76_n_0 ),
        .I3(\badr[31]_INST_0_i_77_n_0 ),
        .I4(ir[12]),
        .I5(ir[11]),
        .O(\badr[31]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h55F70000FFFFFFFF)) 
    \badr[31]_INST_0_i_51 
       (.I0(ir[9]),
        .I1(ir[11]),
        .I2(ir[14]),
        .I3(ctl_fetch_inferred_i_17_n_0),
        .I4(ir[15]),
        .I5(\iv[15]_i_122_0 ),
        .O(\badr[31]_INST_0_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h8088808080888088)) 
    \badr[31]_INST_0_i_52 
       (.I0(ir[11]),
        .I1(ir[12]),
        .I2(\badr[31]_INST_0_i_78_n_0 ),
        .I3(\bcmd[3]_INST_0_i_16_n_0 ),
        .I4(\badr[31]_INST_0_i_79_n_0 ),
        .I5(\badr[31]_INST_0_i_80_n_0 ),
        .O(\badr[31]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h00000B00FFFFFFFF)) 
    \badr[31]_INST_0_i_53 
       (.I0(\badr[31]_INST_0_i_81_n_0 ),
        .I1(\ccmd[3]_INST_0_i_24_n_0 ),
        .I2(\badr[31]_INST_0_i_82_n_0 ),
        .I3(\badr[31]_INST_0_i_83_n_0 ),
        .I4(\badr[31]_INST_0_i_84_n_0 ),
        .I5(\badr[31]_INST_0_i_85_n_0 ),
        .O(\badr[31]_INST_0_i_53_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \badr[31]_INST_0_i_54 
       (.I0(ir[14]),
        .I1(ir[13]),
        .I2(ir[15]),
        .O(\badr[31]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'hAEAEAEAEFFAEAEAE)) 
    \badr[31]_INST_0_i_55 
       (.I0(\tr[31]_i_30_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(\badr[31]_INST_0_i_86_n_0 ),
        .I3(ir[15]),
        .I4(ir[8]),
        .I5(\badr[31]_INST_0_i_87_n_0 ),
        .O(\badr[31]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455545554)) 
    \badr[31]_INST_0_i_56 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\badr[31]_INST_0_i_88_n_0 ),
        .I2(\tr[31]_i_9_n_0 ),
        .I3(\badr[31]_INST_0_i_89_n_0 ),
        .I4(\iv[15]_i_43_n_0 ),
        .I5(\badr[31]_INST_0_i_90_n_0 ),
        .O(\badr[31]_INST_0_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFD7FFF)) 
    \badr[31]_INST_0_i_57 
       (.I0(\badr[31]_INST_0_i_91_n_0 ),
        .I1(ir[6]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[7]),
        .I5(\badr[31]_INST_0_i_92_n_0 ),
        .O(\badr[31]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'h888B88888B8B8B8B)) 
    \badr[31]_INST_0_i_58 
       (.I0(\badr[31]_INST_0_i_93_n_0 ),
        .I1(ir[11]),
        .I2(\bcmd[3]_INST_0_i_16_n_0 ),
        .I3(ir[6]),
        .I4(ir[2]),
        .I5(\bcmd[1]_INST_0_i_5_n_0 ),
        .O(\badr[31]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \badr[31]_INST_0_i_59 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(ir[10]),
        .I2(\tr[31]_i_22_n_0 ),
        .I3(\badr[31]_INST_0_i_94_n_0 ),
        .I4(ir[15]),
        .I5(\iv_reg[0]_0 ),
        .O(\badr[31]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000F2)) 
    \badr[31]_INST_0_i_60 
       (.I0(\badr[31]_INST_0_i_95_n_0 ),
        .I1(\badr[31]_INST_0_i_96_n_0 ),
        .I2(\bcmd[3]_INST_0_i_16_n_0 ),
        .I3(\badr[31]_INST_0_i_97_n_0 ),
        .I4(\badr[31]_INST_0_i_93_n_0 ),
        .I5(\badr[31]_INST_0_i_98_n_0 ),
        .O(\badr[31]_INST_0_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hFF40F8F0C840C840)) 
    \badr[31]_INST_0_i_61 
       (.I0(ir[6]),
        .I1(\ccmd[3]_INST_0_i_24_n_0 ),
        .I2(ir[5]),
        .I3(ir[2]),
        .I4(ir[8]),
        .I5(\badr[31]_INST_0_i_99_n_0 ),
        .O(\badr[31]_INST_0_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h000000003AFFFAFF)) 
    \badr[31]_INST_0_i_62 
       (.I0(\badr[31]_INST_0_i_100_n_0 ),
        .I1(ir[10]),
        .I2(ir[9]),
        .I3(ir[5]),
        .I4(ir[6]),
        .I5(\badr[31]_INST_0_i_101_n_0 ),
        .O(\badr[31]_INST_0_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hBAFBFFBFAAAAAAAA)) 
    \badr[31]_INST_0_i_63 
       (.I0(\bcmd[0] ),
        .I1(ir[14]),
        .I2(ir[11]),
        .I3(ir[13]),
        .I4(ir[12]),
        .I5(\iv_reg[0] ),
        .O(\badr[31]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \badr[31]_INST_0_i_64 
       (.I0(\ccmd[3]_INST_0_i_18_n_0 ),
        .I1(\bcmd[0]_INST_0_i_6_n_0 ),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(\iv[15]_i_78_n_0 ),
        .I4(\ccmd[0]_INST_0_i_9_n_0 ),
        .I5(\stat_reg[2]_12 [0]),
        .O(\badr[31]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hF000F2F3F0F0F2F3)) 
    \badr[31]_INST_0_i_65 
       (.I0(\badr[31]_INST_0_i_102_n_0 ),
        .I1(\badr[31]_INST_0_i_103_n_0 ),
        .I2(\badr[31]_INST_0_i_104_n_0 ),
        .I3(ir[10]),
        .I4(ir[11]),
        .I5(\badr[31]_INST_0_i_105_n_0 ),
        .O(\badr[31]_INST_0_i_65_n_0 ));
  LUT5 #(
    .INIT(32'h00000080)) 
    \badr[31]_INST_0_i_66 
       (.I0(\ccmd[2]_INST_0_i_15_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(ir[0]),
        .I3(ir[11]),
        .I4(ir[8]),
        .O(\badr[31]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hAA08080808080808)) 
    \badr[31]_INST_0_i_67 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\badr[31]_INST_0_i_106_n_0 ),
        .I2(\badr[31]_INST_0_i_107_n_0 ),
        .I3(\ccmd[3]_INST_0_i_9_n_0 ),
        .I4(ir[0]),
        .I5(ir[3]),
        .O(\badr[31]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h8AAA8A8A8AAA8AAA)) 
    \badr[31]_INST_0_i_68 
       (.I0(\ccmd[3]_INST_0_i_19_n_0 ),
        .I1(\bdatw[15]_INST_0_i_12_n_0 ),
        .I2(\stat_reg[2]_13 ),
        .I3(\ccmd[4]_INST_0_i_4_n_0 ),
        .I4(\badr[31]_INST_0_i_108_n_0 ),
        .I5(\badr[31]_INST_0_i_109_n_0 ),
        .O(\badr[31]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hFF22FF220000FFF0)) 
    \badr[31]_INST_0_i_69 
       (.I0(\badr[31]_INST_0_i_110_n_0 ),
        .I1(\badr[31]_INST_0_i_111_n_0 ),
        .I2(\badr[31]_INST_0_i_36_0 ),
        .I3(\stat_reg[2]_12 [1]),
        .I4(\badr[31]_INST_0_i_113_n_0 ),
        .I5(ir[13]),
        .O(\badr[31]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00000000AAAABBFB)) 
    \badr[31]_INST_0_i_70 
       (.I0(\badr[31]_INST_0_i_34_n_0 ),
        .I1(\stat[0]_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_114_n_0 ),
        .I3(\badr[31]_INST_0_i_115_n_0 ),
        .I4(\badr[31]_INST_0_i_116_n_0 ),
        .I5(\badr[31]_INST_0_i_31_n_0 ),
        .O(\badr[31]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFFFFF700FFFF)) 
    \badr[31]_INST_0_i_71 
       (.I0(ir[3]),
        .I1(ir[10]),
        .I2(\badr[31]_INST_0_i_117_n_0 ),
        .I3(ir[6]),
        .I4(ir[1]),
        .I5(\badr[31]_INST_0_i_118_n_0 ),
        .O(\badr[31]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h0000080000000000)) 
    \badr[31]_INST_0_i_72 
       (.I0(ir[9]),
        .I1(\bcmd[1]_INST_0_i_5_n_0 ),
        .I2(ir[6]),
        .I3(ir[1]),
        .I4(ir[11]),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001101)) 
    \badr[31]_INST_0_i_73 
       (.I0(\ccmd[1]_INST_0_i_1_0 ),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .I2(\badr[31]_INST_0_i_94_n_0 ),
        .I3(\badr[31]_INST_0_i_119_n_0 ),
        .I4(\stat[1]_i_16_n_0 ),
        .I5(\tr[31]_i_74_n_0 ),
        .O(\badr[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEEEEEEE)) 
    \badr[31]_INST_0_i_74 
       (.I0(\badr[31]_INST_0_i_120_n_0 ),
        .I1(\badr[31]_INST_0_i_121_n_0 ),
        .I2(\badr[31]_INST_0_i_122_n_0 ),
        .I3(\badr[31]_INST_0_i_123_n_0 ),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(div_crdy_reg_1),
        .O(\badr[31]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h00E0FFFF00E000E0)) 
    \badr[31]_INST_0_i_75 
       (.I0(\badr[31]_INST_0_i_124_n_0 ),
        .I1(\badr[31]_INST_0_i_125_n_0 ),
        .I2(\badr[31]_INST_0_i_126_n_0 ),
        .I3(rst_n_fl_reg_17),
        .I4(\badr[31]_INST_0_i_100_n_0 ),
        .I5(\badr[31]_INST_0_i_127_n_0 ),
        .O(\badr[31]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF7FF7FFF77FF)) 
    \badr[31]_INST_0_i_76 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[7]),
        .I3(ir[8]),
        .I4(\badr[31]_INST_0_i_128_n_0 ),
        .I5(\badr[31]_INST_0_i_129_n_0 ),
        .O(\badr[31]_INST_0_i_76_n_0 ));
  LUT6 #(
    .INIT(64'h545454FF54545454)) 
    \badr[31]_INST_0_i_77 
       (.I0(\stat[0]_i_34_n_0 ),
        .I1(ir[4]),
        .I2(\badr[31]_INST_0_i_130_n_0 ),
        .I3(\badr[31]_INST_0_i_131_n_0 ),
        .I4(\badr[31]_INST_0_i_132_n_0 ),
        .I5(\badr[31]_INST_0_i_133_n_0 ),
        .O(\badr[31]_INST_0_i_77_n_0 ));
  LUT6 #(
    .INIT(64'h1F1F1F1111111111)) 
    \badr[31]_INST_0_i_78 
       (.I0(\badr[31]_INST_0_i_134_n_0 ),
        .I1(ir[10]),
        .I2(\stat[0]_i_34_n_0 ),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(ir[6]),
        .I5(ir[3]),
        .O(\badr[31]_INST_0_i_78_n_0 ));
  LUT6 #(
    .INIT(64'hA80A0A8000000088)) 
    \badr[31]_INST_0_i_79 
       (.I0(\tr[31]_i_71_n_0 ),
        .I1(ir[0]),
        .I2(ir[3]),
        .I3(ir[4]),
        .I4(ir[5]),
        .I5(ir[6]),
        .O(\badr[31]_INST_0_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hFCFE5677FFFFFFFF)) 
    \badr[31]_INST_0_i_80 
       (.I0(ir[6]),
        .I1(ir[5]),
        .I2(ir[4]),
        .I3(ir[0]),
        .I4(ir[3]),
        .I5(\ccmd[3]_INST_0_i_23_n_0 ),
        .O(\badr[31]_INST_0_i_80_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \badr[31]_INST_0_i_81 
       (.I0(ir[3]),
        .I1(ir[0]),
        .I2(ir[6]),
        .O(\badr[31]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'h5555404400004044)) 
    \badr[31]_INST_0_i_82 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(ir[0]),
        .I2(ir[8]),
        .I3(ir[7]),
        .I4(ir[6]),
        .I5(ir[3]),
        .O(\badr[31]_INST_0_i_82_n_0 ));
  LUT6 #(
    .INIT(64'hFDFDFFFDFDFFFFFF)) 
    \badr[31]_INST_0_i_83 
       (.I0(div_crdy_reg_1),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\badr[31]_INST_0_i_123_n_0 ),
        .I3(ir[8]),
        .I4(ir[0]),
        .I5(ir[3]),
        .O(\badr[31]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h00000000838F0000)) 
    \badr[31]_INST_0_i_84 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[8]),
        .I3(\stat[1]_i_10_0 ),
        .I4(ir[10]),
        .I5(\badr[31]_INST_0_i_135_n_0 ),
        .O(\badr[31]_INST_0_i_84_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[31]_INST_0_i_85 
       (.I0(ir[12]),
        .I1(ir[11]),
        .O(\badr[31]_INST_0_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \badr[31]_INST_0_i_86 
       (.I0(\eir_fl_reg[31]_0 ),
        .I1(ir[7]),
        .I2(\bdatw[31]_INST_0_i_78_n_0 ),
        .I3(\stat[1]_i_16_n_0 ),
        .I4(\tr[31]_i_23_n_0 ),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_86_n_0 ));
  LUT4 #(
    .INIT(16'h8088)) 
    \badr[31]_INST_0_i_87 
       (.I0(ir[12]),
        .I1(ir[13]),
        .I2(ir[14]),
        .I3(ir[11]),
        .O(\badr[31]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h0000310000000000)) 
    \badr[31]_INST_0_i_88 
       (.I0(\badr[31]_INST_0_i_94_n_0 ),
        .I1(\tr[31]_i_22_n_0 ),
        .I2(\tr[31]_i_23_n_0 ),
        .I3(\iv_reg[0]_0 ),
        .I4(\badr[31]_INST_0_i_136_n_0 ),
        .I5(\fch_irq_lev[1]_i_4_n_0 ),
        .O(\badr[31]_INST_0_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \badr[31]_INST_0_i_89 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\ccmd[2]_INST_0_i_8_n_0 ),
        .I2(\iv[15]_i_85_n_0 ),
        .I3(ir[10]),
        .I4(\tr[31]_i_23_n_0 ),
        .I5(\tr[31]_i_22_n_0 ),
        .O(\badr[31]_INST_0_i_89_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \badr[31]_INST_0_i_9 
       (.I0(ir[14]),
        .I1(ir[15]),
        .I2(ir[12]),
        .O(\badr[31]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h757500007575FF00)) 
    \badr[31]_INST_0_i_90 
       (.I0(\badr[31]_INST_0_i_137_n_0 ),
        .I1(\badr[31]_INST_0_i_138_n_0 ),
        .I2(\badr[31]_INST_0_i_139_n_0 ),
        .I3(\badr[31]_INST_0_i_140_n_0 ),
        .I4(ir[11]),
        .I5(\bcmd[3]_INST_0_i_16_n_0 ),
        .O(\badr[31]_INST_0_i_90_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \badr[31]_INST_0_i_91 
       (.I0(ir[2]),
        .I1(ir[3]),
        .I2(ir[8]),
        .I3(ir[9]),
        .O(\badr[31]_INST_0_i_91_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \badr[31]_INST_0_i_92 
       (.I0(ir[9]),
        .I1(ir[7]),
        .I2(ir[8]),
        .O(\badr[31]_INST_0_i_92_n_0 ));
  LUT5 #(
    .INIT(32'h00000800)) 
    \badr[31]_INST_0_i_93 
       (.I0(ir[2]),
        .I1(ir[8]),
        .I2(ir[6]),
        .I3(ir[9]),
        .I4(ir[10]),
        .O(\badr[31]_INST_0_i_93_n_0 ));
  LUT4 #(
    .INIT(16'hFFFB)) 
    \badr[31]_INST_0_i_94 
       (.I0(ir[2]),
        .I1(ir[3]),
        .I2(ir[0]),
        .I3(ir[1]),
        .O(\badr[31]_INST_0_i_94_n_0 ));
  LUT6 #(
    .INIT(64'h5DD7FFF57DDFFFFF)) 
    \badr[31]_INST_0_i_95 
       (.I0(\tr[31]_i_71_n_0 ),
        .I1(ir[3]),
        .I2(ir[4]),
        .I3(ir[5]),
        .I4(ir[6]),
        .I5(ir[2]),
        .O(\badr[31]_INST_0_i_95_n_0 ));
  LUT6 #(
    .INIT(64'h000000A288888020)) 
    \badr[31]_INST_0_i_96 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(ir[6]),
        .I2(ir[2]),
        .I3(ir[4]),
        .I4(ir[5]),
        .I5(ir[3]),
        .O(\badr[31]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h8088AAA88088AAAA)) 
    \badr[31]_INST_0_i_97 
       (.I0(ir[5]),
        .I1(\badr[31]_INST_0_i_141_n_0 ),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(\stat[0]_i_34_n_0 ),
        .I5(ir[7]),
        .O(\badr[31]_INST_0_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DD88EC4C)) 
    \badr[31]_INST_0_i_98 
       (.I0(ir[7]),
        .I1(ir[5]),
        .I2(ir[6]),
        .I3(ir[2]),
        .I4(ir[8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\badr[31]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \badr[31]_INST_0_i_99 
       (.I0(ir[11]),
        .I1(ir[9]),
        .I2(\ccmd[4]_INST_0_i_4_n_0 ),
        .I3(crdy),
        .I4(div_crdy),
        .I5(ir[10]),
        .O(\badr[31]_INST_0_i_99_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[3]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[3]),
        .O(badr[3]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[3]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [3]),
        .I5(\mul_a_reg[15] [3]),
        .O(\tr_reg[3] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[4]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[4]),
        .O(badr[4]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[4]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [4]),
        .I5(\mul_a_reg[15] [4]),
        .O(\tr_reg[4] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[5]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[5]),
        .O(badr[5]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[5]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [5]),
        .I5(\mul_a_reg[15] [5]),
        .O(\tr_reg[5] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[6]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[6]),
        .O(badr[6]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[6]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [6]),
        .I5(\mul_a_reg[15] [6]),
        .O(\tr_reg[6] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[7]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[7]),
        .O(badr[7]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[7]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [7]),
        .I5(\mul_a_reg[15] [7]),
        .O(\tr_reg[7] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[8]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[8]),
        .O(badr[8]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[8]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [8]),
        .I5(\mul_a_reg[15] [8]),
        .O(\tr_reg[8] ));
  LUT3 #(
    .INIT(8'hE0)) 
    \badr[9]_INST_0 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[9]),
        .O(badr[9]));
  LUT6 #(
    .INIT(64'h0407000304040000)) 
    \badr[9]_INST_0_i_2 
       (.I0(\badr[31]_INST_0_i_11_n_0 ),
        .I1(\badr[31]_INST_0_i_12_n_0 ),
        .I2(\badr[31]_INST_0_i_13_n_0 ),
        .I3(\badr[15]_INST_0_i_7_n_0 ),
        .I4(\badr[31]_INST_0_i_1 [9]),
        .I5(\mul_a_reg[15] [9]),
        .O(\tr_reg[9] ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[0]_i_1 
       (.I0(cbus[16]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[0]),
        .O(\sr_reg[8]_72 [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[10]_i_1 
       (.I0(cbus[23]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[10]),
        .O(\sr_reg[8]_72 [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[14]_i_1 
       (.I0(cbus[24]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[14]),
        .O(\sr_reg[8]_72 [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[1]_i_1 
       (.I0(cbus[17]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[1]),
        .O(\sr_reg[8]_72 [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[2]_i_1 
       (.I0(cbus[18]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[2]),
        .O(\sr_reg[8]_72 [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[4]_i_1 
       (.I0(cbus[19]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[4]),
        .O(\sr_reg[8]_72 [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[6]_i_1 
       (.I0(cbus[20]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[6]),
        .O(\sr_reg[8]_72 [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[8]_i_1 
       (.I0(cbus[21]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[8]),
        .O(\sr_reg[8]_72 [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[9]_i_1 
       (.I0(cbus[22]),
        .I1(\sr_reg[13] [8]),
        .I2(cbus[9]),
        .O(\sr_reg[8]_72 [6]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[10]_INST_0 
       (.I0(bbus_0[8]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[11]_INST_0 
       (.I0(bbus_0[9]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[12]_INST_0 
       (.I0(bbus_0[10]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[13]_INST_0 
       (.I0(bbus_0[11]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[14]_INST_0 
       (.I0(bbus_0[12]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[15]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[13]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[16]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_14),
        .O(bbus_o[14]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[17]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_13),
        .O(bbus_o[15]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[18]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_12),
        .O(bbus_o[16]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[19]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_11),
        .O(bbus_o[17]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[1]_INST_0 
       (.I0(bbus_0[0]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[20]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_10),
        .O(bbus_o[18]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[21]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_9),
        .O(bbus_o[19]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[22]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_8),
        .O(bbus_o[20]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[23]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_7),
        .O(bbus_o[21]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[24]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_6),
        .O(bbus_o[22]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[25]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_16),
        .O(bbus_o[23]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[26]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_5),
        .O(bbus_o[24]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[27]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_4),
        .O(bbus_o[25]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[28]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_3),
        .O(bbus_o[26]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[29]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_2),
        .O(bbus_o[27]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[2]_INST_0 
       (.I0(bbus_0[1]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[30]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_1),
        .O(bbus_o[28]));
  LUT2 #(
    .INIT(4'h2)) 
    \bbus_o[31]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(rst_n_fl_reg_0),
        .O(bbus_o[29]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[3]_INST_0 
       (.I0(bbus_0[2]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[4]_INST_0 
       (.I0(bbus_0[3]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[6]_INST_0 
       (.I0(bbus_0[4]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[7]_INST_0 
       (.I0(bbus_0[5]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[8]_INST_0 
       (.I0(bbus_0[6]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[9]_INST_0 
       (.I0(bbus_0[7]),
        .I1(\stat_reg[0]_3 ),
        .O(bbus_o[7]));
  LUT6 #(
    .INIT(64'h00000000BABABABB)) 
    \bcmd[0]_INST_0 
       (.I0(\bcmd[0]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_2_n_0 ),
        .I2(\bcmd[0]_INST_0_i_3_n_0 ),
        .I3(\stat_reg[2]_12 [0]),
        .I4(ir[7]),
        .I5(\bcmd[0]_INST_0_i_4_n_0 ),
        .O(\stat_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h11FF111011101110)) 
    \bcmd[0]_INST_0_i_1 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(\bcmd[0]_INST_0_i_5_n_0 ),
        .I3(\bcmd[0]_INST_0_i_6_n_0 ),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(\bcmd[0]_INST_0_i_8_n_0 ),
        .O(\bcmd[0]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hBB2F)) 
    \bcmd[0]_INST_0_i_11 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(ir[0]),
        .I2(ir[1]),
        .I3(ir[3]),
        .O(\bcmd[0]_INST_0_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[0]_INST_0_i_12 
       (.I0(ir[4]),
        .I1(ir[5]),
        .O(\bcmd[0]_INST_0_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hBF)) 
    \bcmd[0]_INST_0_i_2 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(ir[9]),
        .O(\bcmd[0]_INST_0_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0800)) 
    \bcmd[0]_INST_0_i_3 
       (.I0(ir[7]),
        .I1(rst_n_fl_reg_17),
        .I2(ir[8]),
        .I3(\stat_reg[2]_12 [0]),
        .O(\bcmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hBFABFFFFFFFEFFFF)) 
    \bcmd[0]_INST_0_i_4 
       (.I0(\bcmd[0]_INST_0_i_9_n_0 ),
        .I1(ir[11]),
        .I2(ir[10]),
        .I3(ir[6]),
        .I4(\bcmd[0] ),
        .I5(ir[12]),
        .O(\bcmd[0]_INST_0_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h9A000000)) 
    \bcmd[0]_INST_0_i_5 
       (.I0(ir[5]),
        .I1(ir[7]),
        .I2(ir[4]),
        .I3(ir[3]),
        .I4(ir[6]),
        .O(\bcmd[0]_INST_0_i_5_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[0]_INST_0_i_6 
       (.I0(ir[11]),
        .I1(ir[10]),
        .O(\bcmd[0]_INST_0_i_6_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_7 
       (.I0(ir[6]),
        .I1(ir[8]),
        .I2(ir[9]),
        .O(\bcmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF00000400000004)) 
    \bcmd[0]_INST_0_i_8 
       (.I0(\bcmd[0]_INST_0_i_11_n_0 ),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(ir[2]),
        .I3(ir[10]),
        .I4(ir[7]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\bcmd[0]_INST_0_i_8_n_0 ));
  LUT3 #(
    .INIT(8'h7E)) 
    \bcmd[0]_INST_0_i_9 
       (.I0(ir[12]),
        .I1(ir[13]),
        .I2(ir[14]),
        .O(\bcmd[0]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h5454545454555454)) 
    \bcmd[1]_INST_0 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[1]_INST_0_i_2_n_0 ),
        .I2(\bcmd[1]_INST_0_i_3_n_0 ),
        .I3(\bcmd[1]_INST_0_i_4_n_0 ),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(ir[11]),
        .O(\stat_reg[2]_6 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bcmd[1]_INST_0_i_1 
       (.I0(ir[15]),
        .I1(\stat_reg[2]_12 [2]),
        .O(\bcmd[1]_INST_0_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \bcmd[1]_INST_0_i_10 
       (.I0(ir[13]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(ir[14]),
        .I3(ir[12]),
        .O(\bcmd[1]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000000B05000000)) 
    \bcmd[1]_INST_0_i_11 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\eir_fl_reg[31]_0 ),
        .I2(\bcmd[1]_INST_0_i_15_n_0 ),
        .I3(\stat_reg[2]_12 [1]),
        .I4(ir[3]),
        .I5(ir[0]),
        .O(\bcmd[1]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \bcmd[1]_INST_0_i_12 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[3]),
        .I3(ir[6]),
        .O(\bcmd[1]_INST_0_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[1]_INST_0_i_13 
       (.I0(ir[6]),
        .I1(ir[8]),
        .I2(ir[9]),
        .O(\bcmd[1]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \bcmd[1]_INST_0_i_15 
       (.I0(ir[8]),
        .I1(ir[10]),
        .I2(ir[9]),
        .I3(ir[1]),
        .I4(\bcmd[1]_INST_0_i_16_n_0 ),
        .I5(\bcmd[3]_INST_0_i_2_n_0 ),
        .O(\bcmd[1]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \bcmd[1]_INST_0_i_16 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[2]),
        .I3(ir[6]),
        .O(\bcmd[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \bcmd[1]_INST_0_i_2 
       (.I0(ir[11]),
        .I1(rst_n_fl_reg_17),
        .I2(\iv_reg[0]_1 ),
        .I3(ir[6]),
        .I4(ir[9]),
        .I5(\bcmd[1]_INST_0_i_7_n_0 ),
        .O(\bcmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h000000E000E00000)) 
    \bcmd[1]_INST_0_i_3 
       (.I0(\bcmd[1]_INST_0_i_8_n_0 ),
        .I1(\bcmd[1]_INST_0_i_9_n_0 ),
        .I2(ir[11]),
        .I3(\bcmd[1]_INST_0_i_10_n_0 ),
        .I4(\stat_reg[2]_12 [0]),
        .I5(ir[9]),
        .O(\bcmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFFF7FF)) 
    \bcmd[1]_INST_0_i_4 
       (.I0(ir[6]),
        .I1(ir[9]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[10]),
        .I4(\bcmd[1]_INST_0_i_10_n_0 ),
        .I5(\bcmd[1]_INST_0_i_11_n_0 ),
        .O(\bcmd[1]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bcmd[1]_INST_0_i_5 
       (.I0(ir[8]),
        .I1(ir[7]),
        .O(\bcmd[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \bcmd[1]_INST_0_i_7 
       (.I0(ir[12]),
        .I1(ir[13]),
        .I2(ir[14]),
        .I3(ir[10]),
        .I4(ir[8]),
        .I5(ir[7]),
        .O(\bcmd[1]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hC000202000000000)) 
    \bcmd[1]_INST_0_i_8 
       (.I0(ir[6]),
        .I1(ir[9]),
        .I2(ir[10]),
        .I3(\bcmd[1]_INST_0_i_12_n_0 ),
        .I4(ir[8]),
        .I5(ir[7]),
        .O(\bcmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h20208220AAAAAAAA)) 
    \bcmd[1]_INST_0_i_9 
       (.I0(\bcmd[1]_INST_0_i_13_n_0 ),
        .I1(ir[3]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[7]),
        .I5(ir[10]),
        .O(\bcmd[1]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000100010000000)) 
    \bcmd[2]_INST_0 
       (.I0(\bcmd[2] ),
        .I1(ir[7]),
        .I2(ir[8]),
        .I3(ir[9]),
        .I4(ir[11]),
        .I5(ir[10]),
        .O(\stat_reg[1] ));
  LUT3 #(
    .INIT(8'h80)) 
    \bcmd[2]_INST_0_i_2 
       (.I0(ir[14]),
        .I1(ir[13]),
        .I2(ir[12]),
        .O(rst_n_fl_reg_20));
  LUT6 #(
    .INIT(64'h000000000000AAEA)) 
    \bcmd[3]_INST_0 
       (.I0(\bcmd[3]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_2_n_0 ),
        .I2(\bcmd[3] ),
        .I3(\bcmd[3]_INST_0_i_4_n_0 ),
        .I4(\bcmd[3]_INST_0_i_5_n_0 ),
        .I5(\bcmd[3]_INST_0_i_6_n_0 ),
        .O(\stat_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h000000005444DCCC)) 
    \bcmd[3]_INST_0_i_1 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(rst_n_fl_reg_17),
        .I2(crdy),
        .I3(div_crdy),
        .I4(ir[11]),
        .I5(\bcmd[3]_INST_0_i_8_n_0 ),
        .O(\bcmd[3]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[3]_INST_0_i_10 
       (.I0(ir[0]),
        .I1(\stat_reg[2]_12 [1]),
        .O(\bcmd[3]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF40)) 
    \bcmd[3]_INST_0_i_11 
       (.I0(\bcmd[3]_INST_0_i_14_n_0 ),
        .I1(\bcmd[3]_INST_0_i_15_n_0 ),
        .I2(ir[8]),
        .I3(\bcmd[3]_INST_0_i_16_n_0 ),
        .I4(\stat_reg[2]_12 [0]),
        .I5(ir[7]),
        .O(\bcmd[3]_INST_0_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00000001)) 
    \bcmd[3]_INST_0_i_12 
       (.I0(ir[7]),
        .I1(ir[10]),
        .I2(ir[4]),
        .I3(ir[5]),
        .I4(ir[2]),
        .O(\bcmd[3]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[3]_INST_0_i_13 
       (.I0(ir[1]),
        .I1(ir[0]),
        .O(\bcmd[3]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bcmd[3]_INST_0_i_14 
       (.I0(ir[4]),
        .I1(ir[5]),
        .O(\bcmd[3]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[3]_INST_0_i_15 
       (.I0(ir[3]),
        .I1(ir[5]),
        .O(\bcmd[3]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bcmd[3]_INST_0_i_16 
       (.I0(ir[9]),
        .I1(ir[10]),
        .O(\bcmd[3]_INST_0_i_16_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[3]_INST_0_i_2 
       (.I0(ir[12]),
        .I1(ir[13]),
        .I2(ir[14]),
        .O(\bcmd[3]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \bcmd[3]_INST_0_i_4 
       (.I0(ir[8]),
        .I1(ir[10]),
        .I2(ir[11]),
        .O(\bcmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAABAA)) 
    \bcmd[3]_INST_0_i_5 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\bcmd[3]_INST_0_i_9_n_0 ),
        .I2(ir[2]),
        .I3(ir[3]),
        .I4(\bcmd[3]_INST_0_i_10_n_0 ),
        .I5(ir[5]),
        .O(\bcmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h2A002AAA2AAA2AAA)) 
    \bcmd[3]_INST_0_i_6 
       (.I0(\bcmd[3]_INST_0_i_11_n_0 ),
        .I1(ir[7]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[9]),
        .I4(\bcmd[3]_INST_0_i_12_n_0 ),
        .I5(ir[3]),
        .O(\bcmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEFFFFFFFFFFF)) 
    \bcmd[3]_INST_0_i_7 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(ir[13]),
        .I3(ir[12]),
        .I4(ir[15]),
        .I5(ir[14]),
        .O(rst_n_fl_reg_17));
  LUT5 #(
    .INIT(32'hBFFBFFFB)) 
    \bcmd[3]_INST_0_i_8 
       (.I0(\bcmd[1]_INST_0_i_10_n_0 ),
        .I1(ir[10]),
        .I2(ir[8]),
        .I3(ir[11]),
        .I4(ir[6]),
        .O(\bcmd[3]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bcmd[3]_INST_0_i_9 
       (.I0(ir[7]),
        .I1(ir[4]),
        .I2(ir[9]),
        .I3(ir[6]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\bcmd[3]_INST_0_i_13_n_0 ),
        .O(\bcmd[3]_INST_0_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[0]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(\bdatw[5] [0]),
        .O(bdatw[0]));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[10]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(bbus_0[1]),
        .I4(bbus_0[8]),
        .O(bdatw[10]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAE)) 
    \bdatw[10]_INST_0_i_1 
       (.I0(\bdatw[10]_INST_0_i_3_n_0 ),
        .I1(eir[2]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\mul_b_reg[2] ),
        .I4(\mul_b_reg[2]_0 ),
        .I5(\mul_b_reg[2]_1 ),
        .O(bbus_0[1]));
  LUT4 #(
    .INIT(16'h0100)) 
    \bdatw[10]_INST_0_i_10 
       (.I0(ir[2]),
        .I1(ir[3]),
        .I2(ir[0]),
        .I3(ir[1]),
        .O(\bdatw[10]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[10]_INST_0_i_2 
       (.I0(\bdatw[10]_INST_0_i_7_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(eir[10]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\mul_b_reg[10] ),
        .I5(\mul_b_reg[10]_0 ),
        .O(bbus_0[8]));
  LUT6 #(
    .INIT(64'h5505045450000454)) 
    \bdatw[10]_INST_0_i_3 
       (.I0(\sr_reg[6]_2 ),
        .I1(ir[1]),
        .I2(ctl_selb_0),
        .I3(\bdatw[10]_INST_0_i_10_n_0 ),
        .I4(\stat_reg[0]_5 ),
        .I5(ir[2]),
        .O(\bdatw[10]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h9AAAAAAA9AAAFFFF)) 
    \bdatw[10]_INST_0_i_7 
       (.I0(\stat_reg[0]_5 ),
        .I1(ir[2]),
        .I2(ir[3]),
        .I3(\bdatw[14]_INST_0_i_9_n_0 ),
        .I4(ctl_selb_0),
        .I5(ir[9]),
        .O(\bdatw[10]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[11]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(bbus_0[2]),
        .I4(bbus_0[9]),
        .O(bdatw[11]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF2)) 
    \bdatw[11]_INST_0_i_1 
       (.I0(eir[3]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\mul_b_reg[3] ),
        .I3(\mul_b_reg[3]_0 ),
        .I4(\mul_b_reg[3]_1 ),
        .I5(\bdatw[11]_INST_0_i_6_n_0 ),
        .O(bbus_0[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[11]_INST_0_i_19 
       (.I0(ir[3]),
        .I1(ir[2]),
        .O(\bdatw[11]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    \bdatw[11]_INST_0_i_2 
       (.I0(\bdatw[11]_INST_0_i_7_n_0 ),
        .I1(eir[11]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\mul_b_reg[11] ),
        .I4(\mul_b_reg[11]_0 ),
        .O(bbus_0[9]));
  LUT6 #(
    .INIT(64'h1112111132103210)) 
    \bdatw[11]_INST_0_i_6 
       (.I0(\stat_reg[0]_5 ),
        .I1(\sr_reg[6]_2 ),
        .I2(ir[2]),
        .I3(ir[3]),
        .I4(\bdatw[15]_INST_0_i_10_n_0 ),
        .I5(ctl_selb_0),
        .O(\bdatw[11]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000C2323232)) 
    \bdatw[11]_INST_0_i_7 
       (.I0(ir[10]),
        .I1(\stat_reg[0]_5 ),
        .I2(ctl_selb_0),
        .I3(\bdatw[11]_INST_0_i_19_n_0 ),
        .I4(\bdatw[15]_INST_0_i_10_n_0 ),
        .I5(\sr_reg[6]_2 ),
        .O(\bdatw[11]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[12]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(bbus_0[3]),
        .I4(bbus_0[10]),
        .O(bdatw[12]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF2)) 
    \bdatw[12]_INST_0_i_1 
       (.I0(\bdatw[12]_INST_0_i_3_n_0 ),
        .I1(\bdatw[12]_INST_0_i_4_n_0 ),
        .I2(\mul_b_reg[4] ),
        .I3(\mul_b_reg[4]_0 ),
        .I4(\mul_b_reg[4]_1 ),
        .I5(rst_n_fl_reg_15),
        .O(bbus_0[3]));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    \bdatw[12]_INST_0_i_2 
       (.I0(\bdatw[12]_INST_0_i_9_n_0 ),
        .I1(eir[12]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\mul_b_reg[12] ),
        .I4(\mul_b_reg[12]_0 ),
        .O(bbus_0[10]));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[12]_INST_0_i_21 
       (.I0(\stat_reg[0]_5 ),
        .I1(ctl_selb_0),
        .I2(\sr_reg[6]_2 ),
        .I3(ctl_selb_rn[1]),
        .I4(\stat_reg[2]_8 ),
        .I5(ctl_selb_rn[0]),
        .O(bbus_sel_cr[1]));
  LUT4 #(
    .INIT(16'h0010)) 
    \bdatw[12]_INST_0_i_22 
       (.I0(ir[0]),
        .I1(ir[1]),
        .I2(ir[2]),
        .I3(ir[3]),
        .O(\bdatw[12]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[12]_INST_0_i_23 
       (.I0(ir[3]),
        .I1(ir[2]),
        .O(\bdatw[12]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \bdatw[12]_INST_0_i_3 
       (.I0(ir[0]),
        .I1(ir[1]),
        .I2(ir[2]),
        .I3(ir[3]),
        .I4(ctl_selb_0),
        .I5(ir[4]),
        .O(\bdatw[12]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[12]_INST_0_i_4 
       (.I0(\sr_reg[6]_2 ),
        .I1(\stat_reg[0]_5 ),
        .O(\bdatw[12]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4444444444)) 
    \bdatw[12]_INST_0_i_8 
       (.I0(\bdatw[31]_INST_0_i_2_n_0 ),
        .I1(eir[4]),
        .I2(\bdatw[12]_INST_0_i_22_n_0 ),
        .I3(ctl_selb_0),
        .I4(ir[3]),
        .I5(\bdatw[31]_INST_0_i_8_n_0 ),
        .O(rst_n_fl_reg_15));
  LUT6 #(
    .INIT(64'h00000000C2323232)) 
    \bdatw[12]_INST_0_i_9 
       (.I0(ir[10]),
        .I1(\stat_reg[0]_5 ),
        .I2(ctl_selb_0),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\bdatw[12]_INST_0_i_23_n_0 ),
        .I5(\sr_reg[6]_2 ),
        .O(\bdatw[12]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[13]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(\bdatw[5] [1]),
        .I4(bbus_0[11]),
        .O(bdatw[13]));
  LUT4 #(
    .INIT(16'h0040)) 
    \bdatw[13]_INST_0_i_12 
       (.I0(ir[1]),
        .I1(ir[0]),
        .I2(ir[2]),
        .I3(ir[3]),
        .O(\bdatw[13]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[13]_INST_0_i_2 
       (.I0(\bdatw[13]_INST_0_i_9_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(eir[13]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\mul_b_reg[13] ),
        .I5(\mul_b_reg[13]_0 ),
        .O(bbus_0[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[13]_INST_0_i_26 
       (.I0(bbus_sel_cr[0]),
        .I1(\sr_reg[13] [5]),
        .O(bbus_sr[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_27 
       (.I0(ir[0]),
        .I1(ir[1]),
        .O(\bdatw[13]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'h5505045450000454)) 
    \bdatw[13]_INST_0_i_3 
       (.I0(\sr_reg[6]_2 ),
        .I1(ir[4]),
        .I2(ctl_selb_0),
        .I3(\bdatw[13]_INST_0_i_12_n_0 ),
        .I4(\stat_reg[0]_5 ),
        .I5(ir[5]),
        .O(rst_n_fl_reg_23));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[13]_INST_0_i_4 
       (.I0(eir[5]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .O(rst_n_fl_reg_22));
  LUT6 #(
    .INIT(64'hFF0D0000FFFFFFFF)) 
    \bdatw[13]_INST_0_i_67 
       (.I0(\bdatw[31]_INST_0_i_69_n_0 ),
        .I1(\bdatw[31]_INST_0_i_68_n_0 ),
        .I2(\bdatw[31]_INST_0_i_67_n_0 ),
        .I3(\bdatw[31]_INST_0_i_66_n_0 ),
        .I4(\stat_reg[0]_10 ),
        .I5(\stat_reg[2]_8 ),
        .O(\stat_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h6AAAAAAA6AAAFFFF)) 
    \bdatw[13]_INST_0_i_9 
       (.I0(\stat_reg[0]_5 ),
        .I1(ir[2]),
        .I2(ir[3]),
        .I3(\bdatw[13]_INST_0_i_27_n_0 ),
        .I4(ctl_selb_0),
        .I5(ir[10]),
        .O(\bdatw[13]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[14]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(bbus_0[4]),
        .I4(bbus_0[12]),
        .O(bdatw[14]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[14]_INST_0_i_1 
       (.I0(\bdatw[14]_INST_0_i_3_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(eir[6]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\mul_b_reg[6] ),
        .I5(\mul_b_reg[6]_0 ),
        .O(bbus_0[4]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[14]_INST_0_i_2 
       (.I0(\bdatw[14]_INST_0_i_6_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(eir[14]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\mul_b_reg[14] ),
        .I5(\mul_b_reg[14]_0 ),
        .O(bbus_0[12]));
  LUT6 #(
    .INIT(64'hCC3C4444CC3C7777)) 
    \bdatw[14]_INST_0_i_3 
       (.I0(ir[6]),
        .I1(\stat_reg[0]_5 ),
        .I2(\bdatw[14]_INST_0_i_9_n_0 ),
        .I3(\bdatw[15]_INST_0_i_11_n_0 ),
        .I4(ctl_selb_0),
        .I5(ir[5]),
        .O(\bdatw[14]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h6AAAAAAA6AAAFFFF)) 
    \bdatw[14]_INST_0_i_6 
       (.I0(\stat_reg[0]_5 ),
        .I1(ir[2]),
        .I2(ir[3]),
        .I3(\bdatw[14]_INST_0_i_9_n_0 ),
        .I4(ctl_selb_0),
        .I5(ir[10]),
        .O(\bdatw[14]_INST_0_i_6_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[14]_INST_0_i_9 
       (.I0(ir[1]),
        .I1(ir[0]),
        .O(\bdatw[14]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[15]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(bbus_0[5]),
        .I4(bbus_0[13]),
        .O(bdatw[15]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[15]_INST_0_i_1 
       (.I0(\bdatw[15]_INST_0_i_3_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(eir[7]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\mul_b_reg[7] ),
        .I5(\mul_b_reg[7]_0 ),
        .O(bbus_0[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[15]_INST_0_i_10 
       (.I0(ir[1]),
        .I1(ir[0]),
        .O(\bdatw[15]_INST_0_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \bdatw[15]_INST_0_i_11 
       (.I0(ir[3]),
        .I1(ir[2]),
        .O(\bdatw[15]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h2AAA)) 
    \bdatw[15]_INST_0_i_12 
       (.I0(ir[15]),
        .I1(ir[12]),
        .I2(ir[13]),
        .I3(ir[14]),
        .O(\bdatw[15]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055D55555)) 
    \bdatw[15]_INST_0_i_13 
       (.I0(ir[14]),
        .I1(\bcmd[3]_INST_0_i_14_n_0 ),
        .I2(\bdatw[15]_INST_0_i_28_n_0 ),
        .I3(\bcmd[3]_INST_0_i_16_n_0 ),
        .I4(ir[7]),
        .I5(\bdatw[15]_INST_0_i_29_n_0 ),
        .O(\bdatw[15]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h04FF)) 
    \bdatw[15]_INST_0_i_14 
       (.I0(ir[14]),
        .I1(\sr_reg[13] [6]),
        .I2(ir[12]),
        .I3(ir[13]),
        .O(\bdatw[15]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \bdatw[15]_INST_0_i_18 
       (.I0(\stat_reg[0]_5 ),
        .I1(ctl_selb_0),
        .I2(\sr_reg[6]_2 ),
        .I3(ctl_selb_rn[1]),
        .I4(ctl_selb_rn[0]),
        .I5(\stat_reg[2]_8 ),
        .O(bbus_sel_cr[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[15]_INST_0_i_2 
       (.I0(\bdatw[15]_INST_0_i_7_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(eir[15]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\mul_b_reg[15] ),
        .I5(\mul_b_reg[15]_0 ),
        .O(bbus_0[13]));
  LUT6 #(
    .INIT(64'h0000000000000080)) 
    \bdatw[15]_INST_0_i_22 
       (.I0(\stat_reg[0]_5 ),
        .I1(ctl_selb_0),
        .I2(\sr_reg[6]_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_cr[0]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[15]_INST_0_i_28 
       (.I0(ir[8]),
        .I1(ir[6]),
        .O(\bdatw[15]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFBFBEEE)) 
    \bdatw[15]_INST_0_i_29 
       (.I0(ir[15]),
        .I1(ir[11]),
        .I2(ir[12]),
        .I3(\sr_reg[13] [7]),
        .I4(ir[14]),
        .I5(\bdatw[15]_INST_0_i_14_n_0 ),
        .O(\bdatw[15]_INST_0_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hCC3C4444CC3C7777)) 
    \bdatw[15]_INST_0_i_3 
       (.I0(ir[7]),
        .I1(\stat_reg[0]_5 ),
        .I2(\bdatw[15]_INST_0_i_10_n_0 ),
        .I3(\bdatw[15]_INST_0_i_11_n_0 ),
        .I4(ctl_selb_0),
        .I5(ir[6]),
        .O(\bdatw[15]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h01111101FFFFFFFF)) 
    \bdatw[15]_INST_0_i_4 
       (.I0(\bdatw[15]_INST_0_i_12_n_0 ),
        .I1(\bdatw[15]_INST_0_i_13_n_0 ),
        .I2(\bdatw[15]_INST_0_i_14_n_0 ),
        .I3(\mul_b_reg[15]_1 ),
        .I4(ir[11]),
        .I5(\iv_reg[0] ),
        .O(\sr_reg[6]_2 ));
  LUT6 #(
    .INIT(64'hFFFFCCDF00000000)) 
    \bdatw[15]_INST_0_i_61 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[31]_INST_0_i_66_n_0 ),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_70_n_0 ),
        .I5(\stat_reg[0]_10 ),
        .O(\stat_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h3322FFF2FFFFFFFF)) 
    \bdatw[15]_INST_0_i_62 
       (.I0(\bdatw[15]_INST_0_i_70_n_0 ),
        .I1(\bdatw[31]_INST_0_i_66_n_0 ),
        .I2(\bdatw[15]_INST_0_i_71_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_70_n_0 ),
        .I5(\stat_reg[0]_10 ),
        .O(\stat_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h5555FF5DFFFFFFFF)) 
    \bdatw[15]_INST_0_i_68 
       (.I0(\stat_reg[2]_8 ),
        .I1(\bdatw[31]_INST_0_i_69_n_0 ),
        .I2(\bdatw[31]_INST_0_i_68_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_66_n_0 ),
        .I5(\stat_reg[0]_10 ),
        .O(\stat_reg[2]_10 ));
  LUT6 #(
    .INIT(64'h5555FF5DFFFFFFFF)) 
    \bdatw[15]_INST_0_i_69 
       (.I0(\stat_reg[2]_8 ),
        .I1(\bdatw[31]_INST_0_i_72_n_0 ),
        .I2(\bdatw[31]_INST_0_i_71_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_70_n_0 ),
        .I5(\stat_reg[0]_10 ),
        .O(\stat_reg[2]_11 ));
  LUT6 #(
    .INIT(64'h6AAAAAAA6AAAFFFF)) 
    \bdatw[15]_INST_0_i_7 
       (.I0(\stat_reg[0]_5 ),
        .I1(ir[2]),
        .I2(ir[3]),
        .I3(\bdatw[15]_INST_0_i_10_n_0 ),
        .I4(ctl_selb_0),
        .I5(ir[10]),
        .O(\bdatw[15]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0E0EFFFFFF00FFFF)) 
    \bdatw[15]_INST_0_i_70 
       (.I0(\bdatw[15]_INST_0_i_72_n_0 ),
        .I1(\bdatw[31]_INST_0_i_88_n_0 ),
        .I2(\bdatw[15]_INST_0_i_73_n_0 ),
        .I3(\bdatw[15]_INST_0_i_74_n_0 ),
        .I4(ir[12]),
        .I5(ir[11]),
        .O(\bdatw[15]_INST_0_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h4C0FFFFF4CFFFFFF)) 
    \bdatw[15]_INST_0_i_71 
       (.I0(\bdatw[31]_INST_0_i_93_n_0 ),
        .I1(\bdatw[15]_INST_0_i_75_n_0 ),
        .I2(ir[0]),
        .I3(ir[11]),
        .I4(ir[12]),
        .I5(\bdatw[15]_INST_0_i_76_n_0 ),
        .O(\bdatw[15]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h5555555555155555)) 
    \bdatw[15]_INST_0_i_72 
       (.I0(ir[1]),
        .I1(ir[10]),
        .I2(ir[6]),
        .I3(ir[9]),
        .I4(ir[7]),
        .I5(ir[8]),
        .O(\bdatw[15]_INST_0_i_72_n_0 ));
  LUT6 #(
    .INIT(64'h0040555500400040)) 
    \bdatw[15]_INST_0_i_73 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(ir[1]),
        .I2(ir[6]),
        .I3(\bdatw[31]_INST_0_i_95_n_0 ),
        .I4(\bdatw[15]_INST_0_i_77_n_0 ),
        .I5(\ccmd[3]_INST_0_i_23_n_0 ),
        .O(\bdatw[15]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hA200A2A2AAAAAAAA)) 
    \bdatw[15]_INST_0_i_74 
       (.I0(\bdatw[15]_INST_0_i_78_n_0 ),
        .I1(ir[10]),
        .I2(\bdatw[31]_INST_0_i_97_n_0 ),
        .I3(\badr[31]_INST_0_i_149_n_0 ),
        .I4(\bdatw[15]_INST_0_i_79_n_0 ),
        .I5(ir[1]),
        .O(\bdatw[15]_INST_0_i_74_n_0 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \bdatw[15]_INST_0_i_75 
       (.I0(ir[9]),
        .I1(ir[8]),
        .I2(ir[10]),
        .I3(\bdatw[31]_INST_0_i_92_n_0 ),
        .O(\bdatw[15]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'h4040404040FF4040)) 
    \bdatw[15]_INST_0_i_76 
       (.I0(\bdatw[31]_INST_0_i_97_n_0 ),
        .I1(ir[10]),
        .I2(\bdatw[31]_INST_0_i_98_n_0 ),
        .I3(\badr[31]_INST_0_i_149_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(\bdatw[31]_INST_0_i_57_n_0 ),
        .O(\bdatw[15]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'h8FBF7FBF)) 
    \bdatw[15]_INST_0_i_77 
       (.I0(ir[3]),
        .I1(ir[6]),
        .I2(ir[1]),
        .I3(ir[4]),
        .I4(ir[5]),
        .O(\bdatw[15]_INST_0_i_77_n_0 ));
  LUT5 #(
    .INIT(32'hFF7FFFFF)) 
    \bdatw[15]_INST_0_i_78 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(ir[7]),
        .O(\bdatw[15]_INST_0_i_78_n_0 ));
  LUT5 #(
    .INIT(32'h01010111)) 
    \bdatw[15]_INST_0_i_79 
       (.I0(ir[8]),
        .I1(ir[11]),
        .I2(ir[9]),
        .I3(ir[6]),
        .I4(ir[10]),
        .O(\bdatw[15]_INST_0_i_79_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[16]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_14),
        .O(bdatw[16]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[16]_INST_0_i_1 
       (.I0(eir[16]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_16_sn_1),
        .I4(\bbus_o[16]_0 ),
        .O(rst_n_fl_reg_14));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[17]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_13),
        .O(bdatw[17]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[17]_INST_0_i_1 
       (.I0(eir[17]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_17_sn_1),
        .I4(\bbus_o[17]_0 ),
        .O(rst_n_fl_reg_13));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[18]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_12),
        .O(bdatw[18]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[18]_INST_0_i_1 
       (.I0(eir[18]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_18_sn_1),
        .I4(\bbus_o[18]_0 ),
        .O(rst_n_fl_reg_12));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[19]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_11),
        .O(bdatw[19]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[19]_INST_0_i_1 
       (.I0(eir[19]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_19_sn_1),
        .I4(\bbus_o[19]_0 ),
        .O(rst_n_fl_reg_11));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[1]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(bbus_0[0]),
        .O(bdatw[1]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[20]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_10),
        .O(bdatw[20]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[20]_INST_0_i_1 
       (.I0(eir[20]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_20_sn_1),
        .I4(\bbus_o[20]_0 ),
        .O(rst_n_fl_reg_10));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[21]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_9),
        .O(bdatw[21]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[21]_INST_0_i_1 
       (.I0(eir[21]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_21_sn_1),
        .I4(\bbus_o[21]_0 ),
        .O(rst_n_fl_reg_9));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[22]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_8),
        .O(bdatw[22]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[22]_INST_0_i_1 
       (.I0(eir[22]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_22_sn_1),
        .I4(\bbus_o[22]_0 ),
        .O(rst_n_fl_reg_8));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[23]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_7),
        .O(bdatw[23]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[23]_INST_0_i_1 
       (.I0(eir[23]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_23_sn_1),
        .I4(\bbus_o[23]_0 ),
        .O(rst_n_fl_reg_7));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[24]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_6),
        .O(bdatw[24]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[24]_INST_0_i_1 
       (.I0(eir[24]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_24_sn_1),
        .I4(\bbus_o[24]_0 ),
        .O(rst_n_fl_reg_6));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[25]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_16),
        .O(bdatw[25]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[25]_INST_0_i_1 
       (.I0(eir[25]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_25_sn_1),
        .I4(\bbus_o[25]_0 ),
        .O(rst_n_fl_reg_16));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[26]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_5),
        .O(bdatw[26]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[26]_INST_0_i_1 
       (.I0(eir[26]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_26_sn_1),
        .I4(\bbus_o[26]_0 ),
        .O(rst_n_fl_reg_5));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[27]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_4),
        .O(bdatw[27]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[27]_INST_0_i_1 
       (.I0(eir[27]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_27_sn_1),
        .I4(\bbus_o[27]_0 ),
        .O(rst_n_fl_reg_4));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[28]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_3),
        .O(bdatw[28]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[28]_INST_0_i_1 
       (.I0(eir[28]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_28_sn_1),
        .I4(\bbus_o[28]_0 ),
        .O(rst_n_fl_reg_3));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[29]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_2),
        .O(bdatw[29]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[29]_INST_0_i_1 
       (.I0(eir[29]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(bbus_o_29_sn_1),
        .I4(\bbus_o[29]_0 ),
        .O(rst_n_fl_reg_2));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[2]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(bbus_0[1]),
        .O(bdatw[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[30]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_1),
        .O(bdatw[30]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[30]_INST_0_i_1 
       (.I0(eir[30]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\bbus_o[30] ),
        .I4(\bbus_o[30]_0 ),
        .O(rst_n_fl_reg_1));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[31]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(rst_n_fl_reg_0),
        .O(bdatw[31]));
  LUT5 #(
    .INIT(32'h0000000D)) 
    \bdatw[31]_INST_0_i_1 
       (.I0(eir[31]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .I2(\bdatw[31]_INST_0_i_3_n_0 ),
        .I3(\mul_b_reg[31] ),
        .I4(\mul_b_reg[31]_0 ),
        .O(rst_n_fl_reg_0));
  LUT5 #(
    .INIT(32'h00B00000)) 
    \bdatw[31]_INST_0_i_100 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(ir[7]),
        .O(\bdatw[31]_INST_0_i_100_n_0 ));
  LUT4 #(
    .INIT(16'h4044)) 
    \bdatw[31]_INST_0_i_101 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[8]),
        .O(\bdatw[31]_INST_0_i_101_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFF2C)) 
    \bdatw[31]_INST_0_i_102 
       (.I0(ir[6]),
        .I1(ir[8]),
        .I2(ir[7]),
        .I3(ir[9]),
        .I4(ir[10]),
        .O(\bdatw[31]_INST_0_i_102_n_0 ));
  LUT3 #(
    .INIT(8'h9C)) 
    \bdatw[31]_INST_0_i_103 
       (.I0(ir[5]),
        .I1(ir[3]),
        .I2(ir[4]),
        .O(\bdatw[31]_INST_0_i_103_n_0 ));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[31]_INST_0_i_13 
       (.I0(\stat_reg[0]_5 ),
        .I1(ctl_selb_0),
        .I2(\sr_reg[6]_2 ),
        .I3(ctl_selb_rn[1]),
        .I4(ctl_selb_rn[0]),
        .I5(\stat_reg[2]_8 ),
        .O(bbus_sel_cr[4]));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \bdatw[31]_INST_0_i_14 
       (.I0(\stat_reg[0]_5 ),
        .I1(ctl_selb_0),
        .I2(\sr_reg[6]_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_cr[5]));
  LUT6 #(
    .INIT(64'h0000008000000000)) 
    \bdatw[31]_INST_0_i_15 
       (.I0(\stat_reg[0]_5 ),
        .I1(ctl_selb_0),
        .I2(\sr_reg[6]_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_cr[2]));
  LUT6 #(
    .INIT(64'h000CAA000000AA00)) 
    \bdatw[31]_INST_0_i_18 
       (.I0(\bdatw[31]_INST_0_i_46_n_0 ),
        .I1(ir[11]),
        .I2(\ccmd[4]_INST_0_i_2_n_0 ),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\stat[0]_i_24_n_0 ),
        .O(\bdatw[31]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h1040401050000050)) 
    \bdatw[31]_INST_0_i_19 
       (.I0(ir[13]),
        .I1(ir[12]),
        .I2(\iv[15]_i_122_0 ),
        .I3(ir[11]),
        .I4(\sr_reg[13] [5]),
        .I5(\sr_reg[13] [7]),
        .O(\bdatw[31]_INST_0_i_19_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \bdatw[31]_INST_0_i_2 
       (.I0(\stat_reg[0]_5 ),
        .I1(\sr_reg[6]_2 ),
        .I2(ctl_selb_0),
        .O(\bdatw[31]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h01001111FFFFFFFF)) 
    \bdatw[31]_INST_0_i_20 
       (.I0(\bdatw[31]_INST_0_i_47_n_0 ),
        .I1(\bdatw[31]_INST_0_i_48_n_0 ),
        .I2(\bdatw[31]_INST_0_i_49_n_0 ),
        .I3(\bdatw[31]_INST_0_i_50_n_0 ),
        .I4(\iv[15]_i_35_n_0 ),
        .I5(\iv[15]_i_122_0 ),
        .O(\bdatw[31]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \bdatw[31]_INST_0_i_21 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(ir[14]),
        .I2(ir[15]),
        .O(\bdatw[31]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000AE)) 
    \bdatw[31]_INST_0_i_22 
       (.I0(\bdatw[31]_INST_0_i_51_n_0 ),
        .I1(\stat[1]_i_9_n_0 ),
        .I2(\bdatw[31]_INST_0_i_52_n_0 ),
        .I3(ir[14]),
        .I4(ir[15]),
        .I5(\bdatw[31]_INST_0_i_53_n_0 ),
        .O(\bdatw[31]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hDFDD)) 
    \bdatw[31]_INST_0_i_23 
       (.I0(ir[13]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(\bdatw[31]_INST_0_i_46_n_0 ),
        .I3(\stat_reg[2]_12 [0]),
        .O(\bdatw[31]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h10111111FFFFFFFF)) 
    \bdatw[31]_INST_0_i_24 
       (.I0(\bdatw[31]_INST_0_i_54_n_0 ),
        .I1(\bdatw[31]_INST_0_i_55_n_0 ),
        .I2(\bdatw[31]_INST_0_i_56_n_0 ),
        .I3(ir[8]),
        .I4(ir[7]),
        .I5(ir[11]),
        .O(\bdatw[31]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000000011105510)) 
    \bdatw[31]_INST_0_i_25 
       (.I0(ir[8]),
        .I1(ir[7]),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .I3(ir[10]),
        .I4(\stat[1]_i_10_0 ),
        .I5(\bdatw[31]_INST_0_i_57_n_0 ),
        .O(\bdatw[31]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFD0D0DDD0)) 
    \bdatw[31]_INST_0_i_26 
       (.I0(\bdatw[31]_INST_0_i_58_n_0 ),
        .I1(\bdatw[31]_INST_0_i_59_n_0 ),
        .I2(\ccmd[4]_INST_0_i_1_n_0 ),
        .I3(ir[10]),
        .I4(ir[11]),
        .I5(\bdatw[31]_INST_0_i_60_n_0 ),
        .O(\bdatw[31]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000000A8)) 
    \bdatw[31]_INST_0_i_27 
       (.I0(\iv[15]_i_14_n_0 ),
        .I1(\bdatw[31]_INST_0_i_7_0 ),
        .I2(\bdatw[31]_INST_0_i_7_1 ),
        .I3(\bdatw[31]_INST_0_i_63_n_0 ),
        .I4(\bdatw[31]_INST_0_i_64_n_0 ),
        .I5(\bdatw[31]_INST_0_i_65_n_0 ),
        .O(\bdatw[31]_INST_0_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEFFEFFFFFFFEF)) 
    \bdatw[31]_INST_0_i_28 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(ir[15]),
        .I2(\bdatw[31]_INST_0_i_27_n_0 ),
        .I3(ir[2]),
        .I4(ir[14]),
        .I5(ir[12]),
        .O(\bdatw[31]_INST_0_i_28_n_0 ));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_29 
       (.I0(ctl_selb_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\sr_reg[6]_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_0[3]));
  LUT3 #(
    .INIT(8'hA8)) 
    \bdatw[31]_INST_0_i_3 
       (.I0(\bdatw[31]_INST_0_i_8_n_0 ),
        .I1(ctl_selb_0),
        .I2(ir[10]),
        .O(\bdatw[31]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bdatw[31]_INST_0_i_30 
       (.I0(ctl_selb_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\sr_reg[6]_2 ),
        .I3(ctl_selb_rn[0]),
        .I4(\stat_reg[2]_8 ),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_0[4]));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bdatw[31]_INST_0_i_31 
       (.I0(ctl_selb_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\sr_reg[6]_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_0[1]));
  LUT6 #(
    .INIT(64'h0000000000200000)) 
    \bdatw[31]_INST_0_i_32 
       (.I0(ctl_selb_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\sr_reg[6]_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(ctl_selb_rn[1]),
        .I5(ctl_selb_rn[0]),
        .O(bbus_sel_0[2]));
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \bdatw[31]_INST_0_i_33 
       (.I0(\stat_reg[2]_8 ),
        .I1(ctl_selb_0),
        .I2(\stat_reg[0]_5 ),
        .I3(\sr_reg[6]_2 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_0[7]));
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    \bdatw[31]_INST_0_i_34 
       (.I0(ctl_selb_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\sr_reg[6]_2 ),
        .I3(\stat_reg[2]_8 ),
        .I4(ctl_selb_rn[0]),
        .I5(ctl_selb_rn[1]),
        .O(bbus_sel_0[0]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_35 
       (.I0(ctl_selb_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\sr_reg[6]_2 ),
        .I3(ctl_selb_rn[1]),
        .I4(ctl_selb_rn[0]),
        .I5(\stat_reg[2]_8 ),
        .O(bbus_sel_0[5]));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \bdatw[31]_INST_0_i_36 
       (.I0(ctl_selb_0),
        .I1(\stat_reg[0]_5 ),
        .I2(\sr_reg[6]_2 ),
        .I3(ctl_selb_rn[0]),
        .I4(ctl_selb_rn[1]),
        .I5(\stat_reg[2]_8 ),
        .O(bbus_sel_0[6]));
  LUT6 #(
    .INIT(64'h1011101010111011)) 
    \bdatw[31]_INST_0_i_37 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(\bdatw[31]_INST_0_i_66_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_68_n_0 ),
        .I5(\bdatw[31]_INST_0_i_69_n_0 ),
        .O(ctl_selb_rn[1]));
  LUT6 #(
    .INIT(64'h1011101010111011)) 
    \bdatw[31]_INST_0_i_38 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(\bdatw[31]_INST_0_i_70_n_0 ),
        .I3(\bdatw[31]_INST_0_i_67_n_0 ),
        .I4(\bdatw[31]_INST_0_i_71_n_0 ),
        .I5(\bdatw[31]_INST_0_i_72_n_0 ),
        .O(ctl_selb_rn[0]));
  LUT6 #(
    .INIT(64'h4544454445454544)) 
    \bdatw[31]_INST_0_i_39 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\badr[31]_INST_0_i_59_n_0 ),
        .I2(\bdatw[31]_INST_0_i_73_n_0 ),
        .I3(\bdatw[31]_INST_0_i_74_n_0 ),
        .I4(\bdatw[31]_INST_0_i_75_n_0 ),
        .I5(\bdatw[31]_INST_0_i_76_n_0 ),
        .O(\stat_reg[2]_8 ));
  LUT6 #(
    .INIT(64'h0020000020000000)) 
    \bdatw[31]_INST_0_i_46 
       (.I0(ir[6]),
        .I1(ir[8]),
        .I2(ir[7]),
        .I3(ir[9]),
        .I4(ir[10]),
        .I5(ir[11]),
        .O(\bdatw[31]_INST_0_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h4444444544454445)) 
    \bdatw[31]_INST_0_i_47 
       (.I0(ir[11]),
        .I1(\bdatw[31]_INST_0_i_77_n_0 ),
        .I2(\bdatw[31]_INST_0_i_78_n_0 ),
        .I3(\stat[1]_i_10_0 ),
        .I4(\bdatw[31]_INST_0_i_79_n_0 ),
        .I5(rst_n_fl_reg_17),
        .O(\bdatw[31]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF1400)) 
    \bdatw[31]_INST_0_i_48 
       (.I0(rst_n_fl_reg_17),
        .I1(ir[6]),
        .I2(ir[9]),
        .I3(\bdatw[31]_INST_0_i_80_n_0 ),
        .I4(\bdatw[31]_INST_0_i_81_n_0 ),
        .O(\bdatw[31]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h383338FF30CC30CC)) 
    \bdatw[31]_INST_0_i_49 
       (.I0(ir[5]),
        .I1(ir[10]),
        .I2(ir[6]),
        .I3(ir[9]),
        .I4(\stat[1]_i_10_0 ),
        .I5(ir[7]),
        .O(\bdatw[31]_INST_0_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hF7FFFF77FFFFF7FF)) 
    \bdatw[31]_INST_0_i_50 
       (.I0(ir[6]),
        .I1(ir[9]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[3]),
        .I5(ir[7]),
        .O(\bdatw[31]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hEEFFFBAAAAAAAAAA)) 
    \bdatw[31]_INST_0_i_51 
       (.I0(ir[12]),
        .I1(\sr_reg[13] [6]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[13]),
        .I4(ir[11]),
        .I5(\iv_reg[0] ),
        .O(\bdatw[31]_INST_0_i_51_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFDDDB)) 
    \bdatw[31]_INST_0_i_52 
       (.I0(ir[0]),
        .I1(ir[3]),
        .I2(\stat_reg[2]_12 [2]),
        .I3(\stat_reg[2]_12 [1]),
        .I4(\bdatw[31]_INST_0_i_82_n_0 ),
        .O(\bdatw[31]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h22288828AAAAAAAA)) 
    \bdatw[31]_INST_0_i_53 
       (.I0(ir[12]),
        .I1(ir[11]),
        .I2(\sr_reg[13] [4]),
        .I3(ir[13]),
        .I4(\sr_reg[13] [7]),
        .I5(\iv_reg[0] ),
        .O(\bdatw[31]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000860000)) 
    \bdatw[31]_INST_0_i_54 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[3]),
        .I3(ir[7]),
        .I4(ir[6]),
        .I5(\ccmd[4]_INST_0_i_2_n_0 ),
        .O(\bdatw[31]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h03F00FF3073F0F33)) 
    \bdatw[31]_INST_0_i_55 
       (.I0(\stat[1]_i_10_0 ),
        .I1(ir[8]),
        .I2(ir[9]),
        .I3(ir[10]),
        .I4(ir[7]),
        .I5(ir[6]),
        .O(\bdatw[31]_INST_0_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hE6EE66666E66666E)) 
    \bdatw[31]_INST_0_i_56 
       (.I0(ir[9]),
        .I1(ir[10]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[6]),
        .I5(ir[3]),
        .O(\bdatw[31]_INST_0_i_56_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[31]_INST_0_i_57 
       (.I0(ir[10]),
        .I1(ir[6]),
        .I2(ir[9]),
        .O(\bdatw[31]_INST_0_i_57_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEAFAFAFAE)) 
    \bdatw[31]_INST_0_i_58 
       (.I0(\bcmd[1]_INST_0_i_5_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(ir[9]),
        .I3(ir[10]),
        .I4(ir[11]),
        .I5(ir[6]),
        .O(\bdatw[31]_INST_0_i_58_n_0 ));
  LUT6 #(
    .INIT(64'hF080808080808080)) 
    \bdatw[31]_INST_0_i_59 
       (.I0(ir[9]),
        .I1(ir[10]),
        .I2(ir[6]),
        .I3(ir[7]),
        .I4(ir[8]),
        .I5(rst_n_fl_reg_17),
        .O(\bdatw[31]_INST_0_i_59_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF33FF10)) 
    \bdatw[31]_INST_0_i_6 
       (.I0(\bdatw[31]_INST_0_i_18_n_0 ),
        .I1(\bdatw[31]_INST_0_i_19_n_0 ),
        .I2(\bdatw[31]_INST_0_i_20_n_0 ),
        .I3(\bdatw[31]_INST_0_i_21_n_0 ),
        .I4(ctl_fetch_inferred_i_17_n_0),
        .I5(\bdatw[31]_INST_0_i_22_n_0 ),
        .O(\stat_reg[0]_5 ));
  LUT6 #(
    .INIT(64'hAAAAAAAABAAAAAAA)) 
    \bdatw[31]_INST_0_i_60 
       (.I0(\bdatw[31]_INST_0_i_46_n_0 ),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[7]),
        .I4(ir[10]),
        .I5(\stat[1]_i_10_0 ),
        .O(\bdatw[31]_INST_0_i_60_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[31]_INST_0_i_63 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(ir[13]),
        .O(\bdatw[31]_INST_0_i_63_n_0 ));
  LUT3 #(
    .INIT(8'hE7)) 
    \bdatw[31]_INST_0_i_64 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[3]),
        .I2(ir[0]),
        .O(\bdatw[31]_INST_0_i_64_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \bdatw[31]_INST_0_i_65 
       (.I0(ir[1]),
        .I1(ir[7]),
        .I2(ir[5]),
        .I3(ir[4]),
        .O(\bdatw[31]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \bdatw[31]_INST_0_i_66 
       (.I0(\tr[31]_i_49_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(ir[8]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(ir[1]),
        .I5(\bdatw[31]_INST_0_i_83_n_0 ),
        .O(\bdatw[31]_INST_0_i_66_n_0 ));
  LUT4 #(
    .INIT(16'hFFF7)) 
    \bdatw[31]_INST_0_i_67 
       (.I0(ir[14]),
        .I1(ir[13]),
        .I2(ir[15]),
        .I3(\stat_reg[2]_12 [0]),
        .O(\bdatw[31]_INST_0_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h808880888088AAAA)) 
    \bdatw[31]_INST_0_i_68 
       (.I0(\badr[31]_INST_0_i_85_n_0 ),
        .I1(ir[1]),
        .I2(\bdatw[31]_INST_0_i_84_n_0 ),
        .I3(\bdatw[31]_INST_0_i_85_n_0 ),
        .I4(\bcmd[3]_INST_0_i_16_n_0 ),
        .I5(\bdatw[31]_INST_0_i_86_n_0 ),
        .O(\bdatw[31]_INST_0_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0EEFFFFFFFF)) 
    \bdatw[31]_INST_0_i_69 
       (.I0(\bcmd[3]_INST_0_i_16_n_0 ),
        .I1(\bdatw[31]_INST_0_i_87_n_0 ),
        .I2(\bdatw[31]_INST_0_i_88_n_0 ),
        .I3(\bdatw[31]_INST_0_i_89_n_0 ),
        .I4(ir[1]),
        .I5(\bdatw[31]_INST_0_i_90_n_0 ),
        .O(\bdatw[31]_INST_0_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF5551)) 
    \bdatw[31]_INST_0_i_7 
       (.I0(\bdatw[31]_INST_0_i_23_n_0 ),
        .I1(\bdatw[31]_INST_0_i_24_n_0 ),
        .I2(\bdatw[31]_INST_0_i_25_n_0 ),
        .I3(\bdatw[31]_INST_0_i_26_n_0 ),
        .I4(\bdatw[31]_INST_0_i_27_n_0 ),
        .I5(\bdatw[31]_INST_0_i_28_n_0 ),
        .O(ctl_selb_0));
  LUT6 #(
    .INIT(64'h40400000404000FF)) 
    \bdatw[31]_INST_0_i_70 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(ir[0]),
        .I2(\bdatw[31]_INST_0_i_46_n_0 ),
        .I3(\badr[31]_INST_0_i_32_n_0 ),
        .I4(\stat_reg[2]_12 [0]),
        .I5(ir[15]),
        .O(\bdatw[31]_INST_0_i_70_n_0 ));
  LUT5 #(
    .INIT(32'h00E00000)) 
    \bdatw[31]_INST_0_i_71 
       (.I0(\bdatw[31]_INST_0_i_84_n_0 ),
        .I1(\bdatw[31]_INST_0_i_91_n_0 ),
        .I2(ir[12]),
        .I3(ir[11]),
        .I4(ir[0]),
        .O(\bdatw[31]_INST_0_i_71_n_0 ));
  LUT6 #(
    .INIT(64'h5555DFFFDFFFDFFF)) 
    \bdatw[31]_INST_0_i_72 
       (.I0(\bdatw[31]_INST_0_i_90_n_0 ),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(ir[10]),
        .I3(\bdatw[31]_INST_0_i_92_n_0 ),
        .I4(\bdatw[31]_INST_0_i_93_n_0 ),
        .I5(ir[0]),
        .O(\bdatw[31]_INST_0_i_72_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFDFCC)) 
    \bdatw[31]_INST_0_i_73 
       (.I0(\bdatw[31]_INST_0_i_46_n_0 ),
        .I1(\stat_reg[2]_12 [1]),
        .I2(ir[2]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\bdatw[31]_INST_0_i_73_n_0 ));
  LUT6 #(
    .INIT(64'hAEFFAEAEAAAAAAAA)) 
    \bdatw[31]_INST_0_i_74 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\bdatw[31]_INST_0_i_94_n_0 ),
        .I2(\bdatw[31]_INST_0_i_95_n_0 ),
        .I3(\bdatw[31]_INST_0_i_96_n_0 ),
        .I4(\ccmd[3]_INST_0_i_23_n_0 ),
        .I5(\iv[15]_i_30_n_0 ),
        .O(\bdatw[31]_INST_0_i_74_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF4040FF40)) 
    \bdatw[31]_INST_0_i_75 
       (.I0(\bdatw[31]_INST_0_i_97_n_0 ),
        .I1(ir[10]),
        .I2(\bdatw[31]_INST_0_i_98_n_0 ),
        .I3(\badr[31]_INST_0_i_54_n_0 ),
        .I4(\bdatw[31]_INST_0_i_99_n_0 ),
        .I5(ir[11]),
        .O(\bdatw[31]_INST_0_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hBAAA0000FFFFFFFF)) 
    \bdatw[31]_INST_0_i_76 
       (.I0(\bdatw[31]_INST_0_i_100_n_0 ),
        .I1(\bdatw[31]_INST_0_i_101_n_0 ),
        .I2(\stat[0]_i_34_n_0 ),
        .I3(\bdatw[31]_INST_0_i_102_n_0 ),
        .I4(ir[11]),
        .I5(ir[2]),
        .O(\bdatw[31]_INST_0_i_76_n_0 ));
  LUT5 #(
    .INIT(32'hA8006000)) 
    \bdatw[31]_INST_0_i_77 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[9]),
        .I3(ir[10]),
        .I4(ir[8]),
        .O(\bdatw[31]_INST_0_i_77_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[31]_INST_0_i_78 
       (.I0(ir[9]),
        .I1(ir[8]),
        .O(\bdatw[31]_INST_0_i_78_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[31]_INST_0_i_79 
       (.I0(ir[10]),
        .I1(ir[7]),
        .O(\bdatw[31]_INST_0_i_79_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[31]_INST_0_i_8 
       (.I0(\sr_reg[6]_2 ),
        .I1(\stat_reg[0]_5 ),
        .O(\bdatw[31]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0830000000000000)) 
    \bdatw[31]_INST_0_i_80 
       (.I0(ir[7]),
        .I1(ir[8]),
        .I2(ir[9]),
        .I3(ir[10]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\bdatw[31]_INST_0_i_80_n_0 ));
  LUT6 #(
    .INIT(64'h1100110005045504)) 
    \bdatw[31]_INST_0_i_81 
       (.I0(ir[8]),
        .I1(ir[10]),
        .I2(ir[7]),
        .I3(ir[11]),
        .I4(ir[6]),
        .I5(ir[9]),
        .O(\bdatw[31]_INST_0_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFEFFFEFF)) 
    \bdatw[31]_INST_0_i_82 
       (.I0(ir[2]),
        .I1(ir[1]),
        .I2(ir[13]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\stat_reg[2]_12 [1]),
        .O(\bdatw[31]_INST_0_i_82_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \bdatw[31]_INST_0_i_83 
       (.I0(ir[7]),
        .I1(ir[6]),
        .O(\bdatw[31]_INST_0_i_83_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001F00)) 
    \bdatw[31]_INST_0_i_84 
       (.I0(ir[10]),
        .I1(ir[6]),
        .I2(ir[9]),
        .I3(\ccmd[3]_INST_0_i_10_n_0 ),
        .I4(\stat[1]_i_10_0 ),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\bdatw[31]_INST_0_i_84_n_0 ));
  LUT6 #(
    .INIT(64'h1022BAEEFFFFFFFF)) 
    \bdatw[31]_INST_0_i_85 
       (.I0(ir[8]),
        .I1(ir[9]),
        .I2(\stat[1]_i_10_0 ),
        .I3(ir[7]),
        .I4(ir[6]),
        .I5(ir[10]),
        .O(\bdatw[31]_INST_0_i_85_n_0 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \bdatw[31]_INST_0_i_86 
       (.I0(ir[7]),
        .I1(ir[8]),
        .I2(ir[6]),
        .O(\bdatw[31]_INST_0_i_86_n_0 ));
  LUT6 #(
    .INIT(64'hDD00F5F5FFFFFFFF)) 
    \bdatw[31]_INST_0_i_87 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(\bdatw[31]_INST_0_i_103_n_0 ),
        .I2(\stat[0]_i_32_n_0 ),
        .I3(\bdatw[31]_INST_0_i_95_n_0 ),
        .I4(ir[6]),
        .I5(ir[1]),
        .O(\bdatw[31]_INST_0_i_87_n_0 ));
  LUT6 #(
    .INIT(64'hA8999988ECDD8888)) 
    \bdatw[31]_INST_0_i_88 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(\stat[1]_i_10_0 ),
        .I3(ir[7]),
        .I4(ir[8]),
        .I5(ir[6]),
        .O(\bdatw[31]_INST_0_i_88_n_0 ));
  LUT5 #(
    .INIT(32'h04000000)) 
    \bdatw[31]_INST_0_i_89 
       (.I0(ir[8]),
        .I1(ir[7]),
        .I2(ir[9]),
        .I3(ir[6]),
        .I4(ir[10]),
        .O(\bdatw[31]_INST_0_i_89_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_90 
       (.I0(ir[12]),
        .I1(ir[11]),
        .O(\bdatw[31]_INST_0_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h8888808028280AAA)) 
    \bdatw[31]_INST_0_i_91 
       (.I0(ir[10]),
        .I1(ir[6]),
        .I2(ir[7]),
        .I3(\stat[1]_i_10_0 ),
        .I4(ir[9]),
        .I5(ir[8]),
        .O(\bdatw[31]_INST_0_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h2822C220A00C0000)) 
    \bdatw[31]_INST_0_i_92 
       (.I0(ir[0]),
        .I1(ir[3]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[7]),
        .I5(ir[6]),
        .O(\bdatw[31]_INST_0_i_92_n_0 ));
  LUT6 #(
    .INIT(64'h00001FDFBBBBD3D3)) 
    \bdatw[31]_INST_0_i_93 
       (.I0(ir[6]),
        .I1(ir[8]),
        .I2(ir[7]),
        .I3(\stat[1]_i_10_0 ),
        .I4(ir[9]),
        .I5(ir[10]),
        .O(\bdatw[31]_INST_0_i_93_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[31]_INST_0_i_94 
       (.I0(ir[6]),
        .I1(ir[2]),
        .O(\bdatw[31]_INST_0_i_94_n_0 ));
  LUT5 #(
    .INIT(32'hFFEBFFFF)) 
    \bdatw[31]_INST_0_i_95 
       (.I0(ir[3]),
        .I1(ir[4]),
        .I2(ir[5]),
        .I3(ir[7]),
        .I4(ir[8]),
        .O(\bdatw[31]_INST_0_i_95_n_0 ));
  LUT5 #(
    .INIT(32'h9C5FFFFF)) 
    \bdatw[31]_INST_0_i_96 
       (.I0(ir[5]),
        .I1(ir[3]),
        .I2(ir[4]),
        .I3(ir[6]),
        .I4(ir[2]),
        .O(\bdatw[31]_INST_0_i_96_n_0 ));
  LUT6 #(
    .INIT(64'h5555777711110CCC)) 
    \bdatw[31]_INST_0_i_97 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(div_crdy),
        .I3(crdy),
        .I4(ir[9]),
        .I5(ir[8]),
        .O(\bdatw[31]_INST_0_i_97_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7777F777)) 
    \bdatw[31]_INST_0_i_98 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(div_crdy),
        .I3(crdy),
        .I4(ir[9]),
        .I5(ir[8]),
        .O(\bdatw[31]_INST_0_i_98_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFA8FFFFFF)) 
    \bdatw[31]_INST_0_i_99 
       (.I0(ir[9]),
        .I1(ir[6]),
        .I2(ir[10]),
        .I3(crdy),
        .I4(div_crdy),
        .I5(ir[8]),
        .O(\bdatw[31]_INST_0_i_99_n_0 ));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[3]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(bbus_0[2]),
        .O(bdatw[3]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[4]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(bbus_0[3]),
        .O(bdatw[4]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[5]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(\bdatw[5] [1]),
        .O(bdatw[5]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[6]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(bbus_0[4]),
        .O(bdatw[6]));
  LUT3 #(
    .INIT(8'hE0)) 
    \bdatw[7]_INST_0 
       (.I0(\stat_reg[0]_4 ),
        .I1(\stat_reg[2]_6 ),
        .I2(bbus_0[5]),
        .O(bdatw[7]));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[8]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(\bdatw[5] [0]),
        .I4(bbus_0[6]),
        .O(bdatw[8]));
  LUT5 #(
    .INIT(32'hFFFFFFAE)) 
    \bdatw[8]_INST_0_i_2 
       (.I0(\bdatw[8]_INST_0_i_9_n_0 ),
        .I1(eir[8]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\mul_b_reg[8] ),
        .I4(\mul_b_reg[8]_0 ),
        .O(bbus_0[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \bdatw[8]_INST_0_i_21 
       (.I0(bbus_sel_cr[0]),
        .I1(\sr_reg[13] [0]),
        .O(bbus_sr[0]));
  LUT6 #(
    .INIT(64'h000000000F2DF000)) 
    \bdatw[8]_INST_0_i_3 
       (.I0(\bdatw[9]_INST_0_i_10_n_0 ),
        .I1(ir[1]),
        .I2(\stat_reg[0]_5 ),
        .I3(ir[0]),
        .I4(ctl_selb_0),
        .I5(\sr_reg[6]_2 ),
        .O(rst_n_fl_reg_18));
  LUT2 #(
    .INIT(4'h2)) 
    \bdatw[8]_INST_0_i_4 
       (.I0(eir[0]),
        .I1(\bdatw[31]_INST_0_i_2_n_0 ),
        .O(rst_n_fl_reg_21));
  LUT6 #(
    .INIT(64'h3000000002323232)) 
    \bdatw[8]_INST_0_i_9 
       (.I0(ir[7]),
        .I1(\sr_reg[6]_2 ),
        .I2(ctl_selb_0),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\bdatw[11]_INST_0_i_19_n_0 ),
        .I5(\stat_reg[0]_5 ),
        .O(\bdatw[8]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hDC548800)) 
    \bdatw[9]_INST_0 
       (.I0(\stat_reg[1] ),
        .I1(\stat_reg[2]_6 ),
        .I2(\stat_reg[0]_4 ),
        .I3(bbus_0[0]),
        .I4(bbus_0[7]),
        .O(bdatw[9]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFAE)) 
    \bdatw[9]_INST_0_i_1 
       (.I0(\bdatw[9]_INST_0_i_3_n_0 ),
        .I1(eir[1]),
        .I2(\bdatw[31]_INST_0_i_2_n_0 ),
        .I3(\mul_b_reg[1] ),
        .I4(\mul_b_reg[1]_0 ),
        .I5(\mul_b_reg[1]_1 ),
        .O(bbus_0[0]));
  LUT2 #(
    .INIT(4'h1)) 
    \bdatw[9]_INST_0_i_10 
       (.I0(ir[3]),
        .I1(ir[2]),
        .O(\bdatw[9]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF11F1)) 
    \bdatw[9]_INST_0_i_2 
       (.I0(\bdatw[9]_INST_0_i_7_n_0 ),
        .I1(\sr_reg[6]_2 ),
        .I2(eir[9]),
        .I3(\bdatw[31]_INST_0_i_2_n_0 ),
        .I4(\mul_b_reg[9] ),
        .I5(\mul_b_reg[9]_0 ),
        .O(bbus_0[7]));
  LUT2 #(
    .INIT(4'hE)) 
    \bdatw[9]_INST_0_i_20 
       (.I0(ir[2]),
        .I1(ir[1]),
        .O(\bdatw[9]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0540050054145454)) 
    \bdatw[9]_INST_0_i_3 
       (.I0(\sr_reg[6]_2 ),
        .I1(ir[0]),
        .I2(ctl_selb_0),
        .I3(ir[1]),
        .I4(\bdatw[9]_INST_0_i_10_n_0 ),
        .I5(\stat_reg[0]_5 ),
        .O(\bdatw[9]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAA6AAAAAAA6AFFFF)) 
    \bdatw[9]_INST_0_i_7 
       (.I0(\stat_reg[0]_5 ),
        .I1(ir[0]),
        .I2(ir[3]),
        .I3(\bdatw[9]_INST_0_i_20_n_0 ),
        .I4(ctl_selb_0),
        .I5(ir[8]),
        .O(\bdatw[9]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[0]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(ccmd[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF55555504)) 
    \ccmd[0]_INST_0_i_1 
       (.I0(\ccmd[0]_INST_0_i_2_n_0 ),
        .I1(\sr_reg[13] [6]),
        .I2(ir[12]),
        .I3(ir[15]),
        .I4(\ccmd[0]_INST_0_i_3_n_0 ),
        .I5(\ccmd[0]_INST_0_i_4_n_0 ),
        .O(\ccmd[0]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'hAAA2AAAAAAAAAAAA)) 
    \ccmd[0]_INST_0_i_10 
       (.I0(\ccmd[3]_INST_0_i_16_n_0 ),
        .I1(ir[6]),
        .I2(ir[9]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\ccmd[3]_INST_0_i_13_n_0 ),
        .I5(\niho_dsp_a[32]_INST_0_i_9_0 ),
        .O(\ccmd[0]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEEEAFFFFFEFA)) 
    \ccmd[0]_INST_0_i_11 
       (.I0(\ccmd[0]_INST_0_i_17_n_0 ),
        .I1(ir[8]),
        .I2(\stat[1]_i_10_0 ),
        .I3(ir[9]),
        .I4(ir[11]),
        .I5(rst_n_fl_reg_17),
        .O(\ccmd[0]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hBABBBBBBBBBABBBA)) 
    \ccmd[0]_INST_0_i_12 
       (.I0(\ccmd[0]_INST_0_i_18_n_0 ),
        .I1(\ccmd[0]_INST_0_i_19_n_0 ),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(ir[10]),
        .I5(ir[7]),
        .O(\ccmd[0]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hDFDFDFDFDFDDDFDF)) 
    \ccmd[0]_INST_0_i_13 
       (.I0(\ccmd[3]_INST_0_i_9_n_0 ),
        .I1(ir[2]),
        .I2(\ccmd[0]_INST_0_i_20_n_0 ),
        .I3(\ccmd[3]_INST_0_i_12_n_0 ),
        .I4(\ccmd[0]_INST_0_i_21_n_0 ),
        .I5(\bcmd[3]_INST_0_i_4_n_0 ),
        .O(\ccmd[0]_INST_0_i_13_n_0 ));
  LUT4 #(
    .INIT(16'h8000)) 
    \ccmd[0]_INST_0_i_15 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(ir[8]),
        .I3(ir[9]),
        .O(\ccmd[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h3FFF3FFB2EEA2EEA)) 
    \ccmd[0]_INST_0_i_17 
       (.I0(ir[6]),
        .I1(ir[10]),
        .I2(ir[9]),
        .I3(ir[7]),
        .I4(ir[8]),
        .I5(rst_n_fl_reg_17),
        .O(\ccmd[0]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h002008A002000020)) 
    \ccmd[0]_INST_0_i_18 
       (.I0(\ccmd[0]_INST_0_i_15_n_0 ),
        .I1(ir[4]),
        .I2(ir[7]),
        .I3(ir[6]),
        .I4(ir[3]),
        .I5(ir[5]),
        .O(\ccmd[0]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hDFDDDDDDDFDDDFDD)) 
    \ccmd[0]_INST_0_i_19 
       (.I0(ir[11]),
        .I1(ir[9]),
        .I2(\ccmd[0]_INST_0_i_22_n_0 ),
        .I3(ir[6]),
        .I4(\stat[1]_i_10_0 ),
        .I5(ir[7]),
        .O(\ccmd[0]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h0505FFFF0040FFFF)) 
    \ccmd[0]_INST_0_i_2 
       (.I0(ir[12]),
        .I1(\sr_reg[13] [6]),
        .I2(ir[11]),
        .I3(ir[14]),
        .I4(ir[13]),
        .I5(ir[15]),
        .O(\ccmd[0]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h4000000000000000)) 
    \ccmd[0]_INST_0_i_20 
       (.I0(ir[6]),
        .I1(ir[3]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\iv[15]_i_122_0 ),
        .I5(\ccmd[3]_INST_0_i_18_n_0 ),
        .O(\ccmd[0]_INST_0_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \ccmd[0]_INST_0_i_21 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[0]),
        .I2(ir[3]),
        .O(\ccmd[0]_INST_0_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[0]_INST_0_i_22 
       (.I0(ir[10]),
        .I1(ir[8]),
        .O(\ccmd[0]_INST_0_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hAAFF3CCCAAFFFFFF)) 
    \ccmd[0]_INST_0_i_3 
       (.I0(\ccmd[0]_INST_0_i_5_n_0 ),
        .I1(ir[11]),
        .I2(\sr_reg[13] [7]),
        .I3(ir[12]),
        .I4(ir[14]),
        .I5(\iv[15]_i_122_0 ),
        .O(\ccmd[0]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAEFFFAAAAAAAA)) 
    \ccmd[0]_INST_0_i_4 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(ir[15]),
        .I2(ir[12]),
        .I3(\stat_reg[1]_0 ),
        .I4(\ccmd[0]_INST_0_i_7_n_0 ),
        .I5(\ccmd[0]_INST_0_i_8_n_0 ),
        .O(\ccmd[0]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hCCCCCCCC888800C0)) 
    \ccmd[0]_INST_0_i_5 
       (.I0(\ccmd[0]_INST_0_i_9_n_0 ),
        .I1(\ccmd[0]_INST_0_i_10_n_0 ),
        .I2(\ccmd[0]_INST_0_i_11_n_0 ),
        .I3(\ccmd[0]_INST_0_i_12_n_0 ),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\stat_reg[2]_12 [1]),
        .O(\ccmd[0]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h5E000000FFFFFFFF)) 
    \ccmd[0]_INST_0_i_7 
       (.I0(ir[14]),
        .I1(ir[12]),
        .I2(ir[11]),
        .I3(\iv[15]_i_122_0 ),
        .I4(ir[15]),
        .I5(\ccmd[0]_INST_0_i_2_n_0 ),
        .O(\ccmd[0]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h00FFB0B0FFFFFFFF)) 
    \ccmd[0]_INST_0_i_8 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\ccmd[3]_INST_0_i_19_n_0 ),
        .I2(\ccmd[0]_INST_0_i_13_n_0 ),
        .I3(\ccmd[0]_INST_0_i_4_0 ),
        .I4(ir[14]),
        .I5(\stat[1]_i_5_n_0 ),
        .O(\ccmd[0]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFF7FEFFFFFFFFFFF)) 
    \ccmd[0]_INST_0_i_9 
       (.I0(ir[4]),
        .I1(ir[5]),
        .I2(ir[3]),
        .I3(ir[7]),
        .I4(ir[6]),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\ccmd[0]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(ccmd[1]));
  LUT6 #(
    .INIT(64'h000000000000EE0E)) 
    \ccmd[1]_INST_0_i_1 
       (.I0(\ccmd[1]_INST_0_i_2_n_0 ),
        .I1(\bcmd[2] ),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(\ccmd[1]_INST_0_i_3_n_0 ),
        .I4(\ccmd[1]_INST_0_i_4_n_0 ),
        .I5(\ccmd[1]_INST_0_i_5_n_0 ),
        .O(\ccmd[1]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[1]_INST_0_i_11 
       (.I0(ir[11]),
        .I1(ir[10]),
        .O(\ccmd[1]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \ccmd[1]_INST_0_i_13 
       (.I0(ir[14]),
        .I1(ir[13]),
        .I2(ir[12]),
        .I3(ir[7]),
        .I4(ir[8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\ccmd[1]_INST_0_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hE7)) 
    \ccmd[1]_INST_0_i_14 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(ir[0]),
        .I2(ir[3]),
        .O(\ccmd[1]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h77779F1F7F7FFF7F)) 
    \ccmd[1]_INST_0_i_15 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(ir[7]),
        .I3(\stat[1]_i_10_0 ),
        .I4(ir[9]),
        .I5(ir[6]),
        .O(\ccmd[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00010100)) 
    \ccmd[1]_INST_0_i_16 
       (.I0(rst_n_fl_reg_17),
        .I1(ir[8]),
        .I2(ir[10]),
        .I3(ir[6]),
        .I4(ir[7]),
        .I5(\ccmd[1]_INST_0_i_18_n_0 ),
        .O(\ccmd[1]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[1]_INST_0_i_17 
       (.I0(ir[9]),
        .I1(ir[10]),
        .O(\ccmd[1]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000F10)) 
    \ccmd[1]_INST_0_i_18 
       (.I0(\iv[15]_i_87_n_0 ),
        .I1(ir[9]),
        .I2(ir[10]),
        .I3(ir[11]),
        .I4(ir[8]),
        .I5(ir[6]),
        .O(\ccmd[1]_INST_0_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hEEE0E0EEEEEEEEEE)) 
    \ccmd[1]_INST_0_i_2 
       (.I0(\ccmd[1]_INST_0_i_6_n_0 ),
        .I1(\ccmd[1]_INST_0_i_7_n_0 ),
        .I2(ir[9]),
        .I3(\ccmd[1]_INST_0_i_8_n_0 ),
        .I4(ir[10]),
        .I5(\ccmd[1]_INST_0_i_9_n_0 ),
        .O(\ccmd[1]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFDFFFFFFFFFF)) 
    \ccmd[1]_INST_0_i_3 
       (.I0(\bcmd[0]_INST_0_i_12_n_0 ),
        .I1(ir[7]),
        .I2(ir[3]),
        .I3(\iv_reg[0]_0 ),
        .I4(\ccmd[1]_INST_0_i_11_n_0 ),
        .I5(\bcmd[1]_INST_0_i_13_n_0 ),
        .O(\ccmd[1]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h0880888008880888)) 
    \ccmd[1]_INST_0_i_4 
       (.I0(ir[15]),
        .I1(\iv_reg[0] ),
        .I2(ir[14]),
        .I3(ir[13]),
        .I4(ir[12]),
        .I5(ir[11]),
        .O(\ccmd[1]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \ccmd[1]_INST_0_i_5 
       (.I0(ir[2]),
        .I1(ir[11]),
        .I2(\ccmd[1]_INST_0_i_1_0 ),
        .I3(\ccmd[1]_INST_0_i_13_n_0 ),
        .I4(\ccmd[1]_INST_0_i_14_n_0 ),
        .I5(\ccmd[3]_INST_0_i_12_n_0 ),
        .O(\ccmd[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DCDB555F)) 
    \ccmd[1]_INST_0_i_6 
       (.I0(ir[4]),
        .I1(ir[3]),
        .I2(ir[5]),
        .I3(ir[7]),
        .I4(ir[6]),
        .I5(\bcmd[3]_INST_0_i_16_n_0 ),
        .O(\ccmd[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF80FF)) 
    \ccmd[1]_INST_0_i_7 
       (.I0(ir[7]),
        .I1(ir[9]),
        .I2(ir[5]),
        .I3(ir[8]),
        .I4(\ccmd[1]_INST_0_i_15_n_0 ),
        .I5(\ccmd[1]_INST_0_i_16_n_0 ),
        .O(\ccmd[1]_INST_0_i_7_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \ccmd[1]_INST_0_i_8 
       (.I0(ir[7]),
        .I1(ir[6]),
        .O(\ccmd[1]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h30D5300030003000)) 
    \ccmd[1]_INST_0_i_9 
       (.I0(rst_n_fl_reg_17),
        .I1(ir[7]),
        .I2(ir[10]),
        .I3(ir[11]),
        .I4(div_crdy),
        .I5(crdy),
        .O(\ccmd[1]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[2]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(ccmd[2]));
  LUT6 #(
    .INIT(64'hA8A008A0AAAAAAAA)) 
    \ccmd[2]_INST_0_i_1 
       (.I0(\ccmd[2]_INST_0_i_2_n_0 ),
        .I1(ir[11]),
        .I2(ir[13]),
        .I3(ir[12]),
        .I4(ir[14]),
        .I5(ccmd_2_sn_1),
        .O(\ccmd[2]_INST_0_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h00000000509E559E)) 
    \ccmd[2]_INST_0_i_10 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[6]),
        .I2(ir[9]),
        .I3(ir[7]),
        .I4(\stat[1]_i_10_0 ),
        .I5(\ccmd[2]_INST_0_i_16_n_0 ),
        .O(\ccmd[2]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF0FF7070F0FF7F7F)) 
    \ccmd[2]_INST_0_i_11 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(ir[7]),
        .I3(rst_n_fl_reg_17),
        .I4(\stat_reg[2]_12 [1]),
        .I5(ir[6]),
        .O(\ccmd[2]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h0220FFFFAAAAFFFF)) 
    \ccmd[2]_INST_0_i_12 
       (.I0(ir[9]),
        .I1(ir[5]),
        .I2(ir[7]),
        .I3(ir[4]),
        .I4(ir[10]),
        .I5(\ccmd[2]_INST_0_i_17_n_0 ),
        .O(\ccmd[2]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \ccmd[2]_INST_0_i_15 
       (.I0(ir[7]),
        .I1(ir[6]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(ir[3]),
        .I4(ir[2]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\ccmd[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hD000FFFFFFFFFFFF)) 
    \ccmd[2]_INST_0_i_16 
       (.I0(ir[7]),
        .I1(ir[6]),
        .I2(ir[9]),
        .I3(ir[5]),
        .I4(ir[8]),
        .I5(ir[11]),
        .O(\ccmd[2]_INST_0_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h27F7FF2F)) 
    \ccmd[2]_INST_0_i_17 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[6]),
        .I3(\stat_reg[2]_12 [1]),
        .I4(ir[3]),
        .O(\ccmd[2]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFF8A0000FF8AFF8A)) 
    \ccmd[2]_INST_0_i_2 
       (.I0(\ccmd[2]_INST_0_i_4_n_0 ),
        .I1(\ccmd[2]_INST_0_i_5_n_0 ),
        .I2(\ccmd[2]_INST_0_i_6_n_0 ),
        .I3(\ccmd[2]_INST_0_i_7_n_0 ),
        .I4(\ccmd[2]_INST_0_i_8_n_0 ),
        .I5(\ccmd[2]_INST_0_i_9_n_0 ),
        .O(\ccmd[2]_INST_0_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF55555554)) 
    \ccmd[2]_INST_0_i_4 
       (.I0(\ccmd[2]_INST_0_i_10_n_0 ),
        .I1(\ccmd[2]_INST_0_i_11_n_0 ),
        .I2(ir[11]),
        .I3(ir[8]),
        .I4(ir[9]),
        .I5(\ccmd[2]_INST_0_i_12_n_0 ),
        .O(\ccmd[2]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEF6F2FFF2F2F2)) 
    \ccmd[2]_INST_0_i_5 
       (.I0(ir[9]),
        .I1(ir[6]),
        .I2(\ccmd[2]_INST_0_i_2_1 ),
        .I3(ir[11]),
        .I4(ir[8]),
        .I5(ir[7]),
        .O(\ccmd[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBFAABFFFBAAABAAA)) 
    \ccmd[2]_INST_0_i_6 
       (.I0(ir[11]),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(ir[6]),
        .I3(ir[7]),
        .I4(ir[9]),
        .I5(ir[8]),
        .O(\ccmd[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF4F)) 
    \ccmd[2]_INST_0_i_7 
       (.I0(rst_n_fl_reg_17),
        .I1(\stat[1]_i_10_0 ),
        .I2(rst_n_fl_reg_20),
        .I3(\stat_reg[2]_12 [2]),
        .I4(ir[15]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\ccmd[2]_INST_0_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[2]_INST_0_i_8 
       (.I0(ir[14]),
        .I1(ir[13]),
        .I2(ir[11]),
        .I3(ir[12]),
        .O(\ccmd[2]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \ccmd[2]_INST_0_i_9 
       (.I0(\ccmd[2]_INST_0_i_2_0 ),
        .I1(ir[8]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(\ccmd[2]_INST_0_i_15_n_0 ),
        .I4(ir[1]),
        .I5(ir[15]),
        .O(\ccmd[2]_INST_0_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(ccmd[3]));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \ccmd[3]_INST_0_i_1 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\ccmd[3]_INST_0_i_2_n_0 ),
        .I3(\ccmd[3]_INST_0_i_3_n_0 ),
        .I4(\ccmd[3]_INST_0_i_4_n_0 ),
        .I5(\ccmd[3]_INST_0_i_5_n_0 ),
        .O(\ccmd[3]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_10 
       (.I0(ir[11]),
        .I1(ir[8]),
        .O(\ccmd[3]_INST_0_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \ccmd[3]_INST_0_i_11 
       (.I0(ir[13]),
        .I1(ir[2]),
        .I2(ir[14]),
        .O(\ccmd[3]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \ccmd[3]_INST_0_i_12 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[1]),
        .I3(ir[6]),
        .O(\ccmd[3]_INST_0_i_12_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_13 
       (.I0(ir[10]),
        .I1(ir[8]),
        .O(\ccmd[3]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFDFDFFF)) 
    \ccmd[3]_INST_0_i_15 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[10]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\ccmd[3]_INST_0_i_24_n_0 ),
        .O(\ccmd[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF6FFFFFFFFF)) 
    \ccmd[3]_INST_0_i_16 
       (.I0(ir[8]),
        .I1(ir[11]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(ir[9]),
        .I5(ir[10]),
        .O(\ccmd[3]_INST_0_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[3]_INST_0_i_17 
       (.I0(rst_n_fl_reg_17),
        .I1(ir[7]),
        .O(\ccmd[3]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_18 
       (.I0(ir[10]),
        .I1(ir[8]),
        .O(\ccmd[3]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[3]_INST_0_i_19 
       (.I0(ir[11]),
        .I1(\stat_reg[2]_12 [1]),
        .O(\ccmd[3]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h3333032233333322)) 
    \ccmd[3]_INST_0_i_2 
       (.I0(\ccmd[3]_INST_0_i_6_n_0 ),
        .I1(\ccmd[3]_INST_0_i_7_n_0 ),
        .I2(\ccmd[3]_INST_0_i_8_n_0 ),
        .I3(ir[11]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(ir[8]),
        .O(\ccmd[3]_INST_0_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \ccmd[3]_INST_0_i_20 
       (.I0(ir[9]),
        .I1(ir[6]),
        .I2(ir[7]),
        .O(\ccmd[3]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h9FFFFFFF)) 
    \ccmd[3]_INST_0_i_21 
       (.I0(ir[7]),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[4]),
        .I3(ir[9]),
        .I4(ir[10]),
        .O(\ccmd[3]_INST_0_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAAAABAAAAAAAAAAF)) 
    \ccmd[3]_INST_0_i_22 
       (.I0(\ccmd[3]_INST_0_i_25_n_0 ),
        .I1(\stat[1]_i_10_0 ),
        .I2(ir[10]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(ir[9]),
        .I5(ir[7]),
        .O(\ccmd[3]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \ccmd[3]_INST_0_i_23 
       (.I0(ir[7]),
        .I1(ir[8]),
        .O(\ccmd[3]_INST_0_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \ccmd[3]_INST_0_i_24 
       (.I0(ir[8]),
        .I1(ir[9]),
        .I2(ir[10]),
        .I3(div_crdy),
        .I4(crdy),
        .I5(rst_n_fl_reg_17),
        .O(\ccmd[3]_INST_0_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000088400000080)) 
    \ccmd[3]_INST_0_i_25 
       (.I0(ir[3]),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(ir[6]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\bcmd[3]_INST_0_i_16_n_0 ),
        .I5(ir[7]),
        .O(\ccmd[3]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \ccmd[3]_INST_0_i_3 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(ir[10]),
        .I2(\ccmd[3]_INST_0_i_9_n_0 ),
        .I3(\bcmd[1]_INST_0_i_1_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(\ccmd[3]_INST_0_i_11_n_0 ),
        .O(\ccmd[3]_INST_0_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEBF)) 
    \ccmd[3]_INST_0_i_4 
       (.I0(\ccmd[3]_INST_0_i_12_n_0 ),
        .I1(\stat_reg[2]_12 [1]),
        .I2(ir[0]),
        .I3(ir[3]),
        .I4(ir[15]),
        .I5(ir[12]),
        .O(\ccmd[3]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0808800000888000)) 
    \ccmd[3]_INST_0_i_5 
       (.I0(ir[15]),
        .I1(\iv_reg[0] ),
        .I2(ir[12]),
        .I3(ir[13]),
        .I4(ir[14]),
        .I5(ir[11]),
        .O(\ccmd[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFDFFFDFFFFF0000)) 
    \ccmd[3]_INST_0_i_6 
       (.I0(\ccmd[3]_INST_0_i_13_n_0 ),
        .I1(\stat[1]_i_10_0 ),
        .I2(ir[7]),
        .I3(ir[9]),
        .I4(\ccmd[3]_INST_0_i_15_n_0 ),
        .I5(\stat_reg[2]_12 [0]),
        .O(\ccmd[3]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F4444444444444)) 
    \ccmd[3]_INST_0_i_7 
       (.I0(\ccmd[3]_INST_0_i_16_n_0 ),
        .I1(\ccmd[3]_INST_0_i_17_n_0 ),
        .I2(\ccmd[3]_INST_0_i_18_n_0 ),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\ccmd[3]_INST_0_i_19_n_0 ),
        .I5(\ccmd[3]_INST_0_i_20_n_0 ),
        .O(\ccmd[3]_INST_0_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF40000510)) 
    \ccmd[3]_INST_0_i_8 
       (.I0(\ccmd[3]_INST_0_i_21_n_0 ),
        .I1(ir[3]),
        .I2(ir[5]),
        .I3(ir[6]),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\ccmd[3]_INST_0_i_22_n_0 ),
        .O(\ccmd[3]_INST_0_i_8_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[3]_INST_0_i_9 
       (.I0(ir[9]),
        .I1(ir[7]),
        .O(\ccmd[3]_INST_0_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h282A282800000000)) 
    \ccmd[4]_INST_0 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\stat_reg[2]_12 [0]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(ir[10]),
        .I4(\ccmd[4]_INST_0_i_2_n_0 ),
        .I5(\ccmd[4]_INST_0_i_3_n_0 ),
        .O(\stat_reg[0]_3 ));
  LUT5 #(
    .INIT(32'h00001000)) 
    \ccmd[4]_INST_0_i_1 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(crdy),
        .I3(div_crdy),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\ccmd[4]_INST_0_i_1_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \ccmd[4]_INST_0_i_2 
       (.I0(ir[9]),
        .I1(ir[8]),
        .O(\ccmd[4]_INST_0_i_2_n_0 ));
  LUT5 #(
    .INIT(32'h00400000)) 
    \ccmd[4]_INST_0_i_3 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(ir[13]),
        .I2(ir[12]),
        .I3(ir[15]),
        .I4(ir[14]),
        .O(\ccmd[4]_INST_0_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hDFFF)) 
    \ccmd[4]_INST_0_i_4 
       (.I0(ir[14]),
        .I1(ir[15]),
        .I2(ir[12]),
        .I3(ir[13]),
        .O(\ccmd[4]_INST_0_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020000002)) 
    ctl_fetch_ext_fl_i_1
       (.I0(ctl_fetch_ext_fl_i_2_n_0),
        .I1(ctl_fetch_ext_fl_i_3_n_0),
        .I2(ir[10]),
        .I3(ir[8]),
        .I4(ir[9]),
        .I5(ctl_fetch_ext_fl_i_4_n_0),
        .O(ctl_fetch_ext));
  LUT6 #(
    .INIT(64'h0F0F000000000018)) 
    ctl_fetch_ext_fl_i_2
       (.I0(\stat_reg[2]_12 [2]),
        .I1(ir[0]),
        .I2(ir[3]),
        .I3(\bdatw[9]_INST_0_i_20_n_0 ),
        .I4(ir[8]),
        .I5(ir[6]),
        .O(ctl_fetch_ext_fl_i_2_n_0));
  LUT5 #(
    .INIT(32'hFFFE3FFE)) 
    ctl_fetch_ext_fl_i_3
       (.I0(\stat_reg[2]_12 [0]),
        .I1(ir[11]),
        .I2(ir[10]),
        .I3(ir[12]),
        .I4(\stat_reg[2]_12 [2]),
        .O(ctl_fetch_ext_fl_i_3_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFF7E)) 
    ctl_fetch_ext_fl_i_4
       (.I0(ir[14]),
        .I1(ir[13]),
        .I2(ir[12]),
        .I3(ctl_fetch_ext_fl_i_5_n_0),
        .I4(\stat_reg[2]_12 [1]),
        .I5(ir[15]),
        .O(ctl_fetch_ext_fl_i_4_n_0));
  LUT3 #(
    .INIT(8'hFE)) 
    ctl_fetch_ext_fl_i_5
       (.I0(ir[4]),
        .I1(ir[5]),
        .I2(ir[7]),
        .O(ctl_fetch_ext_fl_i_5_n_0));
  FDRE ctl_fetch_ext_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_ext),
        .Q(ctl_fetch_ext_fl),
        .R(\<const0> ));
  FDRE ctl_fetch_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(ctl_fetch_fl_reg_0),
        .Q(ctl_fetch_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h00000000FFFFFF54)) 
    ctl_fetch_inferred_i_1
       (.I0(ctl_fetch_inferred_i_2_n_0),
        .I1(ctl_fetch_fl_reg_1),
        .I2(ctl_fetch_inferred_i_4_n_0),
        .I3(ctl_fetch_inferred_i_5_n_0),
        .I4(ctl_fetch_inferred_i_6_n_0),
        .I5(ctl_fetch_inferred_i_7_n_0),
        .O(in0));
  LUT3 #(
    .INIT(8'h40)) 
    ctl_fetch_inferred_i_10
       (.I0(ir[10]),
        .I1(div_crdy),
        .I2(crdy),
        .O(div_crdy_reg_1));
  LUT6 #(
    .INIT(64'h22A222A222A2A2A2)) 
    ctl_fetch_inferred_i_11
       (.I0(\stat[0]_i_12_n_0 ),
        .I1(ctl_fetch_inferred_i_22_n_0),
        .I2(rst_n_fl_reg_17),
        .I3(ir[12]),
        .I4(ir[10]),
        .I5(ir[8]),
        .O(ctl_fetch_inferred_i_11_n_0));
  LUT5 #(
    .INIT(32'h88888088)) 
    ctl_fetch_inferred_i_12
       (.I0(ctl_fetch_inferred_i_23_n_0),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[6]),
        .I3(ir[10]),
        .I4(ir[8]),
        .O(ctl_fetch_inferred_i_12_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch_inferred_i_13
       (.I0(ir[14]),
        .I1(\sr_reg[13] [5]),
        .O(ctl_fetch_inferred_i_13_n_0));
  LUT6 #(
    .INIT(64'hBABABABBBABABABA)) 
    ctl_fetch_inferred_i_14
       (.I0(ctl_fetch_inferred_i_24_n_0),
        .I1(ctl_fetch_inferred_i_5_0),
        .I2(ctl_fetch_inferred_i_17_n_0),
        .I3(ctl_fetch_inferred_i_26_n_0),
        .I4(ctl_fetch_inferred_i_27_n_0),
        .I5(ctl_fetch_inferred_i_28_n_0),
        .O(ctl_fetch_inferred_i_14_n_0));
  LUT6 #(
    .INIT(64'h0E000E000E000000)) 
    ctl_fetch_inferred_i_15
       (.I0(ctl_fetch_inferred_i_29_n_0),
        .I1(ir[12]),
        .I2(\stat[0]_i_12_n_0 ),
        .I3(\iv_reg[0] ),
        .I4(ctl_fetch_inferred_i_6_0),
        .I5(ctl_fetch_inferred_i_31_n_0),
        .O(ctl_fetch_inferred_i_15_n_0));
  LUT6 #(
    .INIT(64'hC0CC000088888888)) 
    ctl_fetch_inferred_i_16
       (.I0(\sr_reg[13] [6]),
        .I1(ir[13]),
        .I2(\bcmd[3]_INST_0_i_16_n_0 ),
        .I3(\bcmd[3] ),
        .I4(ctl_fetch_inferred_i_32_n_0),
        .I5(ir[12]),
        .O(ctl_fetch_inferred_i_16_n_0));
  LUT2 #(
    .INIT(4'h7)) 
    ctl_fetch_inferred_i_17
       (.I0(ir[13]),
        .I1(ir[12]),
        .O(ctl_fetch_inferred_i_17_n_0));
  LUT6 #(
    .INIT(64'hAABABABAAABAAAAA)) 
    ctl_fetch_inferred_i_18
       (.I0(ctl_fetch_inferred_i_33_n_0),
        .I1(ctl_fetch_inferred_i_34_n_0),
        .I2(\ccmd[4]_INST_0_i_3_n_0 ),
        .I3(ctl_fetch_inferred_i_35_n_0),
        .I4(ctl_fetch_inferred_i_36_n_0),
        .I5(ctl_fetch_inferred_i_37_n_0),
        .O(ctl_fetch_inferred_i_18_n_0));
  LUT2 #(
    .INIT(4'hE)) 
    ctl_fetch_inferred_i_19
       (.I0(ir[7]),
        .I1(ir[3]),
        .O(ctl_fetch_inferred_i_19_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFF82A8)) 
    ctl_fetch_inferred_i_2
       (.I0(\bcmd[3]_INST_0_i_2_n_0 ),
        .I1(ir[0]),
        .I2(ir[1]),
        .I3(ir[3]),
        .I4(ir[9]),
        .I5(ctl_fetch_inferred_i_8_n_0),
        .O(ctl_fetch_inferred_i_2_n_0));
  LUT3 #(
    .INIT(8'h40)) 
    ctl_fetch_inferred_i_20
       (.I0(ir[3]),
        .I1(ir[6]),
        .I2(ir[8]),
        .O(ctl_fetch_inferred_i_20_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFEFA)) 
    ctl_fetch_inferred_i_21
       (.I0(ctl_fetch_inferred_i_38_n_0),
        .I1(\stat_reg[2]_12 [2]),
        .I2(ir[15]),
        .I3(ir[1]),
        .I4(ir[3]),
        .I5(ctl_fetch_inferred_i_39_n_0),
        .O(ctl_fetch_inferred_i_21_n_0));
  LUT6 #(
    .INIT(64'hFF0BFFFFFFBBFFFF)) 
    ctl_fetch_inferred_i_22
       (.I0(ir[7]),
        .I1(ir[9]),
        .I2(\sr_reg[13] [10]),
        .I3(ir[8]),
        .I4(ir[10]),
        .I5(ctl_fetch_inferred_i_11_0),
        .O(ctl_fetch_inferred_i_22_n_0));
  LUT6 #(
    .INIT(64'h7D00FFFFFFFFFFFF)) 
    ctl_fetch_inferred_i_23
       (.I0(ir[10]),
        .I1(ir[5]),
        .I2(ir[4]),
        .I3(ir[9]),
        .I4(ctl_fetch_inferred_i_41_n_0),
        .I5(ctl_fetch_inferred_i_42_n_0),
        .O(ctl_fetch_inferred_i_23_n_0));
  LUT4 #(
    .INIT(16'h0800)) 
    ctl_fetch_inferred_i_24
       (.I0(\sr_reg[13] [7]),
        .I1(ir[12]),
        .I2(ir[14]),
        .I3(ir[13]),
        .O(ctl_fetch_inferred_i_24_n_0));
  LUT6 #(
    .INIT(64'hEB00FFFF00000000)) 
    ctl_fetch_inferred_i_26
       (.I0(ctl_fetch_inferred_i_44_n_0),
        .I1(ir[3]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(ir[9]),
        .I4(ir[10]),
        .I5(ir[6]),
        .O(ctl_fetch_inferred_i_26_n_0));
  LUT6 #(
    .INIT(64'h1F0F00FFFFFFFFFF)) 
    ctl_fetch_inferred_i_27
       (.I0(ir[6]),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(ir[8]),
        .I3(ir[10]),
        .I4(ir[9]),
        .I5(ir[14]),
        .O(ctl_fetch_inferred_i_27_n_0));
  LUT6 #(
    .INIT(64'hAAFC0000FFFFFFFF)) 
    ctl_fetch_inferred_i_28
       (.I0(ir[6]),
        .I1(\sr_reg[13] [8]),
        .I2(\sr_reg[13] [10]),
        .I3(ir[9]),
        .I4(ir[8]),
        .I5(ctl_fetch_inferred_i_45_n_0),
        .O(ctl_fetch_inferred_i_28_n_0));
  LUT6 #(
    .INIT(64'h5101550555055505)) 
    ctl_fetch_inferred_i_29
       (.I0(ir[13]),
        .I1(\bcmd[3]_INST_0_i_12_n_0 ),
        .I2(ir[14]),
        .I3(\sr_reg[13] [5]),
        .I4(\bcmd[0]_INST_0_i_7_n_0 ),
        .I5(ctl_fetch_inferred_i_46_n_0),
        .O(ctl_fetch_inferred_i_29_n_0));
  LUT4 #(
    .INIT(16'hFF4F)) 
    ctl_fetch_inferred_i_31
       (.I0(ir[14]),
        .I1(\sr_reg[13] [4]),
        .I2(ir[12]),
        .I3(ir[13]),
        .O(ctl_fetch_inferred_i_31_n_0));
  LUT6 #(
    .INIT(64'hE0EEE0EEE0EEE0E0)) 
    ctl_fetch_inferred_i_32
       (.I0(ctl_fetch_inferred_i_47_n_0),
        .I1(ir[8]),
        .I2(rst_n_fl_reg_17),
        .I3(\stat[1]_i_10_0 ),
        .I4(\ccmd[1]_INST_0_i_17_n_0 ),
        .I5(\stat_reg[2]_12 [0]),
        .O(ctl_fetch_inferred_i_32_n_0));
  LUT6 #(
    .INIT(64'h00000000000000EA)) 
    ctl_fetch_inferred_i_33
       (.I0(ctl_fetch_inferred_i_48_n_0),
        .I1(\bcmd[3]_INST_0_i_10_n_0 ),
        .I2(\stat[1]_i_9_n_0 ),
        .I3(ir[12]),
        .I4(\bcmd[1]_INST_0_i_1_n_0 ),
        .I5(\ccmd[3]_INST_0_i_11_n_0 ),
        .O(ctl_fetch_inferred_i_33_n_0));
  LUT6 #(
    .INIT(64'hF7F7F7FF007700FF)) 
    ctl_fetch_inferred_i_34
       (.I0(\ccmd[3]_INST_0_i_13_n_0 ),
        .I1(ir[7]),
        .I2(ir[6]),
        .I3(ir[9]),
        .I4(ir[11]),
        .I5(\stat_reg[2]_12 [1]),
        .O(ctl_fetch_inferred_i_34_n_0));
  LUT3 #(
    .INIT(8'h2D)) 
    ctl_fetch_inferred_i_35
       (.I0(ir[4]),
        .I1(ir[7]),
        .I2(ir[5]),
        .O(ctl_fetch_inferred_i_35_n_0));
  LUT4 #(
    .INIT(16'h8000)) 
    ctl_fetch_inferred_i_36
       (.I0(ir[6]),
        .I1(ir[10]),
        .I2(ir[8]),
        .I3(ir[11]),
        .O(ctl_fetch_inferred_i_36_n_0));
  LUT6 #(
    .INIT(64'h0777007770777077)) 
    ctl_fetch_inferred_i_37
       (.I0(ctl_fetch_inferred_i_49_n_0),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[10]),
        .I3(ir[9]),
        .I4(ir[8]),
        .I5(ir[11]),
        .O(ctl_fetch_inferred_i_37_n_0));
  LUT6 #(
    .INIT(64'hFFFEFFFEFAFEFFFE)) 
    ctl_fetch_inferred_i_38
       (.I0(ctl_fetch_inferred_i_21_0),
        .I1(ir[2]),
        .I2(ir[6]),
        .I3(ir[9]),
        .I4(ir[14]),
        .I5(\stat_reg[2]_12 [2]),
        .O(ctl_fetch_inferred_i_38_n_0));
  LUT6 #(
    .INIT(64'hFFFFEEFEAAAAAAAA)) 
    ctl_fetch_inferred_i_39
       (.I0(ctl_fetch_inferred_i_51_n_0),
        .I1(ctl_fetch_inferred_i_17_n_0),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[7]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(ir[9]),
        .O(ctl_fetch_inferred_i_39_n_0));
  LUT6 #(
    .INIT(64'h00000000FFFFBAAA)) 
    ctl_fetch_inferred_i_4
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[8]),
        .I2(ir[9]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(ctl_fetch_inferred_i_11_n_0),
        .I5(ctl_fetch_fl_reg_2),
        .O(ctl_fetch_inferred_i_4_n_0));
  LUT6 #(
    .INIT(64'h4040F0F0F0F0F000)) 
    ctl_fetch_inferred_i_41
       (.I0(ir[5]),
        .I1(ir[3]),
        .I2(ir[8]),
        .I3(\sr_reg[13] [10]),
        .I4(ir[9]),
        .I5(ir[7]),
        .O(ctl_fetch_inferred_i_41_n_0));
  LUT5 #(
    .INIT(32'hFFFFF7FF)) 
    ctl_fetch_inferred_i_42
       (.I0(div_crdy),
        .I1(crdy),
        .I2(ir[9]),
        .I3(ir[7]),
        .I4(\sr_reg[13] [9]),
        .O(ctl_fetch_inferred_i_42_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch_inferred_i_44
       (.I0(ir[7]),
        .I1(ir[5]),
        .O(ctl_fetch_inferred_i_44_n_0));
  LUT2 #(
    .INIT(4'h2)) 
    ctl_fetch_inferred_i_45
       (.I0(ir[10]),
        .I1(ir[7]),
        .O(ctl_fetch_inferred_i_45_n_0));
  LUT5 #(
    .INIT(32'hFF0FF7F0)) 
    ctl_fetch_inferred_i_46
       (.I0(ctl_fetch_inferred_i_29_0),
        .I1(irq),
        .I2(ir[3]),
        .I3(ir[0]),
        .I4(ir[1]),
        .O(ctl_fetch_inferred_i_46_n_0));
  LUT6 #(
    .INIT(64'h0008000000080008)) 
    ctl_fetch_inferred_i_47
       (.I0(\stat_reg[2]_12 [0]),
        .I1(ir[7]),
        .I2(ir[9]),
        .I3(\stat[1]_i_10_0 ),
        .I4(\sr_reg[13] [9]),
        .I5(rst_n_fl_reg_17),
        .O(ctl_fetch_inferred_i_47_n_0));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    ctl_fetch_inferred_i_48
       (.I0(ctl_fetch_inferred_i_53_n_0),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(ctl_fetch_inferred_i_48_n_0));
  LUT3 #(
    .INIT(8'hA6)) 
    ctl_fetch_inferred_i_49
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[8]),
        .O(ctl_fetch_inferred_i_49_n_0));
  LUT6 #(
    .INIT(64'h8A8AAA8AAAAAAAAA)) 
    ctl_fetch_inferred_i_5
       (.I0(ir[11]),
        .I1(ctl_fetch_inferred_i_12_n_0),
        .I2(\stat_reg[0]_10 ),
        .I3(ctl_fetch_inferred_i_13_n_0),
        .I4(ir[12]),
        .I5(ctl_fetch_inferred_i_14_n_0),
        .O(ctl_fetch_inferred_i_5_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFF00FFFFFE)) 
    ctl_fetch_inferred_i_51
       (.I0(ir[4]),
        .I1(ir[5]),
        .I2(ir[7]),
        .I3(ir[9]),
        .I4(ir[10]),
        .I5(ir[8]),
        .O(ctl_fetch_inferred_i_51_n_0));
  LUT2 #(
    .INIT(4'h1)) 
    ctl_fetch_inferred_i_53
       (.I0(ir[7]),
        .I1(ir[6]),
        .O(ctl_fetch_inferred_i_53_n_0));
  LUT6 #(
    .INIT(64'h00000000EEEEEEE0)) 
    ctl_fetch_inferred_i_6
       (.I0(ctl_fetch_inferred_i_15_n_0),
        .I1(ctl_fetch_inferred_i_16_n_0),
        .I2(ctl_fetch_inferred_i_17_n_0),
        .I3(ir[14]),
        .I4(\sr_reg[13] [7]),
        .I5(ir[11]),
        .O(ctl_fetch_inferred_i_6_n_0));
  LUT6 #(
    .INIT(64'h0000222022202220)) 
    ctl_fetch_inferred_i_7
       (.I0(ctl_fetch_inferred_i_18_n_0),
        .I1(brdy),
        .I2(ctl_fetch_inferred_i_19_n_0),
        .I3(ir[9]),
        .I4(ctl_fetch_inferred_i_20_n_0),
        .I5(\stat_reg[2]_12 [0]),
        .O(ctl_fetch_inferred_i_7_n_0));
  LUT6 #(
    .INIT(64'hFFFFFFFFF2220000)) 
    ctl_fetch_inferred_i_8
       (.I0(ir[9]),
        .I1(rst_n_fl_reg_17),
        .I2(ir[1]),
        .I3(\stat_reg[2]_12 [1]),
        .I4(\stat_reg[2]_12 [0]),
        .I5(ctl_fetch_inferred_i_21_n_0),
        .O(ctl_fetch_inferred_i_8_n_0));
  LUT6 #(
    .INIT(64'h8000FFFF80000000)) 
    dctl_sign_f_i_1
       (.I0(\stat_reg[0] ),
        .I1(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_0 ),
        .I4(div_crdy),
        .I5(dctl_sign_f),
        .O(dctl_sign));
  LUT4 #(
    .INIT(16'hFF7F)) 
    \dctl_stat[2]_i_2 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_2 ),
        .O(\stat_reg[2]_4 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[1]_i_1 
       (.I0(irq_vec[0]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(eir[1]),
        .O(\eir_fl[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[2]_i_1 
       (.I0(irq_vec[1]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(eir[2]),
        .O(\eir_fl[2]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hFD)) 
    \eir_fl[31]_i_1 
       (.I0(rst_n),
        .I1(ctl_fetch_fl_reg_0),
        .I2(\eir_fl[31]_i_2_n_0 ),
        .O(\eir_fl[31]_i_1_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000400000)) 
    \eir_fl[31]_i_2 
       (.I0(\eir_fl_reg[31]_1 ),
        .I1(\eir_fl[31]_i_4_n_0 ),
        .I2(\fch_irq_lev[1]_i_5_n_0 ),
        .I3(ir[6]),
        .I4(\eir_fl[31]_i_5_n_0 ),
        .I5(\eir_fl_reg[31]_0 ),
        .O(\eir_fl[31]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \eir_fl[31]_i_4 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[3]),
        .O(\eir_fl[31]_i_4_n_0 ));
  LUT5 #(
    .INIT(32'h00010000)) 
    \eir_fl[31]_i_5 
       (.I0(ir[12]),
        .I1(ir[15]),
        .I2(ir[13]),
        .I3(ir[14]),
        .I4(ir[0]),
        .O(\eir_fl[31]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[3]_i_1 
       (.I0(irq_vec[2]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(eir[3]),
        .O(\eir_fl[3]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[4]_i_1 
       (.I0(irq_vec[3]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(eir[4]),
        .O(\eir_fl[4]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[5]_i_1 
       (.I0(irq_vec[4]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(eir[5]),
        .O(\eir_fl[5]_i_1_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \eir_fl[6]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(rst_n),
        .O(eir_fl0));
  LUT3 #(
    .INIT(8'hB8)) 
    \eir_fl[6]_i_2 
       (.I0(irq_vec[5]),
        .I1(\eir_fl[31]_i_2_n_0 ),
        .I2(eir[6]),
        .O(\eir_fl[6]_i_2_n_0 ));
  FDRE \eir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[0]),
        .Q(\eir_fl_reg_n_0_[0] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[10]),
        .Q(\eir_fl_reg_n_0_[10] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[11]),
        .Q(\eir_fl_reg_n_0_[11] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[12]),
        .Q(\eir_fl_reg_n_0_[12] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[13]),
        .Q(\eir_fl_reg_n_0_[13] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[14]),
        .Q(\eir_fl_reg_n_0_[14] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[15]),
        .Q(\eir_fl_reg_n_0_[15] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[16]),
        .Q(\eir_fl_reg_n_0_[16] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[17]),
        .Q(\eir_fl_reg_n_0_[17] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[18]),
        .Q(\eir_fl_reg_n_0_[18] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[19]),
        .Q(\eir_fl_reg_n_0_[19] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[1]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[1] ),
        .R(eir_fl0));
  FDRE \eir_fl_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[20]),
        .Q(\eir_fl_reg_n_0_[20] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[21]),
        .Q(\eir_fl_reg_n_0_[21] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[22]),
        .Q(\eir_fl_reg_n_0_[22] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[23]),
        .Q(\eir_fl_reg_n_0_[23] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[24]),
        .Q(\eir_fl_reg_n_0_[24] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[25]),
        .Q(\eir_fl_reg_n_0_[25] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[26]),
        .Q(\eir_fl_reg_n_0_[26] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[27]),
        .Q(\eir_fl_reg_n_0_[27] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[28]),
        .Q(\eir_fl_reg_n_0_[28] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[29]),
        .Q(\eir_fl_reg_n_0_[29] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[2]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[2] ),
        .R(eir_fl0));
  FDRE \eir_fl_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[30]),
        .Q(\eir_fl_reg_n_0_[30] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[31]),
        .Q(\eir_fl_reg_n_0_[31] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[3]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[3] ),
        .R(eir_fl0));
  FDRE \eir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[4]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[4] ),
        .R(eir_fl0));
  FDRE \eir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[5]_i_1_n_0 ),
        .Q(\eir_fl_reg_n_0_[5] ),
        .R(eir_fl0));
  FDRE \eir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\eir_fl[6]_i_2_n_0 ),
        .Q(\eir_fl_reg_n_0_[6] ),
        .R(eir_fl0));
  FDRE \eir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[7]),
        .Q(\eir_fl_reg_n_0_[7] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[8]),
        .Q(\eir_fl_reg_n_0_[8] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  FDRE \eir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(eir[9]),
        .Q(\eir_fl_reg_n_0_[9] ),
        .R(\eir_fl[31]_i_1_n_0 ));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_1
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[31] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[15] ),
        .O(eir[31]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_10
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[22] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[6] ),
        .O(eir[22]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_11
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[21] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[5] ),
        .O(eir[21]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_12
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[20] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[4] ),
        .O(eir[20]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_13
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[19] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[3] ),
        .O(eir[19]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_14
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[18] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[2] ),
        .O(eir[18]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_15
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[17] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[1] ),
        .O(eir[17]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_16
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[16] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[0] ),
        .O(eir[16]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_17
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[15] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[15]),
        .O(eir[15]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_18
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[14] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[14]),
        .O(eir[14]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_19
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[13] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[13]),
        .O(eir[13]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_2
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[30] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[14] ),
        .O(eir[30]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_20
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[12] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[12]),
        .O(eir[12]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_21
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[11] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[11]),
        .O(eir[11]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_22
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[10] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[10]),
        .O(eir[10]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_23
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[9] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[9]),
        .O(eir[9]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_24
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[8] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[8]),
        .O(eir[8]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_25
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[7] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[7]),
        .O(eir[7]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_26
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[6] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[6]),
        .O(eir[6]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_27
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[5] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[5]),
        .O(eir[5]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_28
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[4] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[4]),
        .O(eir[4]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_29
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[3] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[3]),
        .O(eir[3]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_3
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[29] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[13] ),
        .O(eir[29]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_30
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[2] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[2]),
        .O(eir[2]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_31
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[1] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[1]),
        .O(eir[1]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_32
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[0] ),
        .I2(ctl_fetch_ext_fl),
        .I3(fdat[0]),
        .O(eir[0]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_4
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[28] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[12] ),
        .O(eir[28]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_5
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[27] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[11] ),
        .O(eir[27]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_6
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[26] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[10] ),
        .O(eir[26]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_7
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[25] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[9] ),
        .O(eir[25]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_8
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[24] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[8] ),
        .O(eir[24]));
  LUT4 #(
    .INIT(16'hA808)) 
    eir_inferred_i_9
       (.I0(rst_n_fl),
        .I1(\eir_fl_reg_n_0_[23] ),
        .I2(ctl_fetch_ext_fl),
        .I3(\eir_fl_reg_n_0_[7] ),
        .O(eir[23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[0]_i_1 
       (.I0(irq_lev[0]),
        .I1(fch_irq_lev0),
        .I2(fch_irq_lev[0]),
        .O(\fch_irq_lev[0]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \fch_irq_lev[1]_i_1 
       (.I0(irq_lev[1]),
        .I1(fch_irq_lev0),
        .I2(fch_irq_lev[1]),
        .O(\fch_irq_lev[1]_i_1_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \fch_irq_lev[1]_i_2 
       (.I0(\fch_irq_lev[1]_i_3_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(ir[0]),
        .I3(\fch_irq_lev[1]_i_5_n_0 ),
        .I4(\eir_fl_reg[31]_0 ),
        .O(fch_irq_lev0));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \fch_irq_lev[1]_i_3 
       (.I0(\fch_irq_lev[1]_i_2_0 ),
        .I1(\stat_reg[0]_10 ),
        .I2(ir[3]),
        .I3(ir[4]),
        .I4(ir[6]),
        .I5(ir[5]),
        .O(\fch_irq_lev[1]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \fch_irq_lev[1]_i_4 
       (.I0(ir[14]),
        .I1(ir[13]),
        .I2(ir[15]),
        .I3(ir[12]),
        .O(\fch_irq_lev[1]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \fch_irq_lev[1]_i_5 
       (.I0(\ccmd[1]_INST_0_i_17_n_0 ),
        .I1(ir[8]),
        .I2(ir[7]),
        .I3(brdy),
        .I4(ir[1]),
        .I5(ir[2]),
        .O(\fch_irq_lev[1]_i_5_n_0 ));
  FDRE \fch_irq_lev_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[0]_i_1_n_0 ),
        .Q(fch_irq_lev[0]),
        .R(p_0_in));
  FDRE \fch_irq_lev_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\fch_irq_lev[1]_i_1_n_0 ),
        .Q(fch_irq_lev[1]),
        .R(p_0_in));
  FDRE fch_irq_req_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(fch_irq_req),
        .Q(fch_irq_req_fl),
        .R(\<const0> ));
  LUT6 #(
    .INIT(64'h0000000001010001)) 
    \grn[15]_i_1__11 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\stat_reg[2]_7 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_3 ));
  LUT6 #(
    .INIT(64'h0101010000000000)) 
    \grn[15]_i_1__12 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\stat_reg[2]_7 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_4 ));
  LUT6 #(
    .INIT(64'h0000000001010100)) 
    \grn[15]_i_1__13 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\stat_reg[2]_7 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_5 ));
  LUT6 #(
    .INIT(64'h0101000100000000)) 
    \grn[15]_i_1__14 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .I2(\stat_reg[2]_7 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_6 ));
  LUT6 #(
    .INIT(64'h0404000400000000)) 
    \grn[15]_i_1__15 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_7 ));
  LUT6 #(
    .INIT(64'h0000000004040400)) 
    \grn[15]_i_1__16 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_8 ));
  LUT6 #(
    .INIT(64'h0404040000000000)) 
    \grn[15]_i_1__17 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_9 ));
  LUT6 #(
    .INIT(64'h0000000004040004)) 
    \grn[15]_i_1__18 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[0]),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_10 ));
  LUT6 #(
    .INIT(64'h0404000400000000)) 
    \grn[15]_i_1__19 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_11 ));
  LUT6 #(
    .INIT(64'h0000000004040400)) 
    \grn[15]_i_1__20 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_12 ));
  LUT6 #(
    .INIT(64'h0404040000000000)) 
    \grn[15]_i_1__21 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_13 ));
  LUT6 #(
    .INIT(64'h0000000004040004)) 
    \grn[15]_i_1__22 
       (.I0(\stat_reg[2]_7 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_14 ));
  LUT6 #(
    .INIT(64'h0404000400000000)) 
    \grn[15]_i_1__23 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_15 ));
  LUT6 #(
    .INIT(64'h0000000004040400)) 
    \grn[15]_i_1__24 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_16 ));
  LUT6 #(
    .INIT(64'h0404040000000000)) 
    \grn[15]_i_1__25 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_17 ));
  LUT6 #(
    .INIT(64'h0000000004040004)) 
    \grn[15]_i_1__26 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(\iv[15]_i_6_n_0 ),
        .I2(ctl_selc_rn[1]),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_18 ));
  LUT6 #(
    .INIT(64'h4040004000000000)) 
    \grn[15]_i_1__27 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_19 ));
  LUT6 #(
    .INIT(64'h0000000040404000)) 
    \grn[15]_i_1__28 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_20 ));
  LUT6 #(
    .INIT(64'h4040400000000000)) 
    \grn[15]_i_1__29 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_21 ));
  LUT6 #(
    .INIT(64'h0202000200000000)) 
    \grn[15]_i_1__3 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\stat_reg[2]_9 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(E));
  LUT6 #(
    .INIT(64'h0000000040400040)) 
    \grn[15]_i_1__30 
       (.I0(\grn[15]_i_2__0_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_22 ));
  LUT6 #(
    .INIT(64'h0000000002020200)) 
    \grn[15]_i_1__4 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\stat_reg[2]_9 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h0202020000000000)) 
    \grn[15]_i_1__5 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\stat_reg[2]_9 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_1 ));
  LUT6 #(
    .INIT(64'h0000000002020002)) 
    \grn[15]_i_1__6 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .I2(\stat_reg[2]_9 ),
        .I3(\sr_reg[13] [1]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[13] [0]),
        .O(\sr_reg[1]_2 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \grn[15]_i_2 
       (.I0(\grn[15]_i_2__2_n_0 ),
        .I1(ctl_selc_rn[1]),
        .I2(ctl_selc_rn[0]),
        .I3(\iv[15]_i_6_n_0 ),
        .O(cbus_sel_0));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_2__0 
       (.I0(ctl_selc_rn[0]),
        .I1(\grn[15]_i_2__2_n_0 ),
        .O(\grn[15]_i_2__0_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \grn[15]_i_2__1 
       (.I0(\iv[15]_i_6_n_0 ),
        .I1(\grn[15]_i_2__2_n_0 ),
        .O(\stat_reg[2]_7 ));
  LUT2 #(
    .INIT(4'h7)) 
    \grn[15]_i_2__2 
       (.I0(ctl_selc[1]),
        .I1(ctl_selc[0]),
        .O(\grn[15]_i_2__2_n_0 ));
  FDRE \ir_fl_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[0]),
        .Q(ir_fl[0]),
        .R(p_0_in));
  FDRE \ir_fl_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[10]),
        .Q(ir_fl[10]),
        .R(p_0_in));
  FDRE \ir_fl_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[11]),
        .Q(ir_fl[11]),
        .R(p_0_in));
  FDRE \ir_fl_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[12]),
        .Q(ir_fl[12]),
        .R(p_0_in));
  FDRE \ir_fl_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[13]),
        .Q(ir_fl[13]),
        .R(p_0_in));
  FDRE \ir_fl_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[14]),
        .Q(ir_fl[14]),
        .R(p_0_in));
  FDRE \ir_fl_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[15]),
        .Q(ir_fl[15]),
        .R(p_0_in));
  FDRE \ir_fl_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[1]),
        .Q(ir_fl[1]),
        .R(p_0_in));
  FDRE \ir_fl_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[2]),
        .Q(ir_fl[2]),
        .R(p_0_in));
  FDRE \ir_fl_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[3]),
        .Q(ir_fl[3]),
        .R(p_0_in));
  FDRE \ir_fl_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[4]),
        .Q(ir_fl[4]),
        .R(p_0_in));
  FDRE \ir_fl_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[5]),
        .Q(ir_fl[5]),
        .R(p_0_in));
  FDRE \ir_fl_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[6]),
        .Q(ir_fl[6]),
        .R(p_0_in));
  FDRE \ir_fl_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[7]),
        .Q(ir_fl[7]),
        .R(p_0_in));
  FDRE \ir_fl_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[8]),
        .Q(ir_fl[8]),
        .R(p_0_in));
  FDRE \ir_fl_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(ir[9]),
        .Q(ir_fl[9]),
        .R(p_0_in));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_1
       (.I0(rst_n_fl),
        .I1(ir_fl[15]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[15]),
        .O(ir[15]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_10
       (.I0(rst_n_fl),
        .I1(ir_fl[6]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[6]),
        .O(ir[6]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_11
       (.I0(rst_n_fl),
        .I1(ir_fl[5]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[5]),
        .O(ir[5]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_12
       (.I0(rst_n_fl),
        .I1(ir_fl[4]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[4]),
        .O(ir[4]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_13
       (.I0(rst_n_fl),
        .I1(ir_fl[3]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[3]),
        .O(ir[3]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_14
       (.I0(rst_n_fl),
        .I1(ir_fl[2]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[2]),
        .O(ir[2]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_15
       (.I0(rst_n_fl),
        .I1(ir_fl[1]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[1]),
        .O(ir[1]));
  LUT5 #(
    .INIT(32'hA8A8A808)) 
    ir_inferred_i_16
       (.I0(rst_n_fl),
        .I1(ir_fl[0]),
        .I2(ctl_fetch_fl),
        .I3(fdat[0]),
        .I4(fch_irq_req_fl),
        .O(ir[0]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_2
       (.I0(rst_n_fl),
        .I1(ir_fl[14]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[14]),
        .O(ir[14]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_3
       (.I0(rst_n_fl),
        .I1(ir_fl[13]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[13]),
        .O(ir[13]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_4
       (.I0(rst_n_fl),
        .I1(ir_fl[12]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[12]),
        .O(ir[12]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_5
       (.I0(rst_n_fl),
        .I1(ir_fl[11]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[11]),
        .O(ir[11]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_6
       (.I0(rst_n_fl),
        .I1(ir_fl[10]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[10]),
        .O(ir[10]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_7
       (.I0(rst_n_fl),
        .I1(ir_fl[9]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[9]),
        .O(ir[9]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_8
       (.I0(rst_n_fl),
        .I1(ir_fl[8]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[8]),
        .O(ir[8]));
  LUT5 #(
    .INIT(32'h08A80808)) 
    ir_inferred_i_9
       (.I0(rst_n_fl),
        .I1(ir_fl[7]),
        .I2(ctl_fetch_fl),
        .I3(fch_irq_req_fl),
        .I4(fdat[7]),
        .O(ir[7]));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[0]_i_1 
       (.I0(\iv[0]_i_2_n_0 ),
        .I1(\iv[0]_i_3_n_0 ),
        .I2(\tr_reg[0]_3 ),
        .I3(\tr_reg[0]_4 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[0]),
        .O(cbus[0]));
  LUT6 #(
    .INIT(64'hAEEAEEAACC000000)) 
    \iv[0]_i_13 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\sr[6]_i_14_n_0 ),
        .I2(\stat_reg[0] ),
        .I3(\stat_reg[0]_0 ),
        .I4(abus_0[0]),
        .I5(\bdatw[5] [0]),
        .O(\iv[0]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[0]_i_15 
       (.I0(\sr_reg[8]_10 ),
        .I1(\iv[8]_i_34_0 ),
        .O(\iv[0]_i_27_0 ));
  LUT6 #(
    .INIT(64'hF0FFF000EEEEEEEE)) 
    \iv[0]_i_19 
       (.I0(\iv[8]_i_34_0 ),
        .I1(\iv[6]_i_8_0 ),
        .I2(\iv[0]_i_9 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\sr[4]_i_66_1 ),
        .I5(\stat_reg[0]_2 ),
        .O(\sr_reg[8]_35 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[0]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[0]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[0]),
        .I4(\iv[0]_i_6_n_0 ),
        .I5(\iv[0]_i_7_n_0 ),
        .O(\iv[0]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h80FF)) 
    \iv[0]_i_20 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr_reg[13] [6]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\bdatw[5] [1]),
        .O(\sr_reg[6]_3 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \iv[0]_i_27 
       (.I0(bbus_0[2]),
        .I1(abus_0[0]),
        .I2(\bdatw[8]_INST_0_i_1 ),
        .O(\iv[8]_i_34_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[0]_i_3 
       (.I0(\stat_reg[2]_2 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I2(\tr_reg[0]_0 ),
        .I3(\tr_reg[0]_1 ),
        .I4(\tr_reg[0]_2 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[0]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[0]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[3]_i_2_1 [0]),
        .I2(\tr[30]_i_2_0 [0]),
        .I3(div_crdy_reg),
        .I4(Q[0]),
        .I5(div_crdy_reg_0),
        .O(\iv[0]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[0]_i_7 
       (.I0(\sr[4]_i_7_3 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_1 ),
        .I2(\sr[4]_i_7_4 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[0]_i_13_n_0 ),
        .O(\iv[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[10]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[10]),
        .I2(bdatr[2]),
        .I3(\tr_reg[15]_3 ),
        .I4(\iv[10]_i_2_n_0 ),
        .I5(\iv[10]_i_3_n_0 ),
        .O(cbus[10]));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[10]_i_11 
       (.I0(\sr_reg[8]_33 ),
        .I1(\iv[10]_i_5 ),
        .O(\iv[10]_i_21 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[10]_i_15 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[10]_i_6_0 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr[4]_i_85_1 ),
        .O(\iv[10]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[10]_i_17 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\iv[10]_i_37_n_0 ),
        .O(\iv[10]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[10]_i_18 
       (.I0(\stat_reg[0]_2 ),
        .I1(bbus_0[8]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\stat_reg[2]_1 ),
        .I4(abus_0[10]),
        .O(\iv[10]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \iv[10]_i_19 
       (.I0(abus_0[2]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(bbus_0[8]),
        .I4(abus_0[10]),
        .I5(\stat_reg[0]_2 ),
        .O(\iv[10]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[10]_i_2 
       (.I0(\stat_reg[2]_2 ),
        .I1(\tr_reg[10]_0 ),
        .I2(\tr_reg[10]_1 ),
        .I3(\iv[10]_i_6_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[10]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[10]_i_20 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[8]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[10]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[10]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[10]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[10]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[10]),
        .I4(\iv[10]_i_7_n_0 ),
        .I5(\iv[10]_i_8_n_0 ),
        .O(\iv[10]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[10]_i_31 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[9]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_62 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[10]_i_36 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[9]),
        .I2(\sr_reg[13] [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\sr_reg[8]_61 ));
  LUT6 #(
    .INIT(64'h1DFF1D331D331DFF)) 
    \iv[10]_i_37 
       (.I0(abus_0[18]),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[1]),
        .I3(\stat_reg[0]_2 ),
        .I4(abus_0[10]),
        .I5(bbus_0[8]),
        .O(\iv[10]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[10]_i_6 
       (.I0(\iv[10]_i_15_n_0 ),
        .I1(\iv[10]_i_21 ),
        .I2(\iv[10]_i_2_0 ),
        .I3(\iv[10]_i_2_1 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\iv[10]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[10]_i_7 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[11]_i_3_0 [2]),
        .I2(\tr[30]_i_2_0 [10]),
        .I3(div_crdy_reg),
        .I4(Q[10]),
        .I5(div_crdy_reg_0),
        .O(\iv[10]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[10]_i_8 
       (.I0(\iv[10]_i_17_n_0 ),
        .I1(\iv[10]_i_18_n_0 ),
        .I2(\stat_reg[0] ),
        .I3(\iv[10]_i_19_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\iv[10]_i_20_n_0 ),
        .O(\iv[10]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[11]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[11]),
        .I2(bdatr[3]),
        .I3(\tr_reg[15]_3 ),
        .I4(\iv[11]_i_2_n_0 ),
        .I5(\iv[11]_i_3_n_0 ),
        .O(cbus[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[11]_i_17 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[10]),
        .O(\iv[11]_i_17_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[11]_i_18 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[11]_i_7_2 ),
        .I2(\sr_reg[8]_18 ),
        .I3(\iv[11]_i_7_0 ),
        .O(\iv[11]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'hDDDF)) 
    \iv[11]_i_19 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[6]_i_8_0 ),
        .I2(\iv[11]_i_7_1 ),
        .I3(\sr_reg[8]_11 ),
        .O(\iv[11]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[11]_i_2 
       (.I0(\stat_reg[2]_2 ),
        .I1(\tr_reg[11]_0 ),
        .I2(\tr_reg[11]_1 ),
        .I3(\tr_reg[11]_2 ),
        .I4(\iv[11]_i_7_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[11]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAFF3C00AA003C00)) 
    \iv[11]_i_20 
       (.I0(bbus_0[2]),
        .I1(abus_0[11]),
        .I2(bbus_0[9]),
        .I3(\stat_reg[0]_1 ),
        .I4(\stat_reg[0]_2 ),
        .I5(abus_0[19]),
        .O(\iv[11]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \iv[11]_i_21 
       (.I0(\stat_reg[0]_0 ),
        .I1(abus_0[11]),
        .I2(\stat_reg[2]_1 ),
        .I3(\sr[6]_i_32_n_0 ),
        .I4(bbus_0[9]),
        .I5(\stat_reg[0]_2 ),
        .O(\iv[11]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[11]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[11]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[11]),
        .I4(\iv[11]_i_8_n_0 ),
        .I5(\iv[11]_i_9_n_0 ),
        .O(\iv[11]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[11]_i_32 
       (.I0(\iv[11]_i_17_n_0 ),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_51 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[11]_i_39 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[9]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[11]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[11]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hEAEEEAEA)) 
    \iv[11]_i_40 
       (.I0(\tr[27]_i_5_1 ),
        .I1(\sr[6]_i_32_n_0 ),
        .I2(abus_0[11]),
        .I3(\stat_reg[0]_2 ),
        .I4(bbus_0[9]),
        .O(\iv[11]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[11]_i_7 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\iv[11]_i_17_n_0 ),
        .I3(\iv[14]_i_18_n_0 ),
        .I4(\iv[11]_i_18_n_0 ),
        .I5(\iv[11]_i_19_n_0 ),
        .O(\iv[11]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[11]_i_8 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[11]_i_3_0 [3]),
        .I2(\tr[30]_i_2_0 [11]),
        .I3(div_crdy_reg),
        .I4(Q[11]),
        .I5(div_crdy_reg_0),
        .O(\iv[11]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h20FFFFFF20FF0000)) 
    \iv[11]_i_9 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\iv[11]_i_20_n_0 ),
        .I3(\iv[11]_i_21_n_0 ),
        .I4(\stat_reg[0] ),
        .I5(\iv_reg[11]_i_22_n_0 ),
        .O(\iv[11]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[12]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[12]),
        .I2(bdatr[4]),
        .I3(\tr_reg[15]_3 ),
        .I4(\iv[12]_i_2_n_0 ),
        .I5(\iv[12]_i_3_n_0 ),
        .O(cbus[12]));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[12]_i_12 
       (.I0(\sr_reg[8]_33 ),
        .I1(\sr_reg[8]_9 ),
        .O(\iv[12]_i_22_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[12]_i_13 
       (.I0(\iv[12]_i_26_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\sr[4]_i_44_0 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\tr[20]_i_7 ),
        .I5(\iv[6]_i_8_0 ),
        .O(\sr_reg[8]_21 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[12]_i_15 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[12]_i_6_0 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr[4]_i_98 ),
        .O(\iv[12]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[12]_i_17 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\iv[12]_i_37_n_0 ),
        .O(\iv[12]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[12]_i_18 
       (.I0(\stat_reg[0]_2 ),
        .I1(bbus_0[10]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\stat_reg[2]_1 ),
        .I4(abus_0[12]),
        .O(\iv[12]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \iv[12]_i_19 
       (.I0(abus_0[4]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(bbus_0[10]),
        .I4(abus_0[12]),
        .I5(\stat_reg[0]_2 ),
        .O(\iv[12]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[12]_i_2 
       (.I0(\stat_reg[2]_2 ),
        .I1(\iv[12]_i_10 ),
        .I2(\tr_reg[12]_0 ),
        .I3(\iv[12]_i_6_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[12]_i_20 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[10]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[12]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[12]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hCFCACFCACFCAC5C0)) 
    \iv[12]_i_22 
       (.I0(\sr_reg[8]_13 ),
        .I1(\sr[4]_i_98 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\iv[4]_i_8 ),
        .I4(bbus_0[0]),
        .I5(\iv[4]_i_8_0 ),
        .O(\sr_reg[8]_9 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[12]_i_26 
       (.I0(\sr_reg[8]_13 ),
        .I1(\tr[28]_i_9_0 ),
        .O(\iv[12]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[12]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[12]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[12]),
        .I4(\iv[12]_i_7_n_0 ),
        .I5(\iv[12]_i_8_n_0 ),
        .O(\iv[12]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[12]_i_31 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[11]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_60 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[12]_i_36 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[11]),
        .I2(\sr_reg[13] [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\sr_reg[8]_59 ));
  LUT6 #(
    .INIT(64'h1DFF1D331D331DFF)) 
    \iv[12]_i_37 
       (.I0(abus_0[20]),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[3]),
        .I3(\stat_reg[0]_2 ),
        .I4(abus_0[12]),
        .I5(bbus_0[10]),
        .O(\iv[12]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[12]_i_4 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I1(\iv[12]_i_9_n_0 ),
        .I2(\sr[4]_i_20 ),
        .O(\iv[12]_i_10 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[12]_i_6 
       (.I0(\iv[12]_i_15_n_0 ),
        .I1(\iv[12]_i_22_0 ),
        .I2(\sr_reg[8]_21 ),
        .I3(\iv[12]_i_2_0 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\iv[12]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[12]_i_7 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[15]_i_9_0 [0]),
        .I2(\tr[30]_i_2_0 [12]),
        .I3(div_crdy_reg),
        .I4(Q[12]),
        .I5(div_crdy_reg_0),
        .O(\iv[12]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[12]_i_8 
       (.I0(\iv[12]_i_17_n_0 ),
        .I1(\iv[12]_i_18_n_0 ),
        .I2(\stat_reg[0] ),
        .I3(\iv[12]_i_19_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\iv[12]_i_20_n_0 ),
        .O(\iv[12]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[12]_i_9 
       (.I0(\sr_reg[8]_7 ),
        .I1(abus_0[31]),
        .I2(\iv[12]_i_4_0 ),
        .I3(\iv[12]_i_4_1 ),
        .I4(\sr_reg[8]_9 ),
        .I5(\sr_reg[8]_10 ),
        .O(\iv[12]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[13]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[13]),
        .I2(bdatr[5]),
        .I3(\tr_reg[15]_3 ),
        .I4(\iv[13]_i_2_n_0 ),
        .I5(\iv[13]_i_3_n_0 ),
        .O(cbus[13]));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[13]_i_12 
       (.I0(\sr_reg[8]_33 ),
        .I1(\iv[13]_i_5 ),
        .O(\iv[13]_i_23 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[13]_i_13 
       (.I0(\iv[13]_i_28_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\sr[4]_i_45_0 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\tr[21]_i_7 ),
        .I5(\iv[6]_i_8_0 ),
        .O(\sr_reg[8]_20 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[13]_i_15 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[13]_i_6_0 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\iv[13]_i_6_1 ),
        .O(\iv[13]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[13]_i_17 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\iv[13]_i_8_0 ),
        .O(\iv[13]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[13]_i_18 
       (.I0(\stat_reg[0]_2 ),
        .I1(bbus_0[11]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\stat_reg[2]_1 ),
        .I4(abus_0[13]),
        .O(\iv[13]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \iv[13]_i_19 
       (.I0(abus_0[5]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(abus_0[13]),
        .I4(\stat_reg[0]_2 ),
        .I5(bbus_0[11]),
        .O(\iv[13]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[13]_i_2 
       (.I0(\stat_reg[2]_2 ),
        .I1(\tr_reg[13]_0 ),
        .I2(\tr_reg[13]_1 ),
        .I3(\iv[13]_i_6_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[13]_i_20 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[11]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[13]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[13]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[13]_i_28 
       (.I0(\sr_reg[8]_13 ),
        .I1(\tr[29]_i_7 ),
        .O(\iv[13]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[13]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[13]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[13]),
        .I4(\iv[13]_i_7_n_0 ),
        .I5(\iv[13]_i_8_n_0 ),
        .O(\iv[13]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[13]_i_33 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[12]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_58 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[13]_i_38 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[12]),
        .I2(\sr_reg[13] [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\sr_reg[8]_57 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[13]_i_6 
       (.I0(\iv[13]_i_15_n_0 ),
        .I1(\iv[13]_i_23 ),
        .I2(\sr_reg[8]_20 ),
        .I3(\iv[13]_i_2_0 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\iv[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[13]_i_7 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[15]_i_9_0 [1]),
        .I2(\tr[30]_i_2_0 [13]),
        .I3(div_crdy_reg),
        .I4(Q[13]),
        .I5(div_crdy_reg_0),
        .O(\iv[13]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[13]_i_8 
       (.I0(\iv[13]_i_17_n_0 ),
        .I1(\iv[13]_i_18_n_0 ),
        .I2(\stat_reg[0] ),
        .I3(\iv[13]_i_19_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\iv[13]_i_20_n_0 ),
        .O(\iv[13]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[14]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[14]),
        .I2(bdatr[6]),
        .I3(\tr_reg[15]_3 ),
        .I4(\iv[14]_i_2_n_0 ),
        .I5(\iv[14]_i_3_n_0 ),
        .O(cbus[14]));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[14]_i_13 
       (.I0(\iv[14]_i_28_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\sr[4]_i_80 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\tr[22]_i_7_0 ),
        .I5(\iv[6]_i_8_0 ),
        .O(\sr_reg[8]_23 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[14]_i_17 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[13]),
        .O(\iv[14]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAA00000002)) 
    \iv[14]_i_18 
       (.I0(bbus_0[3]),
        .I1(bbus_0[1]),
        .I2(bbus_0[0]),
        .I3(\bdatw[5] [0]),
        .I4(bbus_0[2]),
        .I5(\iv[0]_i_21 ),
        .O(\iv[14]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[14]_i_19 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[14]_i_7_1 ),
        .I2(\sr_reg[8]_18 ),
        .I3(\iv[14]_i_7_2 ),
        .O(\iv[14]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[14]_i_2 
       (.I0(\stat_reg[2]_2 ),
        .I1(\tr_reg[14]_0 ),
        .I2(\tr_reg[14]_1 ),
        .I3(\iv[14]_i_6_n_0 ),
        .I4(\iv[14]_i_7_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[14]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hDDDF)) 
    \iv[14]_i_20 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[6]_i_8_0 ),
        .I2(\iv[14]_i_7_0 ),
        .I3(\sr_reg[8]_11 ),
        .O(\iv[14]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hAAFF3C00AA003C00)) 
    \iv[14]_i_21 
       (.I0(bbus_0[4]),
        .I1(abus_0[14]),
        .I2(bbus_0[12]),
        .I3(\stat_reg[0]_1 ),
        .I4(\stat_reg[0]_2 ),
        .I5(abus_0[22]),
        .O(\iv[14]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \iv[14]_i_22 
       (.I0(\stat_reg[0]_0 ),
        .I1(abus_0[14]),
        .I2(\stat_reg[2]_1 ),
        .I3(\sr[6]_i_32_n_0 ),
        .I4(bbus_0[12]),
        .I5(\stat_reg[0]_2 ),
        .O(\iv[14]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[14]_i_28 
       (.I0(\sr_reg[8]_13 ),
        .I1(\tr[30]_i_8 ),
        .O(\iv[14]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[14]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[14]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[14]),
        .I4(\iv[14]_i_8_n_0 ),
        .I5(\iv[14]_i_9_n_0 ),
        .O(\iv[14]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h8F)) 
    \iv[14]_i_31 
       (.I0(\sr_reg[13] [8]),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\stat_reg[0]_2 ),
        .O(\sr_reg[8]_44 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[14]_i_33 
       (.I0(\iv[14]_i_17_n_0 ),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_48 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \iv[14]_i_34 
       (.I0(bbus_0[2]),
        .I1(\bdatw[5] [0]),
        .I2(bbus_0[0]),
        .I3(bbus_0[1]),
        .O(\bdatw[10]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h565656AAAA56AAAA)) 
    \iv[14]_i_37 
       (.I0(bbus_0[1]),
        .I1(\bdatw[5] [0]),
        .I2(bbus_0[0]),
        .I3(\sr_reg[13] [8]),
        .I4(bbus_0[3]),
        .I5(\bdatw[5] [1]),
        .O(\sr_reg[8]_18 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[14]_i_40 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[12]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[14]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[14]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hF222F2F2F222F222)) 
    \iv[14]_i_41 
       (.I0(abus_0[6]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(abus_0[14]),
        .I4(\stat_reg[0]_2 ),
        .I5(bbus_0[12]),
        .O(\iv[14]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[14]_i_6 
       (.I0(\sr_reg[8]_23 ),
        .I1(bbus_0[3]),
        .I2(\iv[14]_i_2_0 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\iv[6]_i_8_0 ),
        .I5(\iv[14]_i_2_1 ),
        .O(\iv[14]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[14]_i_7 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\iv[14]_i_17_n_0 ),
        .I3(\iv[14]_i_18_n_0 ),
        .I4(\iv[14]_i_19_n_0 ),
        .I5(\iv[14]_i_20_n_0 ),
        .O(\iv[14]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[14]_i_8 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[15]_i_9_0 [2]),
        .I2(Q[14]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [14]),
        .I5(div_crdy_reg),
        .O(\iv[14]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h20FFFFFF20FF0000)) 
    \iv[14]_i_9 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\iv[14]_i_21_n_0 ),
        .I3(\iv[14]_i_22_n_0 ),
        .I4(\stat_reg[0] ),
        .I5(\iv_reg[14]_i_23_n_0 ),
        .O(\iv[14]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \iv[15]_i_1 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\stat_reg[2]_9 ),
        .I3(\iv[15]_i_6_n_0 ),
        .O(\stat_reg[2]_0 [1]));
  LUT6 #(
    .INIT(64'h000000000000FF04)) 
    \iv[15]_i_10 
       (.I0(\iv[15]_i_29_n_0 ),
        .I1(\iv[15]_i_30_n_0 ),
        .I2(\iv[15]_i_31_n_0 ),
        .I3(\iv[15]_i_32_n_0 ),
        .I4(\iv[15]_i_33_n_0 ),
        .I5(\stat_reg[2]_12 [0]),
        .O(\iv[15]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h04)) 
    \iv[15]_i_100 
       (.I0(\bdatw[8]_INST_0_i_1 ),
        .I1(abus_0[31]),
        .I2(bbus_0[2]),
        .O(\iv[15]_i_100_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_107 
       (.I0(bbus_0[13]),
        .I1(acmd),
        .O(\iv[15]_i_107_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \iv[15]_i_108 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(acmd),
        .O(\stat_reg[2]_1 ));
  LUT6 #(
    .INIT(64'hFF66F0000066F000)) 
    \iv[15]_i_109 
       (.I0(abus_0[15]),
        .I1(bbus_0[13]),
        .I2(abus_0[23]),
        .I3(\stat_reg[0]_2 ),
        .I4(\stat_reg[0]_1 ),
        .I5(bbus_0[5]),
        .O(\iv[15]_i_109_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000007F)) 
    \iv[15]_i_11 
       (.I0(\iv[15]_i_34_n_0 ),
        .I1(\iv[15]_i_35_n_0 ),
        .I2(ir[10]),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\iv[15]_i_36_n_0 ),
        .I5(\iv[15]_i_37_n_0 ),
        .O(\iv[15]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[15]_i_111 
       (.I0(acmd),
        .I1(bbus_0[5]),
        .I2(\stat_reg[0]_2 ),
        .O(\iv[15]_i_111_n_0 ));
  LUT6 #(
    .INIT(64'hFEFEFFFFEAEAFFFB)) 
    \iv[15]_i_112 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[10]),
        .I2(ir[9]),
        .I3(\sr_reg[13] [8]),
        .I4(ir[11]),
        .I5(ir[7]),
        .O(\iv[15]_i_112_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F0000D2C)) 
    \iv[15]_i_113 
       (.I0(ir[4]),
        .I1(ir[7]),
        .I2(ir[5]),
        .I3(ir[3]),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\iv[15]_i_158_n_0 ),
        .O(\iv[15]_i_113_n_0 ));
  LUT6 #(
    .INIT(64'hBBB7BBBA55555555)) 
    \iv[15]_i_114 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(ir[7]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[3]),
        .I5(ir[10]),
        .O(\iv[15]_i_114_n_0 ));
  LUT6 #(
    .INIT(64'h0000AABAFFFFFFFF)) 
    \iv[15]_i_115 
       (.I0(\ccmd[3]_INST_0_i_18_n_0 ),
        .I1(\iv[15]_i_159_n_0 ),
        .I2(\stat_reg[2]_12 [0]),
        .I3(\bcmd[0]_INST_0_i_12_n_0 ),
        .I4(ir[7]),
        .I5(ir[9]),
        .O(\iv[15]_i_115_n_0 ));
  LUT6 #(
    .INIT(64'h43334333C333F333)) 
    \iv[15]_i_116 
       (.I0(\stat[1]_i_10_0 ),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[8]),
        .I3(ir[10]),
        .I4(\sr_reg[13] [8]),
        .I5(ir[7]),
        .O(\iv[15]_i_116_n_0 ));
  LUT6 #(
    .INIT(64'hBABBABBBBABBBBBB)) 
    \iv[15]_i_117 
       (.I0(\stat[0]_i_15_n_0 ),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[8]),
        .I3(ir[7]),
        .I4(ir[9]),
        .I5(ir[6]),
        .O(\iv[15]_i_117_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA0000AAAA0C00)) 
    \iv[15]_i_118 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\iv[15]_i_73_n_0 ),
        .I2(ir[8]),
        .I3(ir[10]),
        .I4(\stat_reg[2]_12 [0]),
        .I5(ir[9]),
        .O(\iv[15]_i_118_n_0 ));
  LUT6 #(
    .INIT(64'hA22AA2222A22A222)) 
    \iv[15]_i_12 
       (.I0(\bcmd[1]_INST_0_i_1_n_0 ),
        .I1(\iv_reg[0] ),
        .I2(ir[12]),
        .I3(ir[14]),
        .I4(ir[11]),
        .I5(ir[13]),
        .O(\iv[15]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hEFEF0000FFFFF0FF)) 
    \iv[15]_i_120 
       (.I0(ir[3]),
        .I1(ctl_fetch_ext_fl_i_5_n_0),
        .I2(ir[6]),
        .I3(ir[7]),
        .I4(ir[9]),
        .I5(ir[8]),
        .O(\iv[15]_i_120_n_0 ));
  LUT6 #(
    .INIT(64'hAAEAAAAAEAEAEAEA)) 
    \iv[15]_i_121 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(ir[10]),
        .I2(\ccmd[3]_INST_0_i_10_n_0 ),
        .I3(ir[6]),
        .I4(ir[7]),
        .I5(ir[9]),
        .O(\iv[15]_i_121_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000FFFE)) 
    \iv[15]_i_122 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[15]),
        .I2(ir[14]),
        .I3(\iv[15]_i_160_n_0 ),
        .I4(\iv[15]_i_161_n_0 ),
        .I5(\iv[15]_i_162_n_0 ),
        .O(\iv[15]_i_122_n_0 ));
  LUT4 #(
    .INIT(16'hA959)) 
    \iv[15]_i_123 
       (.I0(ir[11]),
        .I1(\sr_reg[13] [4]),
        .I2(ir[13]),
        .I3(\sr_reg[13] [7]),
        .O(\iv[15]_i_123_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \iv[15]_i_124 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[8]),
        .O(\iv[15]_i_124_n_0 ));
  LUT3 #(
    .INIT(8'h01)) 
    \iv[15]_i_125 
       (.I0(\sr_reg[13] [8]),
        .I1(ir[7]),
        .I2(ir[8]),
        .O(\iv[15]_i_125_n_0 ));
  LUT5 #(
    .INIT(32'hFFFBBBBB)) 
    \iv[15]_i_126 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(ir[7]),
        .I3(ir[8]),
        .I4(ir[9]),
        .O(\iv[15]_i_126_n_0 ));
  LUT6 #(
    .INIT(64'h0000000020222020)) 
    \iv[15]_i_13 
       (.I0(\iv[15]_i_38_n_0 ),
        .I1(\stat_reg[2]_12 [2]),
        .I2(\iv[15]_i_39_n_0 ),
        .I3(rst_n_fl_reg_17),
        .I4(ir[9]),
        .I5(\iv[15]_i_40_n_0 ),
        .O(\iv[15]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[15]_i_14 
       (.I0(ir[12]),
        .I1(ir[11]),
        .O(\iv[15]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \iv[15]_i_15 
       (.I0(\iv[15]_i_41_n_0 ),
        .I1(\fch_irq_lev[1]_i_4_n_0 ),
        .I2(ir[7]),
        .I3(ir[3]),
        .I4(ir[9]),
        .I5(\iv[15]_i_42_n_0 ),
        .O(\iv[15]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \iv[15]_i_158 
       (.I0(ir[8]),
        .I1(ir[10]),
        .I2(ir[6]),
        .O(\iv[15]_i_158_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \iv[15]_i_159 
       (.I0(ir[6]),
        .I1(ir[3]),
        .O(\iv[15]_i_159_n_0 ));
  LUT6 #(
    .INIT(64'h08080808AA080808)) 
    \iv[15]_i_16 
       (.I0(\iv[15]_i_43_n_0 ),
        .I1(ir[5]),
        .I2(\iv[15]_i_44_n_0 ),
        .I3(ir[10]),
        .I4(ir[11]),
        .I5(\iv[15]_i_45_n_0 ),
        .O(\iv[15]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFF4B0000FF4BFF4B)) 
    \iv[15]_i_160 
       (.I0(\sr_reg[13] [6]),
        .I1(ir[13]),
        .I2(ir[11]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\iv[15]_i_173_n_0 ),
        .I5(\iv[15]_i_41_n_0 ),
        .O(\iv[15]_i_160_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \iv[15]_i_161 
       (.I0(ir[8]),
        .I1(ir[10]),
        .I2(ir[11]),
        .I3(ir[5]),
        .I4(\iv[15]_i_174_n_0 ),
        .I5(\iv[15]_i_175_n_0 ),
        .O(\iv[15]_i_161_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA008200800080)) 
    \iv[15]_i_162 
       (.I0(\iv[15]_i_122_0 ),
        .I1(ir[11]),
        .I2(\sr_reg[13] [5]),
        .I3(ir[13]),
        .I4(ir[15]),
        .I5(ir[14]),
        .O(\iv[15]_i_162_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000EFBF)) 
    \iv[15]_i_17 
       (.I0(\iv[15]_i_46_n_0 ),
        .I1(ir[11]),
        .I2(ir[10]),
        .I3(ir[9]),
        .I4(\iv[15]_i_47_n_0 ),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\iv[15]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF723FFFFF)) 
    \iv[15]_i_173 
       (.I0(ir[0]),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[1]),
        .I3(ir[3]),
        .I4(ctl_fetch_inferred_i_53_n_0),
        .I5(\iv[15]_i_176_n_0 ),
        .O(\iv[15]_i_173_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEA)) 
    \iv[15]_i_174 
       (.I0(ir[6]),
        .I1(ir[1]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[4]),
        .I4(ir[15]),
        .I5(\iv[15]_i_177_n_0 ),
        .O(\iv[15]_i_174_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEFFF)) 
    \iv[15]_i_175 
       (.I0(ir[3]),
        .I1(ir[7]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(ir[0]),
        .I4(ir[9]),
        .I5(ir[13]),
        .O(\iv[15]_i_175_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[15]_i_176 
       (.I0(ir[9]),
        .I1(ir[13]),
        .O(\iv[15]_i_176_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[15]_i_177 
       (.I0(ir[14]),
        .I1(ir[2]),
        .O(\iv[15]_i_177_n_0 ));
  LUT6 #(
    .INIT(64'hE0EE0000FFFFFFFF)) 
    \iv[15]_i_18 
       (.I0(\iv[15]_i_48_n_0 ),
        .I1(ir[15]),
        .I2(\tr[31]_i_6_n_0 ),
        .I3(ir[10]),
        .I4(\iv[15]_i_49_n_0 ),
        .I5(\iv[15]_i_122_0 ),
        .O(\iv[15]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_19 
       (.I0(acmd),
        .I1(\stat_reg[0]_1 ),
        .O(\stat_reg[2]_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[15]_i_2 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[15]),
        .I2(bdatr[7]),
        .I3(\tr_reg[15]_3 ),
        .I4(\sr_reg[8] ),
        .I5(\iv[15]_i_9_n_0 ),
        .O(cbus[15]));
  LUT3 #(
    .INIT(8'h02)) 
    \iv[15]_i_20 
       (.I0(\stat_reg[0] ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_2 ),
        .O(\niho_dsp_a[32]_INST_0_i_7_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_24 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0] ),
        .O(\niho_dsp_a[15]_INST_0_i_2_0 ));
  LUT4 #(
    .INIT(16'hF7FF)) 
    \iv[15]_i_25 
       (.I0(\stat_reg[0] ),
        .I1(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\stat_reg[0]_1 ),
        .O(\iv[15]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'hD5)) 
    \iv[15]_i_26 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I1(mul_rslt),
        .I2(\sr_reg[13] [8]),
        .O(\iv[15]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[15]_i_27 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[15]_i_9_0 [3]),
        .I2(Q[15]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [15]),
        .I5(div_crdy_reg),
        .O(\iv[15]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0DFDFCFC0D0D0)) 
    \iv[15]_i_28 
       (.I0(\iv[15]_i_67_n_0 ),
        .I1(\iv[15]_i_68_n_0 ),
        .I2(\stat_reg[0] ),
        .I3(\iv[15]_i_69_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\iv[15]_i_70_n_0 ),
        .O(\iv[15]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hDD55DD55D151D114)) 
    \iv[15]_i_29 
       (.I0(ir[4]),
        .I1(ir[6]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(ir[7]),
        .I4(ir[3]),
        .I5(ir[5]),
        .O(\iv[15]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF8A88)) 
    \iv[15]_i_3 
       (.I0(rst_n_fl_reg_20),
        .I1(\iv[15]_i_10_n_0 ),
        .I2(\iv[15]_i_11_n_0 ),
        .I3(\iv_reg[0]_1 ),
        .I4(ir[15]),
        .I5(\iv[15]_i_12_n_0 ),
        .O(ctl_selc[0]));
  LUT3 #(
    .INIT(8'h80)) 
    \iv[15]_i_30 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(ir[9]),
        .O(\iv[15]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0000DD00FD00FF00)) 
    \iv[15]_i_31 
       (.I0(ir[5]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(ir[3]),
        .I3(ir[4]),
        .I4(ir[6]),
        .I5(ir[7]),
        .O(\iv[15]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF0F0F444)) 
    \iv[15]_i_32 
       (.I0(\iv[15]_i_71_n_0 ),
        .I1(\ccmd[3]_INST_0_i_20_n_0 ),
        .I2(\iv[15]_i_72_n_0 ),
        .I3(\iv[15]_i_73_n_0 ),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\iv[15]_i_74_n_0 ),
        .O(\iv[15]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00000000D5FFFDFF)) 
    \iv[15]_i_33 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[9]),
        .I2(ir[11]),
        .I3(ir[10]),
        .I4(\iv[15]_i_75_n_0 ),
        .I5(\iv[15]_i_76_n_0 ),
        .O(\iv[15]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'h1800555500005555)) 
    \iv[15]_i_34 
       (.I0(ir[7]),
        .I1(ir[5]),
        .I2(ir[4]),
        .I3(ir[6]),
        .I4(ir[9]),
        .I5(\iv[15]_i_77_n_0 ),
        .O(\iv[15]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_35 
       (.I0(ir[11]),
        .I1(ir[8]),
        .O(\iv[15]_i_35_n_0 ));
  LUT6 #(
    .INIT(64'h00000F0022000000)) 
    \iv[15]_i_36 
       (.I0(brdy),
        .I1(ir[6]),
        .I2(\stat[1]_i_10_0 ),
        .I3(\iv[15]_i_35_n_0 ),
        .I4(ir[9]),
        .I5(ir[10]),
        .O(\iv[15]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h2222222202000000)) 
    \iv[15]_i_37 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(\iv[15]_i_78_n_0 ),
        .I3(brdy),
        .I4(\bcmd[1]_INST_0_i_5_n_0 ),
        .I5(\iv[15]_i_79_n_0 ),
        .O(\iv[15]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FF0D)) 
    \iv[15]_i_38 
       (.I0(\iv[15]_i_80_n_0 ),
        .I1(\iv[15]_i_81_n_0 ),
        .I2(\iv[15]_i_13_0 ),
        .I3(\iv[15]_i_82_n_0 ),
        .I4(\badr[31]_INST_0_i_9_n_0 ),
        .I5(\iv[15]_i_83_n_0 ),
        .O(\iv[15]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFD0)) 
    \iv[15]_i_39 
       (.I0(ir[1]),
        .I1(ir[14]),
        .I2(\iv[15]_i_84_n_0 ),
        .I3(\iv[15]_i_85_n_0 ),
        .I4(ir[8]),
        .I5(brdy),
        .O(\iv[15]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAAAEAEA)) 
    \iv[15]_i_4 
       (.I0(\iv[15]_i_13_n_0 ),
        .I1(ir[15]),
        .I2(\iv_reg[0] ),
        .I3(\iv[15]_i_14_n_0 ),
        .I4(ir[13]),
        .I5(\iv[15]_i_15_n_0 ),
        .O(ctl_selc[1]));
  LUT6 #(
    .INIT(64'h4040404040404044)) 
    \iv[15]_i_40 
       (.I0(brdy),
        .I1(\stat_reg[2]_12 [0]),
        .I2(\iv[15]_i_86_n_0 ),
        .I3(\bcmd[3]_INST_0_i_13_n_0 ),
        .I4(ir[14]),
        .I5(\stat_reg[2]_12 [1]),
        .O(\iv[15]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \iv[15]_i_41 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(ir[8]),
        .I3(ir[4]),
        .I4(ir[5]),
        .I5(ir[2]),
        .O(\iv[15]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFDFFFFFFFFF)) 
    \iv[15]_i_42 
       (.I0(ir[0]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(\stat_reg[2]_12 [2]),
        .I3(ir[6]),
        .I4(ir[1]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\iv[15]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008000)) 
    \iv[15]_i_43 
       (.I0(ir[12]),
        .I1(ir[13]),
        .I2(ir[14]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(ir[15]),
        .O(\iv[15]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h000000000000EFFF)) 
    \iv[15]_i_44 
       (.I0(\iv[15]_i_78_n_0 ),
        .I1(ir[10]),
        .I2(\iv[15]_i_35_n_0 ),
        .I3(brdy),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\iv[15]_i_37_n_0 ),
        .O(\iv[15]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFFFFFDDDDFFFF)) 
    \iv[15]_i_45 
       (.I0(ir[5]),
        .I1(\iv[15]_i_87_n_0 ),
        .I2(\iv[15]_i_88_n_0 ),
        .I3(\bdatw[12]_INST_0_i_23_n_0 ),
        .I4(ir[8]),
        .I5(ir[9]),
        .O(\iv[15]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h7777F0FF7777FFFF)) 
    \iv[15]_i_46 
       (.I0(ir[2]),
        .I1(\iv[15]_i_72_n_0 ),
        .I2(\iv[15]_i_89_n_0 ),
        .I3(brdy),
        .I4(ir[8]),
        .I5(ir[7]),
        .O(\iv[15]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h08FF080800000000)) 
    \iv[15]_i_47 
       (.I0(\iv[15]_i_90_n_0 ),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(ir[3]),
        .I3(\stat[1]_i_19_n_0 ),
        .I4(\ccmd[3]_INST_0_i_10_n_0 ),
        .I5(ir[2]),
        .O(\iv[15]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFEFFFFFFFFFFFF)) 
    \iv[15]_i_48 
       (.I0(\ccmd[2]_INST_0_i_8_n_0 ),
        .I1(ir[10]),
        .I2(\tr[31]_i_22_n_0 ),
        .I3(ir[2]),
        .I4(ir[3]),
        .I5(\bcmd[3]_INST_0_i_13_n_0 ),
        .O(\iv[15]_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hABAAABAB)) 
    \iv[15]_i_49 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\iv[15]_i_91_n_0 ),
        .I2(\iv[15]_i_92_n_0 ),
        .I3(\iv[15]_i_93_n_0 ),
        .I4(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\iv[15]_i_49_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \iv[15]_i_5 
       (.I0(ctl_selc_rn[1]),
        .I1(ctl_selc_rn[0]),
        .O(\stat_reg[2]_9 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_50 
       (.I0(\bdatw[12]_INST_0_i_1_0 ),
        .I1(\sr_reg[13] [8]),
        .O(\sr_reg[8]_45 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[15]_i_57 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[14]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\iv[15]_i_22 ),
        .O(\sr_reg[8]_56 ));
  LUT6 #(
    .INIT(64'h5151514040405140)) 
    \iv[15]_i_58 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\iv[15]_i_100_n_0 ),
        .I3(\tr[23]_i_3 ),
        .I4(\sr_reg[8]_11 ),
        .I5(\iv[15]_i_22_0 ),
        .O(\sr_reg[8]_43 ));
  LUT6 #(
    .INIT(64'hBAAABABABAAAAAAA)) 
    \iv[15]_i_59 
       (.I0(\bdatw[12]_INST_0_i_1_0 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\stat_reg[0]_2 ),
        .I3(\iv[15]_i_22_0 ),
        .I4(\sr_reg[8]_11 ),
        .I5(\tr[23]_i_3 ),
        .O(\sr_reg[8]_17 ));
  LUT6 #(
    .INIT(64'h4445444455555555)) 
    \iv[15]_i_6 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\iv[15]_i_16_n_0 ),
        .I2(\iv[15]_i_17_n_0 ),
        .I3(\ccmd[4]_INST_0_i_4_n_0 ),
        .I4(\iv_reg[0]_0 ),
        .I5(\iv[15]_i_18_n_0 ),
        .O(\iv[15]_i_6_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[15]_i_63 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[14]),
        .I2(\sr[4]_i_66_0 ),
        .I3(bbus_0[3]),
        .O(\sr_reg[8]_55 ));
  LUT4 #(
    .INIT(16'h7FFF)) 
    \iv[15]_i_65 
       (.I0(\stat_reg[2]_2 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\stat_reg[0]_2 ),
        .I3(div_crdy),
        .O(div_crdy_reg_0));
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \iv[15]_i_66 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\stat_reg[0]_0 ),
        .I3(div_crdy),
        .I4(acmd),
        .I5(\stat_reg[0] ),
        .O(div_crdy_reg));
  LUT5 #(
    .INIT(32'h77007F7F)) 
    \iv[15]_i_67 
       (.I0(\iv[15]_i_107_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_2 ),
        .I3(\stat_reg[2]_1 ),
        .I4(abus_0[15]),
        .O(\iv[15]_i_67_n_0 ));
  LUT3 #(
    .INIT(8'h20)) 
    \iv[15]_i_68 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\iv[15]_i_109_n_0 ),
        .O(\iv[15]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'hEAFFEAEAEAEAEAEA)) 
    \iv[15]_i_69 
       (.I0(\iv[15]_i_28_0 ),
        .I1(\sr[6]_i_32_n_0 ),
        .I2(abus_0[15]),
        .I3(\stat_reg[0]_2 ),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_107_n_0 ),
        .O(\iv[15]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[15]_i_70 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[13]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[15]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[15]_i_70_n_0 ));
  LUT4 #(
    .INIT(16'hABBB)) 
    \iv[15]_i_71 
       (.I0(ir[11]),
        .I1(rst_n_fl_reg_17),
        .I2(crdy),
        .I3(div_crdy),
        .O(\iv[15]_i_71_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[15]_i_72 
       (.I0(ir[9]),
        .I1(ir[10]),
        .I2(ir[11]),
        .O(\iv[15]_i_72_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[15]_i_73 
       (.I0(ir[7]),
        .I1(\sr_reg[13] [8]),
        .O(\iv[15]_i_73_n_0 ));
  LUT5 #(
    .INIT(32'h55FF04FF)) 
    \iv[15]_i_74 
       (.I0(ir[10]),
        .I1(ir[6]),
        .I2(ir[9]),
        .I3(ir[8]),
        .I4(ir[7]),
        .O(\iv[15]_i_74_n_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[15]_i_75 
       (.I0(ir[6]),
        .I1(brdy),
        .I2(ir[7]),
        .O(\iv[15]_i_75_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC4044FFFFFFFF)) 
    \iv[15]_i_76 
       (.I0(ir[7]),
        .I1(ir[8]),
        .I2(ir[9]),
        .I3(ir[6]),
        .I4(ir[10]),
        .I5(\iv[15]_i_112_n_0 ),
        .O(\iv[15]_i_76_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_77 
       (.I0(ir[3]),
        .I1(brdy),
        .O(\iv[15]_i_77_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_78 
       (.I0(ir[6]),
        .I1(ir[9]),
        .O(\iv[15]_i_78_n_0 ));
  LUT5 #(
    .INIT(32'h10001111)) 
    \iv[15]_i_79 
       (.I0(ir[8]),
        .I1(ir[9]),
        .I2(crdy),
        .I3(div_crdy),
        .I4(ir[7]),
        .O(\iv[15]_i_79_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[15]_i_8 
       (.I0(\stat_reg[2]_2 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I2(\tr_reg[15]_0 ),
        .I3(\tr_reg[15]_1 ),
        .I4(\tr_reg[15]_2 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'h00FF45FFFFFF45FF)) 
    \iv[15]_i_80 
       (.I0(\iv[15]_i_113_n_0 ),
        .I1(\iv[15]_i_114_n_0 ),
        .I2(\bdatw[15]_INST_0_i_28_n_0 ),
        .I3(ir[11]),
        .I4(\iv[15]_i_115_n_0 ),
        .I5(\iv[15]_i_116_n_0 ),
        .O(\iv[15]_i_80_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF45455545)) 
    \iv[15]_i_81 
       (.I0(\iv[15]_i_117_n_0 ),
        .I1(\iv[15]_i_79_n_0 ),
        .I2(\stat_reg[2]_12 [0]),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(\iv[15]_i_78_n_0 ),
        .I5(\iv[15]_i_118_n_0 ),
        .O(\iv[15]_i_81_n_0 ));
  LUT6 #(
    .INIT(64'hE2E2E2E2222222E2)) 
    \iv[15]_i_82 
       (.I0(\iv[15]_i_38_0 ),
        .I1(ir[13]),
        .I2(\iv_reg[0]_0 ),
        .I3(\iv[15]_i_120_n_0 ),
        .I4(\ccmd[1]_INST_0_i_11_n_0 ),
        .I5(\iv[15]_i_121_n_0 ),
        .O(\iv[15]_i_82_n_0 ));
  LUT6 #(
    .INIT(64'h0C550C550C550055)) 
    \iv[15]_i_83 
       (.I0(\iv[15]_i_122_n_0 ),
        .I1(\iv[15]_i_122_0 ),
        .I2(ir[14]),
        .I3(ir[12]),
        .I4(ir[15]),
        .I5(\iv[15]_i_123_n_0 ),
        .O(\iv[15]_i_83_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[15]_i_84 
       (.I0(ir[9]),
        .I1(ir[11]),
        .O(\iv[15]_i_84_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_85 
       (.I0(ir[15]),
        .I1(\stat_reg[2]_12 [1]),
        .O(\iv[15]_i_85_n_0 ));
  LUT6 #(
    .INIT(64'hA8A828A82828A8A8)) 
    \iv[15]_i_86 
       (.I0(ir[9]),
        .I1(ir[11]),
        .I2(ir[10]),
        .I3(ir[4]),
        .I4(ir[7]),
        .I5(ir[5]),
        .O(\iv[15]_i_86_n_0 ));
  LUT3 #(
    .INIT(8'h2A)) 
    \iv[15]_i_87 
       (.I0(ir[7]),
        .I1(div_crdy),
        .I2(crdy),
        .O(\iv[15]_i_87_n_0 ));
  LUT5 #(
    .INIT(32'h3FB7FFFF)) 
    \iv[15]_i_88 
       (.I0(ir[4]),
        .I1(ir[6]),
        .I2(ir[5]),
        .I3(ir[7]),
        .I4(brdy),
        .O(\iv[15]_i_88_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_89 
       (.I0(ir[6]),
        .I1(ir[5]),
        .O(\iv[15]_i_89_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[15]_i_9 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[15]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[15]),
        .I4(\iv[15]_i_27_n_0 ),
        .I5(\iv[15]_i_28_n_0 ),
        .O(\iv[15]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080000000)) 
    \iv[15]_i_90 
       (.I0(ir[9]),
        .I1(ir[8]),
        .I2(ir[11]),
        .I3(ir[10]),
        .I4(ir[6]),
        .I5(ir[7]),
        .O(\iv[15]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h000000000FDD0F00)) 
    \iv[15]_i_91 
       (.I0(\iv[15]_i_124_n_0 ),
        .I1(\iv[15]_i_125_n_0 ),
        .I2(\bcmd[1]_INST_0_i_5_n_0 ),
        .I3(ir[9]),
        .I4(ir[5]),
        .I5(\stat[0]_i_15_n_0 ),
        .O(\iv[15]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'h444CFCFC44444444)) 
    \iv[15]_i_92 
       (.I0(\iv[15]_i_126_n_0 ),
        .I1(ir[5]),
        .I2(ir[7]),
        .I3(\sr_reg[13] [8]),
        .I4(ir[8]),
        .I5(\iv[15]_i_72_n_0 ),
        .O(\iv[15]_i_92_n_0 ));
  LUT6 #(
    .INIT(64'hF77FFF3FB77FFF7B)) 
    \iv[15]_i_93 
       (.I0(ir[7]),
        .I1(ir[2]),
        .I2(ir[6]),
        .I3(ir[5]),
        .I4(ir[4]),
        .I5(ir[3]),
        .O(\iv[15]_i_93_n_0 ));
  LUT6 #(
    .INIT(64'h5656565656565655)) 
    \iv[15]_i_96 
       (.I0(bbus_0[2]),
        .I1(\iv[0]_i_21 ),
        .I2(\iv[0]_i_21_0 ),
        .I3(bbus_0[1]),
        .I4(bbus_0[0]),
        .I5(\bdatw[5] [0]),
        .O(\sr_reg[8]_11 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[1]_i_1 
       (.I0(\iv[1]_i_2_n_0 ),
        .I1(\tr_reg[1]_0 ),
        .I2(\tr_reg[1]_1 ),
        .I3(\tr_reg[1]_2 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[1]),
        .O(cbus[1]));
  LUT5 #(
    .INIT(32'h47774744)) 
    \iv[1]_i_12 
       (.I0(bbus_0[0]),
        .I1(\stat_reg[0]_1 ),
        .I2(abus_0[9]),
        .I3(\stat_reg[0]_0 ),
        .I4(abus_0[1]),
        .O(\iv[1]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[1]_i_13 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(bbus_0[0]),
        .I3(abus_0[1]),
        .I4(\stat_reg[0] ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[1]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[1]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[1]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[1]),
        .I4(\iv[1]_i_6_n_0 ),
        .I5(\iv[1]_i_7_n_0 ),
        .O(\iv[1]_i_2_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[1]_i_30 
       (.I0(\badr[0]_INST_0_i_1 ),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_50 ));
  LUT4 #(
    .INIT(16'h0213)) 
    \iv[1]_i_32 
       (.I0(\sr_reg[8]_13 ),
        .I1(\sr_reg[8]_11 ),
        .I2(\iv[1]_i_21_0 ),
        .I3(\iv[1]_i_21_1 ),
        .O(\sr_reg[8]_39 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[1]_i_33 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[1]_i_21 ),
        .O(\iv[10]_i_34 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[1]_i_34 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[0]),
        .O(\badr[0]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[1]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[3]_i_2_1 [1]),
        .I2(\tr[30]_i_2_0 [1]),
        .I3(div_crdy_reg),
        .I4(Q[1]),
        .I5(div_crdy_reg_0),
        .O(\iv[1]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[1]_i_7 
       (.I0(\sr[4]_i_24_2 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_1 ),
        .I2(\iv[1]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[1]_i_13_n_0 ),
        .O(\iv[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[2]_i_1 
       (.I0(\iv[2]_i_2_n_0 ),
        .I1(\tr_reg[2]_0 ),
        .I2(\tr_reg[2]_1 ),
        .I3(\tr_reg[2]_2 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[2]),
        .O(cbus[2]));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[2]_i_12 
       (.I0(abus_0[10]),
        .I1(bbus_0[1]),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_0 ),
        .I4(abus_0[2]),
        .O(\iv[2]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[2]_i_13 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(bbus_0[1]),
        .I3(abus_0[2]),
        .I4(\stat_reg[0] ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[2]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[2]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[2]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[2]),
        .I4(\iv[2]_i_6_n_0 ),
        .I5(\iv[2]_i_7_n_0 ),
        .O(\iv[2]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[2]_i_30 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[1]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_66 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[2]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[3]_i_2_1 [2]),
        .I2(\tr[30]_i_2_0 [2]),
        .I3(div_crdy_reg),
        .I4(Q[2]),
        .I5(div_crdy_reg_0),
        .O(\iv[2]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[2]_i_7 
       (.I0(\sr[4]_i_24_1 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_1 ),
        .I2(\iv[2]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[2]_i_13_n_0 ),
        .O(\iv[2]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[3]_i_1 
       (.I0(\iv[3]_i_2_n_0 ),
        .I1(\iv[3]_i_3_n_0 ),
        .I2(\tr_reg[3]_2 ),
        .I3(\tr_reg[3]_3 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[3]),
        .O(cbus[3]));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[3]_i_13 
       (.I0(abus_0[11]),
        .I1(bbus_0[2]),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_0 ),
        .I4(abus_0[3]),
        .O(\iv[3]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[3]_i_14 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(bbus_0[2]),
        .I3(abus_0[3]),
        .I4(\stat_reg[0] ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[3]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \iv[3]_i_15 
       (.I0(\sr_reg[8]_14 ),
        .I1(\sr_reg[8]_10 ),
        .I2(\sr_reg[8]_7 ),
        .I3(abus_0[31]),
        .I4(\iv[6]_i_8_0 ),
        .I5(\iv[3]_i_8_0 ),
        .O(\iv[3]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[3]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[3]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[3]),
        .I4(\iv[3]_i_6_n_0 ),
        .I5(\iv[3]_i_7_n_0 ),
        .O(\iv[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[3]_i_20 
       (.I0(\sr[4]_i_46 ),
        .I1(\sr_reg[8]_11 ),
        .I2(\sr[4]_i_98 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\iv[3]_i_37_n_0 ),
        .I5(bbus_0[3]),
        .O(\bdatw[12]_INST_0_i_1_2 ));
  LUT6 #(
    .INIT(64'h00000030FFFFFFDD)) 
    \iv[3]_i_22 
       (.I0(\stat_reg[0] ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_0 ),
        .I3(acmd),
        .I4(\stat_reg[0]_2 ),
        .I5(\sr_reg[13] [6]),
        .O(\sr_reg[6]_1 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \iv[3]_i_27 
       (.I0(\sr[4]_i_91_0 ),
        .I1(\sr_reg[8]_13 ),
        .I2(\sr_reg[8]_19 ),
        .O(\sr_reg[8]_14 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[3]_i_3 
       (.I0(\stat_reg[2]_2 ),
        .I1(\iv[3]_i_16 ),
        .I2(\tr_reg[3]_0 ),
        .I3(\tr_reg[3]_1 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[3]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[3]_i_35 
       (.I0(\badr[2]_INST_0_i_1 ),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_49 ));
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \iv[3]_i_37 
       (.I0(\iv[6]_i_8_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\sr_reg[8]_11 ),
        .I3(\sr_reg[8]_13 ),
        .I4(\sr[4]_i_91_0 ),
        .O(\iv[3]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \iv[3]_i_38 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[11]_i_7_2 ),
        .I2(\sr_reg[8]_18 ),
        .I3(\iv[11]_i_7_0 ),
        .O(\sr_reg[8]_41 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[3]_i_39 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[3]_i_21 ),
        .O(\iv[12]_i_34 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[3]_i_40 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[2]),
        .O(\badr[2]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[3]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[3]_i_2_1 [3]),
        .I2(\tr[30]_i_2_0 [3]),
        .I3(div_crdy_reg),
        .I4(Q[3]),
        .I5(div_crdy_reg_0),
        .O(\iv[3]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[3]_i_7 
       (.I0(\iv[3]_i_2_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_1 ),
        .I2(\iv[3]_i_13_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[3]_i_14_n_0 ),
        .O(\iv[3]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[3]_i_8 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I1(\iv[3]_i_15_n_0 ),
        .I2(\sr[4]_i_21 ),
        .O(\iv[3]_i_16 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[4]_i_1 
       (.I0(\iv[4]_i_2_n_0 ),
        .I1(\iv[4]_i_3_n_0 ),
        .I2(\tr_reg[4]_1 ),
        .I3(\tr_reg[4]_0 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[4]),
        .O(cbus[4]));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[4]_i_12 
       (.I0(abus_0[12]),
        .I1(bbus_0[3]),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_0 ),
        .I4(abus_0[4]),
        .O(\iv[4]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF88006A008800)) 
    \iv[4]_i_13 
       (.I0(\stat_reg[0]_0 ),
        .I1(abus_0[4]),
        .I2(\stat_reg[0] ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(bbus_0[3]),
        .I5(\iv[7]_i_34_n_0 ),
        .O(\iv[4]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'h00400040004080C0)) 
    \iv[4]_i_15 
       (.I0(\sr_reg[8]_13 ),
        .I1(\sr_reg[8]_10 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\iv[4]_i_8 ),
        .I4(bbus_0[0]),
        .I5(\iv[4]_i_8_0 ),
        .O(\sr_reg[8]_70 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[4]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[4]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[4]),
        .I4(\iv[4]_i_6_n_0 ),
        .I5(\iv[4]_i_7_n_0 ),
        .O(\iv[4]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[4]_i_3 
       (.I0(\stat_reg[2]_2 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I2(\tr_reg[4]_2 ),
        .I3(\tr_reg[4]_3 ),
        .I4(\tr_reg[4]_4 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[4]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[4]_i_33 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[3]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_65 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[4]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[7]_i_2_0 [0]),
        .I2(\tr[30]_i_2_0 [4]),
        .I3(div_crdy_reg),
        .I4(Q[4]),
        .I5(div_crdy_reg_0),
        .O(\iv[4]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[4]_i_7 
       (.I0(\sr[4]_i_24_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_1 ),
        .I2(\iv[4]_i_12_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[4]_i_13_n_0 ),
        .O(\iv[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[5]_i_1 
       (.I0(\iv[5]_i_2_n_0 ),
        .I1(\iv[5]_i_3_n_0 ),
        .I2(\tr_reg[5]_3 ),
        .I3(\tr_reg[5]_4 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[5]),
        .O(cbus[5]));
  LUT6 #(
    .INIT(64'hFFFF88006A008800)) 
    \iv[5]_i_13 
       (.I0(\stat_reg[0]_0 ),
        .I1(abus_0[5]),
        .I2(\stat_reg[0] ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\bdatw[5] [1]),
        .I5(\iv[7]_i_34_n_0 ),
        .O(\iv[5]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'h004080C0)) 
    \iv[5]_i_16 
       (.I0(\sr_reg[8]_18 ),
        .I1(\sr_reg[8]_10 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\iv[5]_i_8 ),
        .I4(\iv[5]_i_8_0 ),
        .O(\sr_reg[8]_71 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[5]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[5]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[5]),
        .I4(\iv[5]_i_6_n_0 ),
        .I5(\iv[5]_i_7_n_0 ),
        .O(\iv[5]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[5]_i_20 
       (.I0(\iv[13]_i_6_0 ),
        .I1(\sr_reg[8]_19 ),
        .I2(\sr[4]_i_81 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\sr_reg[8]_34 ),
        .I5(bbus_0[3]),
        .O(\bdatw[12]_INST_0_i_1_1 ));
  LUT6 #(
    .INIT(64'hFFFFFEFFFDFFFCFF)) 
    \iv[5]_i_27 
       (.I0(\sr_reg[8]_13 ),
        .I1(\iv[6]_i_8_0 ),
        .I2(\stat_reg[0]_2 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\iv[5]_i_8 ),
        .I5(\iv[5]_i_8_0 ),
        .O(\sr_reg[8]_34 ));
  LUT6 #(
    .INIT(64'hAA08AAAA08080808)) 
    \iv[5]_i_3 
       (.I0(\stat_reg[2]_2 ),
        .I1(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I2(\tr_reg[5]_0 ),
        .I3(\tr_reg[5]_1 ),
        .I4(\tr_reg[5]_2 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[5]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[5]_i_32 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[4]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_64 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[5]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[7]_i_2_0 [1]),
        .I2(Q[5]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [5]),
        .I5(div_crdy_reg),
        .O(\iv[5]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[5]_i_7 
       (.I0(\sr[4]_i_7_1 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_1 ),
        .I2(\sr[4]_i_7_2 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[5]_i_13_n_0 ),
        .O(\iv[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[6]_i_1 
       (.I0(\iv[6]_i_2_n_0 ),
        .I1(\iv[6]_i_3_n_0 ),
        .I2(\tr_reg[6]_1 ),
        .I3(\tr_reg[6]_2 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[6]),
        .O(cbus[6]));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \iv[6]_i_10 
       (.I0(\iv[6]_i_20_n_0 ),
        .I1(\iv[6]_i_21_n_0 ),
        .I2(\iv[6]_i_3_0 ),
        .I3(\iv[6]_i_3_1 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\iv[6]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[6]_i_12 
       (.I0(\stat_reg[0] ),
        .I1(\stat_reg[0]_0 ),
        .I2(\stat_reg[0]_1 ),
        .O(\niho_dsp_a[32]_INST_0_i_5_1 ));
  LUT5 #(
    .INIT(32'h353F3530)) 
    \iv[6]_i_13 
       (.I0(abus_0[14]),
        .I1(bbus_0[4]),
        .I2(\stat_reg[0]_1 ),
        .I3(\stat_reg[0]_0 ),
        .I4(abus_0[6]),
        .O(\iv[6]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[6]_i_14 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(bbus_0[4]),
        .I3(abus_0[6]),
        .I4(\stat_reg[0] ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[6]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[6]_i_15 
       (.I0(\sr_reg[8]_7 ),
        .I1(abus_0[31]),
        .I2(\iv[6]_i_8_0 ),
        .I3(\iv[6]_i_8_1 ),
        .I4(\sr_reg[8]_15 ),
        .I5(\sr_reg[8]_10 ),
        .O(\iv[6]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[6]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[6]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[6]),
        .I4(\iv[6]_i_6_n_0 ),
        .I5(\iv[6]_i_7_n_0 ),
        .O(\iv[6]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \iv[6]_i_20 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[6]_i_10_0 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr[4]_i_78_1 ),
        .O(\iv[6]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[6]_i_21 
       (.I0(\sr_reg[8]_33 ),
        .I1(\sr_reg[8]_15 ),
        .O(\iv[6]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hD8FF)) 
    \iv[6]_i_24 
       (.I0(\sr_reg[8]_13 ),
        .I1(\sr[4]_i_81_0 ),
        .I2(\sr[4]_i_81_1 ),
        .I3(\sr_reg[8]_19 ),
        .O(\sr_reg[8]_15 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[6]_i_3 
       (.I0(\stat_reg[2]_2 ),
        .I1(\iv[6]_i_8_n_0 ),
        .I2(\tr_reg[6]_0 ),
        .I3(\iv[6]_i_10_n_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[6]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[6]_i_31 
       (.I0(\badr[5]_INST_0_i_1 ),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_46 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \iv[6]_i_32 
       (.I0(\sr_reg[8]_19 ),
        .I1(\iv[14]_i_7_1 ),
        .I2(\sr_reg[8]_18 ),
        .I3(\iv[14]_i_7_2 ),
        .O(\sr_reg[6]_4 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[6]_i_33 
       (.I0(\sr_reg[8]_19 ),
        .I1(\iv[6]_i_22 ),
        .O(\iv[15]_i_103 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[6]_i_34 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[5]),
        .O(\badr[5]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[6]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[7]_i_2_0 [2]),
        .I2(Q[6]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [6]),
        .I5(div_crdy_reg),
        .O(\iv[6]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFF4700)) 
    \iv[6]_i_7 
       (.I0(\iv[6]_i_2_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_5_1 ),
        .I2(\iv[6]_i_13_n_0 ),
        .I3(\iv[7]_i_14_n_0 ),
        .I4(\iv[6]_i_14_n_0 ),
        .O(\iv[6]_i_7_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[6]_i_8 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I1(\iv[6]_i_15_n_0 ),
        .I2(\sr[4]_i_18_9 ),
        .O(\iv[6]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \iv[7]_i_1 
       (.I0(\iv[7]_i_2_n_0 ),
        .I1(\iv[7]_i_3_n_0 ),
        .I2(\tr_reg[7]_3 ),
        .I3(\tr_reg[7]_4 ),
        .I4(\stat_reg[0]_3 ),
        .I5(cbus_i[7]),
        .O(cbus[7]));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[7]_i_11 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\badr[6]_INST_0_i_1 ),
        .I3(\iv[6]_i_8_0 ),
        .I4(\iv[7]_i_27_n_0 ),
        .I5(\iv[7]_i_28_n_0 ),
        .O(\iv[7]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[7]_i_14 
       (.I0(\stat_reg[0]_2 ),
        .I1(acmd),
        .O(\iv[7]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hBCE0ECE0A0A0A0A0)) 
    \iv[7]_i_15 
       (.I0(\iv[7]_i_34_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(bbus_0[5]),
        .I3(abus_0[7]),
        .I4(\stat_reg[0] ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\iv[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[7]_i_2 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[7]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[7]),
        .I4(\iv[7]_i_6_n_0 ),
        .I5(\iv[7]_i_7_n_0 ),
        .O(\iv[7]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[7]_i_24 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[6]_i_8_0 ),
        .O(\sr_reg[8]_33 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \iv[7]_i_25 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_91_3 ),
        .I2(\sr_reg[8]_13 ),
        .I3(\iv[7]_i_10_0 ),
        .I4(\sr_reg[8]_19 ),
        .I5(\iv[7]_i_10 ),
        .O(\sr_reg[6]_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[7]_i_26 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[6]),
        .O(\badr[6]_INST_0_i_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[7]_i_27 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[7]_i_11_1 ),
        .O(\iv[7]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDDDDDDFDDDFFF)) 
    \iv[7]_i_28 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[6]_i_8_0 ),
        .I2(\iv[7]_i_11_0 ),
        .I3(\sr_reg[8]_18 ),
        .I4(\iv[11]_i_7_0 ),
        .I5(\sr_reg[8]_11 ),
        .O(\iv[7]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[7]_i_3 
       (.I0(\stat_reg[2]_2 ),
        .I1(\tr_reg[7]_0 ),
        .I2(\tr_reg[7]_1 ),
        .I3(\tr_reg[7]_2 ),
        .I4(\iv[7]_i_11_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[7]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hF0DD)) 
    \iv[7]_i_33 
       (.I0(abus_0[7]),
        .I1(\stat_reg[0]_0 ),
        .I2(bbus_0[5]),
        .I3(\stat_reg[0]_1 ),
        .O(\niho_dsp_a[32]_INST_0_i_5_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \iv[7]_i_34 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .O(\iv[7]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[7]_i_40 
       (.I0(\badr[6]_INST_0_i_1 ),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_52 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[7]_i_6 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[7]_i_2_0 [3]),
        .I2(\tr[30]_i_2_0 [7]),
        .I3(div_crdy_reg),
        .I4(Q[7]),
        .I5(div_crdy_reg_0),
        .O(\iv[7]_i_6_n_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \iv[7]_i_7 
       (.I0(\sr[4]_i_7_0 ),
        .I1(\iv[7]_i_14_n_0 ),
        .I2(\iv[7]_i_15_n_0 ),
        .O(\iv[7]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[8]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[8]),
        .I2(bdatr[0]),
        .I3(\tr_reg[15]_3 ),
        .I4(\iv[8]_i_2_n_0 ),
        .I5(\iv[8]_i_3_n_0 ),
        .O(cbus[8]));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[8]_i_10 
       (.I0(\sr_reg[8]_7 ),
        .I1(abus_0[31]),
        .I2(\iv[6]_i_8_0 ),
        .I3(\iv[8]_i_4_0 ),
        .I4(\sr[7]_i_20_0 ),
        .I5(\sr_reg[8]_10 ),
        .O(\iv[8]_i_10_n_0 ));
  LUT4 #(
    .INIT(16'hF0BB)) 
    \iv[8]_i_15 
       (.I0(\bdatw[8]_INST_0_i_1 ),
        .I1(abus_0[0]),
        .I2(\sr[4]_i_77 ),
        .I3(\sr_reg[8]_19 ),
        .O(\sr[7]_i_20_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[8]_i_17 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[7]),
        .I2(\sr_reg[13] [8]),
        .I3(\iv[14]_i_18_n_0 ),
        .O(\iv[8]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \iv[8]_i_18 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[8]_i_7_1 ),
        .O(\iv[8]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[8]_i_19 
       (.I0(\sr_reg[8]_11 ),
        .I1(\iv[8]_i_7_0 ),
        .O(\iv[8]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[8]_i_2 
       (.I0(\stat_reg[2]_2 ),
        .I1(\iv[8]_i_4_n_0 ),
        .I2(\tr_reg[8]_0 ),
        .I3(\tr_reg[8]_1 ),
        .I4(\iv[8]_i_7_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[8]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hAAFBFBFBBBFBFBFB)) 
    \iv[8]_i_22 
       (.I0(\stat_reg[0]_0 ),
        .I1(abus_0[8]),
        .I2(\stat_reg[2]_1 ),
        .I3(\sr[6]_i_32_n_0 ),
        .I4(bbus_0[6]),
        .I5(\stat_reg[0]_2 ),
        .O(\iv[8]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[8]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[8]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[8]),
        .I4(\iv[8]_i_8_n_0 ),
        .I5(\iv[8]_i_9_n_0 ),
        .O(\iv[8]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \iv[8]_i_33 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[7]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_63 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[8]_i_34 
       (.I0(bbus_0[1]),
        .I1(bbus_0[0]),
        .I2(\bdatw[5] [0]),
        .O(\bdatw[8]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[8]_i_39 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[6]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[8]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[8]_i_39_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[8]_i_4 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I1(\iv[8]_i_10_n_0 ),
        .I2(\iv[8]_i_2_0 ),
        .O(\iv[8]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hF2F22222F2F2F222)) 
    \iv[8]_i_40 
       (.I0(abus_0[0]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(bbus_0[6]),
        .I4(abus_0[8]),
        .I5(\stat_reg[0]_2 ),
        .O(\iv[8]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \iv[8]_i_7 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\iv[8]_i_17_n_0 ),
        .I3(\iv[8]_i_18_n_0 ),
        .I4(\iv[8]_i_19_n_0 ),
        .I5(\sr[4]_i_38 ),
        .O(\iv[8]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[8]_i_8 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[11]_i_3_0 [0]),
        .I2(Q[8]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [8]),
        .I5(div_crdy_reg),
        .O(\iv[8]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h02FFFFFF02FF0000)) 
    \iv[8]_i_9 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\sr[4]_i_8_0 ),
        .I3(\iv[8]_i_22_n_0 ),
        .I4(\stat_reg[0] ),
        .I5(\iv_reg[8]_i_23_n_0 ),
        .O(\iv[8]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \iv[9]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[9]),
        .I2(bdatr[1]),
        .I3(\tr_reg[15]_3 ),
        .I4(\iv[9]_i_2_n_0 ),
        .I5(\iv[9]_i_3_n_0 ),
        .O(cbus[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[9]_i_18 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[8]),
        .O(\iv[9]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h084C)) 
    \iv[9]_i_19 
       (.I0(\sr_reg[8]_18 ),
        .I1(\sr_reg[8]_11 ),
        .I2(\iv[1]_i_21_0 ),
        .I3(\iv[1]_i_21_1 ),
        .O(\iv[9]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8A8AA88888888)) 
    \iv[9]_i_2 
       (.I0(\stat_reg[2]_2 ),
        .I1(\tr_reg[9]_0 ),
        .I2(\tr_reg[9]_1 ),
        .I3(\tr_reg[9]_2 ),
        .I4(\iv[9]_i_7_n_0 ),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\iv[9]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'hDDDF)) 
    \iv[9]_i_20 
       (.I0(\stat_reg[0]_2 ),
        .I1(\iv[6]_i_8_0 ),
        .I2(\iv[9]_i_7_0 ),
        .I3(\sr_reg[8]_11 ),
        .O(\iv[9]_i_20_n_0 ));
  LUT3 #(
    .INIT(8'h20)) 
    \iv[9]_i_21 
       (.I0(\stat_reg[0]_0 ),
        .I1(acmd),
        .I2(\iv[9]_i_42_n_0 ),
        .O(\iv[9]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3F007F7F)) 
    \iv[9]_i_22 
       (.I0(\stat_reg[0]_2 ),
        .I1(bbus_0[7]),
        .I2(\sr[6]_i_32_n_0 ),
        .I3(\stat_reg[2]_1 ),
        .I4(abus_0[9]),
        .O(\iv[9]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hEEAAEEEA)) 
    \iv[9]_i_23 
       (.I0(\tr[25]_i_5_1 ),
        .I1(\sr[6]_i_32_n_0 ),
        .I2(bbus_0[7]),
        .I3(abus_0[9]),
        .I4(\stat_reg[0]_2 ),
        .O(\iv[9]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hB888BBBBB888B888)) 
    \iv[9]_i_24 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(bbus_0[7]),
        .I3(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I4(abus_0[9]),
        .I5(\iv[7]_i_14_n_0 ),
        .O(\iv[9]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF404)) 
    \iv[9]_i_3 
       (.I0(\iv[15]_i_25_n_0 ),
        .I1(mulh[9]),
        .I2(\iv[15]_i_26_n_0 ),
        .I3(niho_dsp_c[9]),
        .I4(\iv[9]_i_8_n_0 ),
        .I5(\iv[9]_i_9_n_0 ),
        .O(\iv[9]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'h4F)) 
    \iv[9]_i_34 
       (.I0(\iv[9]_i_18_n_0 ),
        .I1(\bdatw[12]_INST_0_i_1_0 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_47 ));
  LUT6 #(
    .INIT(64'hAAFF3C00AA003C00)) 
    \iv[9]_i_42 
       (.I0(bbus_0[0]),
        .I1(abus_0[9]),
        .I2(bbus_0[7]),
        .I3(\stat_reg[0]_1 ),
        .I4(\stat_reg[0]_2 ),
        .I5(abus_0[17]),
        .O(\iv[9]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hCECCCECCCECCEEEE)) 
    \iv[9]_i_7 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\iv[9]_i_18_n_0 ),
        .I3(\iv[14]_i_18_n_0 ),
        .I4(\iv[9]_i_19_n_0 ),
        .I5(\iv[9]_i_20_n_0 ),
        .O(\iv[9]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \iv[9]_i_8 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\iv[11]_i_3_0 [1]),
        .I2(\tr[30]_i_2_0 [9]),
        .I3(div_crdy_reg),
        .I4(Q[9]),
        .I5(div_crdy_reg_0),
        .O(\iv[9]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0BFBFAFA0B0B0)) 
    \iv[9]_i_9 
       (.I0(\iv[9]_i_21_n_0 ),
        .I1(\iv[9]_i_22_n_0 ),
        .I2(\stat_reg[0] ),
        .I3(\iv[9]_i_23_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\iv[9]_i_24_n_0 ),
        .O(\iv[9]_i_9_n_0 ));
  MUXF7 \iv_reg[11]_i_22 
       (.I0(\iv[11]_i_39_n_0 ),
        .I1(\iv[11]_i_40_n_0 ),
        .O(\iv_reg[11]_i_22_n_0 ),
        .S(\stat_reg[0]_0 ));
  MUXF7 \iv_reg[14]_i_23 
       (.I0(\iv[14]_i_40_n_0 ),
        .I1(\iv[14]_i_41_n_0 ),
        .O(\iv_reg[14]_i_23_n_0 ),
        .S(\stat_reg[0]_0 ));
  MUXF7 \iv_reg[8]_i_23 
       (.I0(\iv[8]_i_39_n_0 ),
        .I1(\iv[8]_i_40_n_0 ),
        .O(\iv_reg[8]_i_23_n_0 ),
        .S(\stat_reg[0]_0 ));
  LUT3 #(
    .INIT(8'h57)) 
    \mul_a[15]_i_1 
       (.I0(rst_n),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(\sr_reg[13] [8]),
        .O(rst_n_2));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[16]_i_1 
       (.I0(rst_n_fl_reg_14),
        .O(bbus_0[14]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[17]_i_1 
       (.I0(rst_n_fl_reg_13),
        .O(bbus_0[15]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[18]_i_1 
       (.I0(rst_n_fl_reg_12),
        .O(bbus_0[16]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[19]_i_1 
       (.I0(rst_n_fl_reg_11),
        .O(bbus_0[17]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[20]_i_1 
       (.I0(rst_n_fl_reg_10),
        .O(bbus_0[18]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[21]_i_1 
       (.I0(rst_n_fl_reg_9),
        .O(bbus_0[19]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[22]_i_1 
       (.I0(rst_n_fl_reg_8),
        .O(bbus_0[20]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[23]_i_1 
       (.I0(rst_n_fl_reg_7),
        .O(bbus_0[21]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[24]_i_1 
       (.I0(rst_n_fl_reg_6),
        .O(bbus_0[22]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[25]_i_1 
       (.I0(rst_n_fl_reg_16),
        .O(bbus_0[23]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[26]_i_1 
       (.I0(rst_n_fl_reg_5),
        .O(bbus_0[24]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[27]_i_1 
       (.I0(rst_n_fl_reg_4),
        .O(bbus_0[25]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[28]_i_1 
       (.I0(rst_n_fl_reg_3),
        .O(bbus_0[26]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[29]_i_1 
       (.I0(rst_n_fl_reg_2),
        .O(bbus_0[27]));
  LUT1 #(
    .INIT(2'h1)) 
    \mul_b[30]_i_1 
       (.I0(rst_n_fl_reg_1),
        .O(bbus_0[28]));
  LUT3 #(
    .INIT(8'h40)) 
    \mul_b[31]_i_1 
       (.I0(rst_n_fl_reg_0),
        .I1(rst_n),
        .I2(\sr_reg[13] [8]),
        .O(rst_n_0[0]));
  LUT4 #(
    .INIT(16'h4000)) 
    \mul_b[32]_i_1 
       (.I0(rst_n_fl_reg_0),
        .I1(rst_n),
        .I2(\sr_reg[13] [8]),
        .I3(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .O(rst_n_0[1]));
  LUT3 #(
    .INIT(8'h75)) 
    \mulh[15]_i_1 
       (.I0(rst_n),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(\sr_reg[13] [8]),
        .O(rst_n_1));
  LUT2 #(
    .INIT(4'h7)) 
    \mulh[15]_i_2 
       (.I0(rst_n),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .O(mul_b));
  LUT4 #(
    .INIT(16'hFD7F)) 
    \niho_dsp_a[15]_INST_0_i_1 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\stat_reg[0]_0 ),
        .I3(\stat_reg[0]_1 ),
        .O(\niho_dsp_a[32]_INST_0_i_5_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[15]_INST_0_i_2 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[0]_INST_0_i_1_n_0 ),
        .O(\stat_reg[0] ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[15]_INST_0_i_3 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[1]_INST_0_i_1_n_0 ),
        .O(\stat_reg[0]_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \niho_dsp_a[32]_INST_0_i_1 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\stat_reg[0]_1 ),
        .O(\niho_dsp_a[32]_INST_0_i_5_3 ));
  LUT6 #(
    .INIT(64'h0000380000000000)) 
    \niho_dsp_a[32]_INST_0_i_10 
       (.I0(ir[11]),
        .I1(ir[12]),
        .I2(ir[13]),
        .I3(ir[14]),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\niho_dsp_a[32]_INST_0_i_6_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \niho_dsp_a[32]_INST_0_i_11 
       (.I0(\ccmd[0]_INST_0_i_15_n_0 ),
        .I1(ir[6]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[7]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\niho_dsp_a[32]_INST_0_i_17_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h9000900090909000)) 
    \niho_dsp_a[32]_INST_0_i_12 
       (.I0(ir[11]),
        .I1(ir[8]),
        .I2(ir[10]),
        .I3(\niho_dsp_a[32]_INST_0_i_9_0 ),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\niho_dsp_a[32]_INST_0_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h00000008)) 
    \niho_dsp_a[32]_INST_0_i_13 
       (.I0(crdy),
        .I1(div_crdy),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[11]),
        .I4(rst_n_fl_reg_17),
        .O(\niho_dsp_a[32]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFBEAF9E8FFFFFFFF)) 
    \niho_dsp_a[32]_INST_0_i_14 
       (.I0(ir[7]),
        .I1(ir[11]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(ir[8]),
        .I4(\stat[1]_i_10_0 ),
        .I5(\niho_dsp_a[32]_INST_0_i_18_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h0000100000000000)) 
    \niho_dsp_a[32]_INST_0_i_15 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(ir[11]),
        .I2(ir[7]),
        .I3(ir[8]),
        .I4(\stat_reg[2]_12 [0]),
        .I5(ir[10]),
        .O(\niho_dsp_a[32]_INST_0_i_15_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \niho_dsp_a[32]_INST_0_i_17 
       (.I0(ir[4]),
        .I1(ir[5]),
        .I2(ir[3]),
        .O(\niho_dsp_a[32]_INST_0_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niho_dsp_a[32]_INST_0_i_18 
       (.I0(ir[10]),
        .I1(\stat_reg[2]_12 [0]),
        .O(\niho_dsp_a[32]_INST_0_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \niho_dsp_a[32]_INST_0_i_3 
       (.I0(acmd),
        .I1(\stat_reg[0]_2 ),
        .O(\niho_dsp_a[32]_INST_0_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[32]_INST_0_i_4 
       (.I0(\stat_reg[0] ),
        .I1(\stat_reg[0]_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[32]_INST_0_i_5 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[2]_INST_0_i_1_n_0 ),
        .O(\stat_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h00000000FFFF1011)) 
    \niho_dsp_a[32]_INST_0_i_6 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\stat_reg[2]_12 [2]),
        .I2(\niho_dsp_a[32]_INST_0_i_8_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_9_n_0 ),
        .I4(\niho_dsp_a[32]_INST_0_i_10_n_0 ),
        .I5(\stat_reg[0]_3 ),
        .O(acmd));
  LUT2 #(
    .INIT(4'h1)) 
    \niho_dsp_a[32]_INST_0_i_7 
       (.I0(\stat_reg[0]_3 ),
        .I1(\ccmd[3]_INST_0_i_1_n_0 ),
        .O(\stat_reg[0]_2 ));
  LUT6 #(
    .INIT(64'hAAFFFFABAAAAAAAA)) 
    \niho_dsp_a[32]_INST_0_i_8 
       (.I0(\niho_dsp_a[32]_INST_0_i_11_n_0 ),
        .I1(ir[10]),
        .I2(ir[8]),
        .I3(\stat_reg[2]_12 [1]),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\ccmd[4]_INST_0_i_1_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FFFFFF1010)) 
    \niho_dsp_a[32]_INST_0_i_9 
       (.I0(\niho_dsp_a[32]_INST_0_i_12_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_13_n_0 ),
        .I2(\niho_dsp_a[32]_INST_0_i_14_n_0 ),
        .I3(ir[6]),
        .I4(ir[9]),
        .I5(\niho_dsp_a[32]_INST_0_i_15_n_0 ),
        .O(\niho_dsp_a[32]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[10]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[8]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_10_sn_1),
        .O(niho_dsp_b[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[11]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[9]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_11_sn_1),
        .O(niho_dsp_b[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[12]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[10]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_12_sn_1),
        .O(niho_dsp_b[9]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[13]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[11]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_13_sn_1),
        .O(niho_dsp_b[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[14]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[12]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_14_sn_1),
        .O(niho_dsp_b[11]));
  LUT5 #(
    .INIT(32'hC000E222)) 
    \niho_dsp_b[15]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(mul_rslt),
        .I3(niho_dsp_b_15_sn_1),
        .I4(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .O(niho_dsp_b[12]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[16]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_16_sn_1),
        .O(niho_dsp_b[13]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[17]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_17_sn_1),
        .O(niho_dsp_b[14]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[18]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_18_sn_1),
        .O(niho_dsp_b[15]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[19]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_19_sn_1),
        .O(niho_dsp_b[16]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[1]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[0]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_1_sn_1),
        .O(niho_dsp_b[0]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[20]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_20_sn_1),
        .O(niho_dsp_b[17]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[21]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_21_sn_1),
        .O(niho_dsp_b[18]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[22]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_22_sn_1),
        .O(niho_dsp_b[19]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[23]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_23_sn_1),
        .O(niho_dsp_b[20]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[24]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_24_sn_1),
        .O(niho_dsp_b[21]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[25]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_25_sn_1),
        .O(niho_dsp_b[22]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[26]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_26_sn_1),
        .O(niho_dsp_b[23]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[27]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_27_sn_1),
        .O(niho_dsp_b[24]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[28]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_28_sn_1),
        .O(niho_dsp_b[25]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[29]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(niho_dsp_b_29_sn_1),
        .O(niho_dsp_b[26]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[2]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[1]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_2_sn_1),
        .O(niho_dsp_b[1]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[30]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(\niho_dsp_b[30] ),
        .O(niho_dsp_b[27]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[31]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(\niho_dsp_b[32] [0]),
        .O(niho_dsp_b[28]));
  LUT5 #(
    .INIT(32'hEC202020)) 
    \niho_dsp_b[32]_INST_0 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\niho_dsp_a[32]_INST_0_i_5_3 ),
        .I3(mul_rslt),
        .I4(\niho_dsp_b[32] [1]),
        .O(niho_dsp_b[29]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[3]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[2]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_3_sn_1),
        .O(niho_dsp_b[2]));
  LUT2 #(
    .INIT(4'h2)) 
    \niho_dsp_b[4]_INST_0_i_1 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .O(\sr_reg[8]_7 ));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[6]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[4]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_6_sn_1),
        .O(niho_dsp_b[3]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[7]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[5]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_7_sn_1),
        .O(niho_dsp_b[4]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[8]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[6]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_8_sn_1),
        .O(niho_dsp_b[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[9]_INST_0 
       (.I0(\sr_reg[13] [8]),
        .I1(\niho_dsp_a[32]_INST_0_i_5_2 ),
        .I2(bbus_0[7]),
        .I3(mul_rslt),
        .I4(niho_dsp_b_9_sn_1),
        .O(niho_dsp_b[6]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[0]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[0]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[0]),
        .I5(rgf_pc[0]),
        .O(\pc_reg[15] [0]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[10]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[10]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[10]),
        .I5(rgf_pc[10]),
        .O(\pc_reg[15] [10]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[11]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[11]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[11]),
        .I5(rgf_pc[11]),
        .O(\pc_reg[15] [11]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[12]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[12]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[12]),
        .I5(rgf_pc[12]),
        .O(\pc_reg[15] [12]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[13]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[13]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[13]),
        .I5(rgf_pc[13]),
        .O(\pc_reg[15] [13]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[14]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[14]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[14]),
        .I5(rgf_pc[14]),
        .O(\pc_reg[15] [14]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[15]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[15]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[15]),
        .I5(rgf_pc[15]),
        .O(\pc_reg[15] [15]));
  LUT5 #(
    .INIT(32'h00040000)) 
    \pc[15]_i_2 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(\iv[15]_i_6_n_0 ),
        .I4(ctl_selc_rn[0]),
        .O(\rgf/cbus_sel_cr ));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[1]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[1]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[1]),
        .I5(rgf_pc[1]),
        .O(\pc_reg[15] [1]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[2]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[2]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[2]),
        .I5(rgf_pc[2]),
        .O(\pc_reg[15] [2]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[3]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[3]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[3]),
        .I5(rgf_pc[3]),
        .O(\pc_reg[15] [3]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[4]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[4]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[4]),
        .I5(rgf_pc[4]),
        .O(\pc_reg[15] [4]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[5]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[5]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[5]),
        .I5(rgf_pc[5]),
        .O(\pc_reg[15] [5]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[6]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[6]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[6]),
        .I5(rgf_pc[6]),
        .O(\pc_reg[15] [6]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[7]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[7]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[7]),
        .I5(rgf_pc[7]),
        .O(\pc_reg[15] [7]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[8]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[8]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[8]),
        .I5(rgf_pc[8]),
        .O(\pc_reg[15] [8]));
  LUT6 #(
    .INIT(64'hF0FFF011F0EEF000)) 
    \pc[9]_i_1 
       (.I0(ctl_fetch_fl_reg_0),
        .I1(ctl_fetch_ext),
        .I2(cbus[9]),
        .I3(\rgf/cbus_sel_cr ),
        .I4(fch_pc[9]),
        .I5(rgf_pc[9]),
        .O(\pc_reg[15] [9]));
  LUT5 #(
    .INIT(32'hE0FFE000)) 
    \read_cyc[0]_i_1 
       (.I0(\stat_reg[2]_6 ),
        .I1(\stat_reg[0]_6 ),
        .I2(abus_0[0]),
        .I3(brdy),
        .I4(read_cyc[0]),
        .O(brdy_1));
  FDRE rst_n_fl_reg
       (.C(clk),
        .CE(\<const1> ),
        .D(rst_n),
        .Q(rst_n_fl),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[0]_i_1 
       (.I0(cbus[0]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(O),
        .I3(ctl_sp_inc),
        .I4(\sp_reg[0] ),
        .O(\cbus_i[30] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF7FFEFFFF)) 
    \sp[0]_i_10 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[11]),
        .I3(ir[13]),
        .I4(brdy),
        .I5(\sp[0]_i_12_n_0 ),
        .O(\sp[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEFFFFFFEEFFFFFFF)) 
    \sp[0]_i_11 
       (.I0(\sp[0]_i_13_n_0 ),
        .I1(\sp[0]_i_14_n_0 ),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(ir[9]),
        .I5(\sp[0]_i_15_n_0 ),
        .O(\sp[0]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h3FFE)) 
    \sp[0]_i_12 
       (.I0(ir[7]),
        .I1(ir[9]),
        .I2(ir[8]),
        .I3(ir[6]),
        .O(\sp[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAEAFAAA)) 
    \sp[0]_i_13 
       (.I0(\sp[0]_i_16_n_0 ),
        .I1(\bcmd[3]_INST_0_i_16_n_0 ),
        .I2(ir[11]),
        .I3(\stat_reg[2]_12 [1]),
        .I4(brdy),
        .I5(\bcmd[0]_INST_0_i_9_n_0 ),
        .O(\sp[0]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hC4C4CC0C)) 
    \sp[0]_i_14 
       (.I0(brdy),
        .I1(\sp[0]_i_15_n_0 ),
        .I2(\stat_reg[2]_12 [1]),
        .I3(ir[1]),
        .I4(ir[0]),
        .O(\sp[0]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \sp[0]_i_15 
       (.I0(ir[2]),
        .I1(ir[5]),
        .I2(ir[3]),
        .I3(ir[4]),
        .O(\sp[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBFFFFBFE)) 
    \sp[0]_i_16 
       (.I0(ir[7]),
        .I1(ir[12]),
        .I2(ir[10]),
        .I3(ir[11]),
        .I4(ir[9]),
        .I5(\sp[0]_i_13_0 ),
        .O(\sp[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h000000000101FF01)) 
    \sp[0]_i_3 
       (.I0(\sp[0]_i_6_n_0 ),
        .I1(\sp[0]_i_7_n_0 ),
        .I2(\bcmd[0]_INST_0_i_11_n_0 ),
        .I3(\bcmd[0]_INST_0_i_5_n_0 ),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\sp[0]_i_8_n_0 ),
        .O(ctl_sp_inc));
  LUT3 #(
    .INIT(8'hBA)) 
    \sp[0]_i_6 
       (.I0(ir[5]),
        .I1(ir[7]),
        .I2(ir[4]),
        .O(\sp[0]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sp[0]_i_7 
       (.I0(ir[6]),
        .I1(ir[2]),
        .O(\sp[0]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF6FF6FFFF)) 
    \sp[0]_i_8 
       (.I0(ir[11]),
        .I1(ir[12]),
        .I2(ir[14]),
        .I3(ir[13]),
        .I4(\bcmd[0] ),
        .I5(\sp[0]_i_10_n_0 ),
        .O(\sp[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h00000000E8FF3CFF)) 
    \sp[0]_i_9 
       (.I0(brdy),
        .I1(ir[4]),
        .I2(ir[5]),
        .I3(ir[6]),
        .I4(ir[3]),
        .I5(\sp[0]_i_11_n_0 ),
        .O(ctl_sp_id4));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[10]_i_1 
       (.I0(cbus[10]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[10] ),
        .O(\cbus_i[30] [10]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[11]_i_1 
       (.I0(cbus[11]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[11] ),
        .O(\cbus_i[30] [11]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[12]_i_1 
       (.I0(cbus[12]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[12] ),
        .O(\cbus_i[30] [12]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[13]_i_1 
       (.I0(cbus[13]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[13] ),
        .O(\cbus_i[30] [13]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[14]_i_1 
       (.I0(cbus[14]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[14] ),
        .O(\cbus_i[30] [14]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[15]_i_1 
       (.I0(cbus[15]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[15] ),
        .O(\cbus_i[30] [15]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[16]_i_1 
       (.I0(cbus[16]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[16] ),
        .O(\cbus_i[30] [16]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[17]_i_1 
       (.I0(cbus[17]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[17] ),
        .O(\cbus_i[30] [17]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[18]_i_1 
       (.I0(cbus[18]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[18] ),
        .O(\cbus_i[30] [18]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[1]_i_1 
       (.I0(cbus[1]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[1] ),
        .O(\cbus_i[30] [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[20]_i_1 
       (.I0(cbus[19]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[20] ),
        .O(\cbus_i[30] [19]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[22]_i_1 
       (.I0(cbus[20]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[22] ),
        .O(\cbus_i[30] [20]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[24]_i_1 
       (.I0(cbus[21]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[24] ),
        .O(\cbus_i[30] [21]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[25]_i_1 
       (.I0(cbus[22]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[25] ),
        .O(\cbus_i[30] [22]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[26]_i_1 
       (.I0(cbus[23]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[26] ),
        .O(\cbus_i[30] [23]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[2]_i_1 
       (.I0(cbus[2]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[2] ),
        .O(\cbus_i[30] [2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[30]_i_1 
       (.I0(cbus[24]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[30] ),
        .O(\cbus_i[30] [24]));
  LUT5 #(
    .INIT(32'hFFFFFFBD)) 
    \sp[31]_i_10 
       (.I0(ir[0]),
        .I1(ir[3]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(ctl_fetch_ext_fl_i_5_n_0),
        .I4(ir[1]),
        .O(\sp[31]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sp[31]_i_11 
       (.I0(ir[0]),
        .I1(ir[3]),
        .O(\sp[31]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \sp[31]_i_2 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(ctl_selc_rn[0]),
        .I4(ctl_selc_rn[1]),
        .O(\stat_reg[2]_0 [0]));
  LUT6 #(
    .INIT(64'h0000000010061007)) 
    \sp[31]_i_5 
       (.I0(\stat_reg[2]_12 [1]),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[11]),
        .I3(ir[12]),
        .I4(\eir_fl_reg[31]_0 ),
        .I5(\sp[31]_i_6_n_0 ),
        .O(ctl_sp_dec));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4FF)) 
    \sp[31]_i_6 
       (.I0(\sp[31]_i_7_n_0 ),
        .I1(\sp[31]_i_8_n_0 ),
        .I2(\bcmd[0]_INST_0_i_9_n_0 ),
        .I3(brdy),
        .I4(\bcmd[1]_INST_0_i_1_n_0 ),
        .I5(\sp[31]_i_9_n_0 ),
        .O(\sp[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h4042844040408440)) 
    \sp[31]_i_7 
       (.I0(ir[3]),
        .I1(ir[6]),
        .I2(ir[5]),
        .I3(ir[4]),
        .I4(ir[7]),
        .I5(ir[8]),
        .O(\sp[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEAEE)) 
    \sp[31]_i_8 
       (.I0(\sp[31]_i_10_n_0 ),
        .I1(ir[8]),
        .I2(\sp[31]_i_11_n_0 ),
        .I3(\stat_reg[2]_12 [1]),
        .I4(ir[6]),
        .I5(ir[2]),
        .O(\sp[31]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'h77FFFFFE)) 
    \sp[31]_i_9 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(ir[9]),
        .O(\sp[31]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[3]_i_1 
       (.I0(cbus[3]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[3] ),
        .O(\cbus_i[30] [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[4]_i_1 
       (.I0(cbus[4]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[4] ),
        .O(\cbus_i[30] [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[5]_i_1 
       (.I0(cbus[5]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[5] ),
        .O(\cbus_i[30] [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[6]_i_1 
       (.I0(cbus[6]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[6] ),
        .O(\cbus_i[30] [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[7]_i_1 
       (.I0(cbus[7]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[7] ),
        .O(\cbus_i[30] [7]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[8]_i_1 
       (.I0(cbus[8]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[8] ),
        .O(\cbus_i[30] [8]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[9]_i_1 
       (.I0(cbus[9]),
        .I1(\stat_reg[2]_0 [0]),
        .I2(\sp_reg[9] ),
        .O(\cbus_i[30] [9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[0]_i_1 
       (.I0(cbus[0]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr_reg[13] [0]),
        .I3(\stat_reg[2] ),
        .O(\sr_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[10]_i_1 
       (.I0(cbus[10]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr_reg[13] [9]),
        .I3(\stat_reg[2] ),
        .O(\sr_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[11]_i_2 
       (.I0(cbus[11]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr_reg[13] [10]),
        .I3(\stat_reg[2] ),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFEEFFFFFAAA0000)) 
    \sr[12]_i_1 
       (.I0(\sr[12]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr_reg[13] [11]),
        .I3(\sr[13]_i_4_n_0 ),
        .I4(rst_n),
        .I5(cpuid[0]),
        .O(D[0]));
  LUT5 #(
    .INIT(32'h0000FEF0)) 
    \sr[12]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(\sr_reg[13] [11]),
        .I3(cpuid[0]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[12]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFEEFFFFFAAA0000)) 
    \sr[13]_i_1 
       (.I0(\sr[13]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr_reg[13] [12]),
        .I3(\sr[13]_i_4_n_0 ),
        .I4(rst_n),
        .I5(cpuid[1]),
        .O(D[1]));
  LUT5 #(
    .INIT(32'h0000FEF0)) 
    \sr[13]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(\sr_reg[13] [12]),
        .I3(cpuid[1]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[13]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'h0000000400000000)) 
    \sr[13]_i_3 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(ctl_selc_rn[0]),
        .I4(ctl_selc_rn[1]),
        .I5(\sr[7]_i_3_n_0 ),
        .O(\sr[13]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h00004000)) 
    \sr[13]_i_4 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(\iv[15]_i_6_n_0 ),
        .I4(ctl_selc_rn[0]),
        .O(\sr[13]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000000001000000)) 
    \sr[13]_i_5 
       (.I0(\sr[13]_i_6_n_0 ),
        .I1(ir[11]),
        .I2(\stat_reg[2]_12 [1]),
        .I3(\bdatw[9]_INST_0_i_10_n_0 ),
        .I4(\sr[13]_i_7_n_0 ),
        .I5(\sr[13]_i_8_n_0 ),
        .O(ctl_sr_ldie));
  LUT6 #(
    .INIT(64'hFFFFFFFFEFFFFFFF)) 
    \sr[13]_i_6 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[0]),
        .I3(brdy),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\stat_reg[2]_12 [2]),
        .O(\sr[13]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[13]_i_7 
       (.I0(ir[12]),
        .I1(ir[15]),
        .I2(ir[13]),
        .I3(ir[14]),
        .I4(ir[6]),
        .I5(ir[7]),
        .O(\sr[13]_i_7_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[13]_i_8 
       (.I0(ir[1]),
        .I1(ir[9]),
        .I2(ir[10]),
        .I3(ir[8]),
        .O(\sr[13]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFB)) 
    \sr[15]_i_2 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(\iv[15]_i_6_n_0 ),
        .I3(ctl_selc_rn[0]),
        .I4(ctl_selc_rn[1]),
        .O(\stat_reg[2] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[1]_i_1 
       (.I0(cbus[1]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr_reg[13] [1]),
        .I3(\stat_reg[2] ),
        .O(\sr_reg[1] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[2]_i_1 
       (.I0(\sr[2]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(cbus[2]),
        .I3(\sr_reg[13] [2]),
        .I4(\sr[13]_i_4_n_0 ),
        .O(\sr_reg[2] ));
  LUT5 #(
    .INIT(32'h0000FB40)) 
    \sr[2]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(fch_irq_lev[0]),
        .I3(\sr_reg[13] [2]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[2]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \sr[3]_i_1 
       (.I0(\sr[3]_i_2_n_0 ),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(cbus[3]),
        .I3(\sr_reg[13] [3]),
        .I4(\sr[13]_i_4_n_0 ),
        .O(\sr_reg[3] ));
  LUT5 #(
    .INIT(32'h0000FB40)) 
    \sr[3]_i_2 
       (.I0(ctl_sr_upd),
        .I1(ctl_sr_ldie),
        .I2(fch_irq_lev[1]),
        .I3(\sr_reg[13] [3]),
        .I4(\sr[7]_i_3_n_0 ),
        .O(\sr[3]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFEAEAEEEA)) 
    \sr[4]_i_1 
       (.I0(\sr[4]_i_2_n_0 ),
        .I1(\sr[6]_i_2_n_0 ),
        .I2(\sr[4]_i_3_n_0 ),
        .I3(\sr_reg[4]_1 ),
        .I4(\sr_reg[4]_2 ),
        .I5(\sr[4]_i_6_n_0 ),
        .O(\sr_reg[4] ));
  LUT5 #(
    .INIT(32'h00000010)) 
    \sr[4]_i_10 
       (.I0(\tr[20]_i_5_n_0 ),
        .I1(\tr[21]_i_14_0 ),
        .I2(\tr[23]_i_15_0 ),
        .I3(\tr[22]_i_5_n_0 ),
        .I4(\sr[4]_i_27_n_0 ),
        .O(\sr[4]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_100 
       (.I0(\sr_reg[8]_20 ),
        .I1(bbus_0[3]),
        .I2(\iv[13]_i_5 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\iv[6]_i_8_0 ),
        .I5(\sr[4]_i_45 ),
        .O(\sr_reg[8]_24 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \sr[4]_i_103 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\sr[4]_i_46_0 ),
        .I3(\iv[12]_i_34 ),
        .I4(\sr_reg[8]_41 ),
        .I5(\sr[4]_i_38 ),
        .O(\sr_reg[8]_40 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \sr[4]_i_115 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_85 ),
        .I2(\sr_reg[8]_13 ),
        .I3(\sr[4]_i_85_0 ),
        .I4(\sr_reg[8]_19 ),
        .I5(\sr[4]_i_66_1 ),
        .O(\sr[4]_i_115_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDFFFDF)) 
    \sr[4]_i_117 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\iv[9]_i_7_0 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\sr[4]_i_66_2 ),
        .I5(\sr[4]_i_157_n_0 ),
        .O(\sr[4]_i_117_n_0 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \sr[4]_i_120 
       (.I0(\sr_reg[8]_10 ),
        .I1(\sr[4]_i_69 ),
        .I2(\sr_reg[8]_11 ),
        .I3(\sr[4]_i_66_1 ),
        .O(\iv[9]_i_35 ));
  LUT6 #(
    .INIT(64'h000002A2AAAA02A2)) 
    \sr[4]_i_124 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_74_0 ),
        .I2(\sr_reg[8]_13 ),
        .I3(\sr[4]_i_74_1 ),
        .I4(\sr_reg[8]_19 ),
        .I5(\sr[4]_i_77 ),
        .O(\sr[4]_i_124_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFBFFF0FFFB)) 
    \sr[4]_i_125 
       (.I0(\bdatw[8]_INST_0_i_1 ),
        .I1(abus_0[0]),
        .I2(\iv[6]_i_8_0 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\sr_reg[8]_19 ),
        .I5(\sr[4]_i_77 ),
        .O(\sr_reg[8]_22 ));
  LUT6 #(
    .INIT(64'h00000000DFDDDFFF)) 
    \sr[4]_i_126 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\iv[8]_i_7_0 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\iv[8]_i_7_1 ),
        .I5(\iv[8]_i_17_n_0 ),
        .O(\sr[4]_i_126_n_0 ));
  LUT5 #(
    .INIT(32'h0040F040)) 
    \sr[4]_i_129 
       (.I0(\bdatw[8]_INST_0_i_1 ),
        .I1(abus_0[0]),
        .I2(\sr_reg[8]_10 ),
        .I3(\sr_reg[8]_11 ),
        .I4(\sr[4]_i_77 ),
        .O(\iv[8]_i_35 ));
  LUT4 #(
    .INIT(16'h02A2)) 
    \sr[4]_i_131 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_78_1 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr[4]_i_81 ),
        .O(\sr[4]_i_131_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDFFFDF)) 
    \sr[4]_i_133 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\iv[14]_i_7_0 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\sr[4]_i_78_0 ),
        .I5(\sr[4]_i_161_n_0 ),
        .O(\sr[4]_i_133_n_0 ));
  LUT6 #(
    .INIT(64'h0000084CCCCC084C)) 
    \sr[4]_i_135 
       (.I0(\sr_reg[8]_13 ),
        .I1(\sr_reg[8]_10 ),
        .I2(\sr[4]_i_81_0 ),
        .I3(\sr[4]_i_81_1 ),
        .I4(\sr_reg[8]_19 ),
        .I5(\sr[4]_i_81 ),
        .O(\sr_reg[8]_69 ));
  LUT6 #(
    .INIT(64'h020202A2A2A202A2)) 
    \sr[4]_i_136 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_85_1 ),
        .I2(\sr_reg[8]_11 ),
        .I3(\sr[4]_i_85 ),
        .I4(\sr_reg[8]_13 ),
        .I5(\sr[4]_i_85_0 ),
        .O(\sr_reg[6] ));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[4]_i_144 
       (.I0(\sr_reg[8]_10 ),
        .I1(\sr_reg[8]_11 ),
        .I2(\iv[7]_i_10 ),
        .O(\sr[7]_i_21 ));
  LUT6 #(
    .INIT(64'h0000084CCCCC084C)) 
    \sr[4]_i_146 
       (.I0(\sr_reg[8]_13 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\sr[4]_i_91_3 ),
        .I3(\sr[4]_i_91_0 ),
        .I4(\sr_reg[8]_19 ),
        .I5(\sr[4]_i_91_1 ),
        .O(\sr[4]_i_146_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DDDFFFDF)) 
    \sr[4]_i_148 
       (.I0(\stat_reg[0]_2 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\iv[11]_i_7_1 ),
        .I3(\sr_reg[8]_19 ),
        .I4(\sr[4]_i_91_2 ),
        .I5(\sr[4]_i_166_n_0 ),
        .O(\sr[4]_i_148_n_0 ));
  LUT5 #(
    .INIT(32'h0002AA02)) 
    \sr[4]_i_151 
       (.I0(\sr_reg[8]_10 ),
        .I1(\sr[4]_i_91_0 ),
        .I2(\sr_reg[8]_13 ),
        .I3(\sr_reg[8]_11 ),
        .I4(\sr[4]_i_91_1 ),
        .O(\sr_reg[8]_12 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_157 
       (.I0(\sr_reg[13] [8]),
        .I1(\iv[9]_i_18_n_0 ),
        .I2(\iv[14]_i_18_n_0 ),
        .O(\sr[4]_i_157_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_161 
       (.I0(\sr_reg[13] [8]),
        .I1(\iv[14]_i_17_n_0 ),
        .I2(\iv[14]_i_18_n_0 ),
        .O(\sr[4]_i_161_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_166 
       (.I0(\sr_reg[13] [8]),
        .I1(\iv[11]_i_17_n_0 ),
        .I2(\iv[14]_i_18_n_0 ),
        .O(\sr[4]_i_166_n_0 ));
  LUT6 #(
    .INIT(64'hF7F5F3FFFFFFFFFF)) 
    \sr[4]_i_17 
       (.I0(\sr[4]_i_5 ),
        .I1(\sr[4]_i_5_0 ),
        .I2(\iv[0]_i_3_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I4(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I5(\stat_reg[2]_2 ),
        .O(\iv[15]_i_19_0 ));
  LUT6 #(
    .INIT(64'hDF00FF00FF00FF00)) 
    \sr[4]_i_18 
       (.I0(\sr[4]_i_37_n_0 ),
        .I1(\iv[6]_i_8_n_0 ),
        .I2(\sr[4]_i_5_1 ),
        .I3(\stat_reg[2]_2 ),
        .I4(\sr[4]_i_39_n_0 ),
        .I5(\sr[4]_i_40_n_0 ),
        .O(\sr[4]_i_40_0 ));
  LUT3 #(
    .INIT(8'h10)) 
    \sr[4]_i_2 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\sr_reg[13] [4]),
        .O(\sr[4]_i_2_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[4]_i_22 
       (.I0(cbus_i[4]),
        .I1(\stat_reg[0]_3 ),
        .O(\sr[4]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFE0037)) 
    \sr[4]_i_23 
       (.I0(\stat_reg[0] ),
        .I1(\stat_reg[0]_1 ),
        .I2(\stat_reg[0]_0 ),
        .I3(\stat_reg[0]_2 ),
        .I4(acmd),
        .I5(\iv[3]_i_7_n_0 ),
        .O(\sr[4]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_24 
       (.I0(\iv[1]_i_7_n_0 ),
        .I1(\iv[2]_i_7_n_0 ),
        .I2(\iv[6]_i_7_n_0 ),
        .I3(\iv[4]_i_7_n_0 ),
        .O(\sr[4]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \sr[4]_i_25 
       (.I0(\iv[13]_i_8_n_0 ),
        .I1(\iv[9]_i_9_n_0 ),
        .O(\sr[4]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_26 
       (.I0(\tr[27]_i_14 ),
        .I1(\tr[26]_i_5_n_0 ),
        .I2(\tr[24]_i_5_n_0 ),
        .I3(\tr[25]_i_5_n_0 ),
        .O(\sr[4]_i_26_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_27 
       (.I0(\tr[19]_i_14_0 ),
        .I1(\tr[18]_i_5_n_0 ),
        .I2(\tr[17]_i_5_n_0 ),
        .I3(\tr[16]_i_7_n_0 ),
        .O(\sr[4]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01001111)) 
    \sr[4]_i_3 
       (.I0(\sr[4]_i_7_n_0 ),
        .I1(\sr[4]_i_8_n_0 ),
        .I2(\sr[4]_i_9_n_0 ),
        .I3(\sr[4]_i_10_n_0 ),
        .I4(\sr_reg[13] [8]),
        .I5(\sr_reg[4]_3 ),
        .O(\sr[4]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'h0000F888)) 
    \sr[4]_i_30 
       (.I0(\sr[6]_i_25_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I4(\sr_reg[13] [4]),
        .O(\sr_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_37 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I1(\sr[4]_i_66_n_0 ),
        .I2(\sr[4]_i_18_6 ),
        .I3(\sr[4]_i_18_7 ),
        .I4(\sr[4]_i_18_8 ),
        .I5(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .O(\sr[4]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_39 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I1(\sr[4]_i_74_n_0 ),
        .I2(\sr[4]_i_18_0 ),
        .I3(\sr[4]_i_18_1 ),
        .I4(\sr[4]_i_18_2 ),
        .I5(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .O(\sr[4]_i_39_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_40 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I1(\sr[4]_i_78_n_0 ),
        .I2(\sr[4]_i_18_3 ),
        .I3(\sr[4]_i_18_4 ),
        .I4(\sr[4]_i_18_5 ),
        .I5(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .O(\sr[4]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_43 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I1(\sr[4]_i_91_n_0 ),
        .I2(\sr[4]_i_19 ),
        .I3(\sr[4]_i_19_0 ),
        .I4(\sr[4]_i_19_1 ),
        .I5(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .O(\sr_reg[8]_1 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAA8)) 
    \sr[4]_i_6 
       (.I0(\sr[7]_i_3_n_0 ),
        .I1(\sr[4]_i_22_n_0 ),
        .I2(\tr_reg[4]_0 ),
        .I3(\tr_reg[4]_1 ),
        .I4(\iv[4]_i_3_n_0 ),
        .I5(\iv[4]_i_2_n_0 ),
        .O(\sr[4]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_66 
       (.I0(\sr[4]_i_115_n_0 ),
        .I1(\sr[4]_i_37_0 ),
        .I2(\sr[4]_i_37_1 ),
        .I3(\sr[4]_i_117_n_0 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\sr[4]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_7 
       (.I0(\iv[0]_i_7_n_0 ),
        .I1(\iv[5]_i_7_n_0 ),
        .I2(\iv[7]_i_7_n_0 ),
        .I3(\iv[10]_i_8_n_0 ),
        .I4(\sr[4]_i_23_n_0 ),
        .I5(\sr[4]_i_24_n_0 ),
        .O(\sr[4]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \sr[4]_i_73 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\sr[4]_i_38_0 ),
        .I3(\iv[15]_i_103 ),
        .I4(\sr_reg[6]_4 ),
        .I5(\sr[4]_i_38 ),
        .O(\sr_reg[8]_42 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_74 
       (.I0(\sr[4]_i_124_n_0 ),
        .I1(\sr_reg[8]_22 ),
        .I2(\sr[4]_i_39_0 ),
        .I3(\sr[4]_i_126_n_0 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\sr[4]_i_74_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_78 
       (.I0(\sr[4]_i_131_n_0 ),
        .I1(\sr[4]_i_40_1 ),
        .I2(\sr_reg[8]_23 ),
        .I3(\sr[4]_i_133_n_0 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\sr[4]_i_78_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_8 
       (.I0(\iv[15]_i_28_n_0 ),
        .I1(\iv[11]_i_9_n_0 ),
        .I2(\iv[14]_i_9_n_0 ),
        .I3(\iv[8]_i_9_n_0 ),
        .I4(\iv[12]_i_8_n_0 ),
        .I5(\sr[4]_i_25_n_0 ),
        .O(\sr[4]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0E0E0E0EE)) 
    \sr[4]_i_86 
       (.I0(bbus_0[3]),
        .I1(\sr_reg[13] [8]),
        .I2(\sr[4]_i_41 ),
        .I3(\iv[10]_i_34 ),
        .I4(\sr_reg[8]_39 ),
        .I5(\sr[4]_i_38 ),
        .O(\sr_reg[8]_38 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_9 
       (.I0(\tr[31]_i_44_0 ),
        .I1(\tr[30]_i_6_n_0 ),
        .I2(\tr[29]_i_14_0 ),
        .I3(\tr[28]_i_13_0 ),
        .I4(\sr[4]_i_26_n_0 ),
        .O(\sr[4]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h50FF50FF44FF4444)) 
    \sr[4]_i_91 
       (.I0(\sr[4]_i_146_n_0 ),
        .I1(\sr[4]_i_43_0 ),
        .I2(\sr[4]_i_43_1 ),
        .I3(\sr[4]_i_148_n_0 ),
        .I4(\sr_reg[13] [8]),
        .I5(bbus_0[3]),
        .O(\sr[4]_i_91_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_96 
       (.I0(\sr_reg[8]_21 ),
        .I1(bbus_0[3]),
        .I2(\sr_reg[8]_9 ),
        .I3(\stat_reg[0]_2 ),
        .I4(\iv[6]_i_8_0 ),
        .I5(\sr[4]_i_44 ),
        .O(\sr_reg[8]_25 ));
  LUT6 #(
    .INIT(64'hFFFF0000EEE4EEE4)) 
    \sr[5]_i_1 
       (.I0(ctl_sr_upd),
        .I1(\sr_reg[13] [5]),
        .I2(\sr_reg[5]_0 ),
        .I3(\sr[5]_i_3_n_0 ),
        .I4(cbus[5]),
        .I5(\sr[7]_i_3_n_0 ),
        .O(\sr_reg[5] ));
  LUT6 #(
    .INIT(64'h141414FF14FF1414)) 
    \sr[5]_i_3 
       (.I0(\sr[5]_i_8_n_0 ),
        .I1(\sr_reg[8] ),
        .I2(\tr_reg[16]_0 ),
        .I3(\sr[5]_i_9_n_0 ),
        .I4(\sr_reg[7]_0 ),
        .I5(\sr_reg[5]_1 ),
        .O(\sr[5]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'hD21E)) 
    \sr[5]_i_4 
       (.I0(bbus_0[13]),
        .I1(\sr_reg[13] [8]),
        .I2(\stat_reg[2]_3 ),
        .I3(rst_n_fl_reg_14),
        .O(\sr_reg[8]_53 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4000)) 
    \sr[5]_i_8 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(acmd),
        .I3(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I4(bbus_0[3]),
        .I5(\sr_reg[13] [8]),
        .O(\sr[5]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF4000FFFFFFFF)) 
    \sr[5]_i_9 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(acmd),
        .I3(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I4(\bdatw[5] [1]),
        .I5(\sr_reg[13] [8]),
        .O(\sr[5]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFDCDCDCFF101010)) 
    \sr[6]_i_1 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\sr_reg[13] [6]),
        .I3(\sr[6]_i_2_n_0 ),
        .I4(alu_sr_flag),
        .I5(cbus[6]),
        .O(\sr_reg[6]_5 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_13 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[0]_1 ),
        .O(\niho_dsp_a[32]_INST_0_i_5_4 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_14 
       (.I0(\sr[6]_i_32_n_0 ),
        .I1(\stat_reg[0]_2 ),
        .O(\sr[6]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_2 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .O(\sr[6]_i_2_n_0 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[6]_i_25 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[0] ),
        .I2(\stat_reg[0]_1 ),
        .I3(acmd),
        .O(\sr[6]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h1F)) 
    \sr[6]_i_31 
       (.I0(\niho_dsp_a[32]_INST_0_i_7_0 ),
        .I1(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I2(\stat_reg[2]_2 ),
        .O(\iv[15]_i_19_1 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_32 
       (.I0(\stat_reg[0]_1 ),
        .I1(acmd),
        .O(\sr[6]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000FFFDFFFDFFFD)) 
    \sr[6]_i_5 
       (.I0(\niho_dsp_a[32]_INST_0_i_5_4 ),
        .I1(acmd),
        .I2(\stat_reg[0]_2 ),
        .I3(\stat_reg[0] ),
        .I4(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\stat_reg[2]_3 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[6]_i_8 
       (.I0(\stat_reg[2]_3 ),
        .I1(\sr[6]_i_25_n_0 ),
        .O(\sr[6]_i_25_0 ));
  LUT5 #(
    .INIT(32'hFFDCFF10)) 
    \sr[7]_i_1 
       (.I0(ctl_sr_upd),
        .I1(\sr[7]_i_3_n_0 ),
        .I2(\sr_reg[13] [7]),
        .I3(\sr[7]_i_4_n_0 ),
        .I4(cbus[7]),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFF01FF01FFFFFF01)) 
    \sr[7]_i_12 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[24]_i_7 ),
        .I3(\sr[7]_i_23_n_0 ),
        .I4(\sr[7]_i_7 ),
        .I5(\sr[7]_i_7_0 ),
        .O(\sr_reg[8]_16 ));
  LUT2 #(
    .INIT(4'h1)) 
    \sr[7]_i_14 
       (.I0(bbus_0[3]),
        .I1(\iv[15]_i_22 ),
        .O(\sr_reg[8]_10 ));
  LUT6 #(
    .INIT(64'h0000000000000089)) 
    \sr[7]_i_15 
       (.I0(ir[11]),
        .I1(ir[9]),
        .I2(ctl_fetch_fl_reg_2),
        .I3(\ccmd[0]_INST_0_i_22_n_0 ),
        .I4(\sr[7]_i_31_n_0 ),
        .I5(\sr[7]_i_32_n_0 ),
        .O(\sr[7]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \sr[7]_i_16 
       (.I0(bbus_0[2]),
        .I1(\bdatw[5] [0]),
        .I2(bbus_0[0]),
        .I3(bbus_0[1]),
        .I4(\bdatw[5] [1]),
        .I5(bbus_0[3]),
        .O(\bdatw[12]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'h0002000200020000)) 
    \sr[7]_i_2 
       (.I0(\sr[7]_i_5_n_0 ),
        .I1(\stat_reg[2]_12 [2]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(\stat_reg[2]_12 [1]),
        .I4(ir[14]),
        .I5(ir[15]),
        .O(ctl_sr_upd));
  LUT6 #(
    .INIT(64'h5656565656565655)) 
    \sr[7]_i_20 
       (.I0(bbus_0[2]),
        .I1(\iv[0]_i_21 ),
        .I2(\iv[0]_i_21_0 ),
        .I3(bbus_0[1]),
        .I4(bbus_0[0]),
        .I5(\bdatw[5] [0]),
        .O(\sr_reg[8]_19 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFBB77FB77)) 
    \sr[7]_i_23 
       (.I0(\stat_reg[0]_0 ),
        .I1(\stat_reg[2]_2 ),
        .I2(\iv[15]_i_22 ),
        .I3(\stat_reg[0] ),
        .I4(abus_0[31]),
        .I5(\sr[7]_i_44_n_0 ),
        .O(\sr[7]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h565656AAAA56AAAA)) 
    \sr[7]_i_29 
       (.I0(bbus_0[1]),
        .I1(\bdatw[5] [0]),
        .I2(bbus_0[0]),
        .I3(\sr_reg[13] [8]),
        .I4(bbus_0[3]),
        .I5(\bdatw[5] [1]),
        .O(\sr_reg[8]_13 ));
  LUT5 #(
    .INIT(32'h00004004)) 
    \sr[7]_i_3 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(\iv[15]_i_6_n_0 ),
        .I4(ctl_selc_rn[0]),
        .O(\sr[7]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'h8880080888888888)) 
    \sr[7]_i_31 
       (.I0(ir[5]),
        .I1(ir[9]),
        .I2(ir[7]),
        .I3(ir[3]),
        .I4(ir[6]),
        .I5(ir[4]),
        .O(\sr[7]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h00000FFF0BFA0FFF)) 
    \sr[7]_i_32 
       (.I0(ir[4]),
        .I1(ir[3]),
        .I2(ir[7]),
        .I3(ir[6]),
        .I4(ir[9]),
        .I5(ir[5]),
        .O(\sr[7]_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hA8AAA888)) 
    \sr[7]_i_4 
       (.I0(\sr[6]_i_2_n_0 ),
        .I1(\sr[7]_i_6_n_0 ),
        .I2(\sr_reg[7]_0 ),
        .I3(\sr_reg[13] [8]),
        .I4(\sr_reg[8] ),
        .O(\sr[7]_i_4_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[7]_i_44 
       (.I0(\stat_reg[0]_2 ),
        .I1(\stat_reg[0] ),
        .I2(\sr_reg[13] [8]),
        .O(\sr[7]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h2CC02C002CCC2CCC)) 
    \sr[7]_i_5 
       (.I0(\sr[7]_i_8_n_0 ),
        .I1(ir[15]),
        .I2(ir[12]),
        .I3(ir[13]),
        .I4(ir[11]),
        .I5(ir[14]),
        .O(\sr[7]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h000000002E222222)) 
    \sr[7]_i_53 
       (.I0(ir[4]),
        .I1(ctl_selb_0),
        .I2(ir[3]),
        .I3(ir[2]),
        .I4(\bcmd[3]_INST_0_i_13_n_0 ),
        .I5(\bdatw[12]_INST_0_i_4_n_0 ),
        .O(rst_n_fl_reg_19));
  LUT6 #(
    .INIT(64'hCFCFAFAACCCCAFAA)) 
    \sr[7]_i_6 
       (.I0(\iv[15]_i_28_n_0 ),
        .I1(\tr[31]_i_44_0 ),
        .I2(\sr[6]_i_25_0 ),
        .I3(\iv[15]_i_9_0 [3]),
        .I4(\sr_reg[13] [8]),
        .I5(\sr[7]_i_4_0 ),
        .O(\sr[7]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0444044C)) 
    \sr[7]_i_8 
       (.I0(ir[10]),
        .I1(ir[11]),
        .I2(ir[9]),
        .I3(ir[8]),
        .I4(ir[7]),
        .I5(\sr[7]_i_15_n_0 ),
        .O(\sr[7]_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \sr[8]_i_1 
       (.I0(cbus[8]),
        .I1(\sr[13]_i_3_n_0 ),
        .I2(\sr_reg[13] [8]),
        .I3(\stat_reg[2] ),
        .O(\sr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'h0D010D010D010101)) 
    \stat[0]_i_1 
       (.I0(\stat[0]_i_2_n_0 ),
        .I1(ir[12]),
        .I2(ir[15]),
        .I3(\stat_reg[0]_10 ),
        .I4(\stat[0]_i_4_n_0 ),
        .I5(\stat[0]_i_5_n_0 ),
        .O(\stat_reg[2]_5 [0]));
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \stat[0]_i_10 
       (.I0(ir[6]),
        .I1(ir[2]),
        .I2(\bcmd[0]_INST_0_i_12_n_0 ),
        .I3(ir[7]),
        .I4(ir[8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\stat[0]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF4FFF4FFFFFFF4FF)) 
    \stat[0]_i_11 
       (.I0(\stat[0]_i_20_n_0 ),
        .I1(\stat[0]_i_21_n_0 ),
        .I2(ctl_fetch_fl_reg_2),
        .I3(\stat_reg[2]_12 [0]),
        .I4(ir[10]),
        .I5(\stat[0]_i_22_n_0 ),
        .O(\stat[0]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \stat[0]_i_12 
       (.I0(ir[13]),
        .I1(ir[14]),
        .O(\stat[0]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hABAAABABABABABAB)) 
    \stat[0]_i_13 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(\stat[0]_i_24_n_0 ),
        .I2(\stat[0]_i_25_n_0 ),
        .I3(\stat[0]_i_26_n_0 ),
        .I4(brdy),
        .I5(ir[3]),
        .O(\stat[0]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF33F70000)) 
    \stat[0]_i_14 
       (.I0(ir[7]),
        .I1(ir[9]),
        .I2(ir[6]),
        .I3(ir[8]),
        .I4(\ccmd[4]_INST_0_i_1_n_0 ),
        .I5(\stat[0]_i_27_n_0 ),
        .O(\stat[0]_i_14_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_15 
       (.I0(ir[11]),
        .I1(ir[10]),
        .O(\stat[0]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FF0AFFF3)) 
    \stat[0]_i_16 
       (.I0(\stat[1]_i_10_0 ),
        .I1(\sr_reg[13] [8]),
        .I2(ir[9]),
        .I3(ir[8]),
        .I4(ir[7]),
        .I5(\stat[0]_i_28_n_0 ),
        .O(\stat[0]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF0000FF20)) 
    \stat[0]_i_18 
       (.I0(\eir_fl_reg[31]_0 ),
        .I1(ir[3]),
        .I2(\stat[0]_i_29_n_0 ),
        .I3(\stat[0]_i_30_n_0 ),
        .I4(ir[11]),
        .I5(\stat[0]_i_31_n_0 ),
        .O(\stat[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hEEEEEEE0EEEEEEEE)) 
    \stat[0]_i_2 
       (.I0(\stat[0]_i_6_n_0 ),
        .I1(\stat_reg[2]_12 [1]),
        .I2(\stat[0]_i_7_n_0 ),
        .I3(\stat[0]_i_8_n_0 ),
        .I4(\stat[0]_i_9_n_0 ),
        .I5(\stat[0]_i_10_n_0 ),
        .O(\stat[0]_i_2_n_0 ));
  LUT6 #(
    .INIT(64'hEFAAEFAAEFAAAFAA)) 
    \stat[0]_i_20 
       (.I0(\stat[0]_i_23_n_0 ),
        .I1(ir[6]),
        .I2(ir[10]),
        .I3(brdy),
        .I4(\stat[0]_i_32_n_0 ),
        .I5(ir[7]),
        .O(\stat[0]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h9999159111111111)) 
    \stat[0]_i_21 
       (.I0(ir[6]),
        .I1(ir[10]),
        .I2(ir[4]),
        .I3(ir[7]),
        .I4(ir[5]),
        .I5(ir[3]),
        .O(\stat[0]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FFFF7D4D)) 
    \stat[0]_i_22 
       (.I0(\stat[1]_i_10_0 ),
        .I1(ir[8]),
        .I2(ir[11]),
        .I3(brdy),
        .I4(\tr[31]_i_29_n_0 ),
        .I5(\stat[0]_i_33_n_0 ),
        .O(\stat[0]_i_22_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \stat[0]_i_23 
       (.I0(ir[8]),
        .I1(ir[9]),
        .I2(ir[11]),
        .O(\stat[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \stat[0]_i_24 
       (.I0(ir[6]),
        .I1(ir[10]),
        .I2(ir[4]),
        .I3(ir[5]),
        .I4(ir[7]),
        .I5(ir[3]),
        .O(\stat[0]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'h0000510050505050)) 
    \stat[0]_i_25 
       (.I0(ir[6]),
        .I1(ir[3]),
        .I2(brdy),
        .I3(ctl_fetch_inferred_i_44_n_0),
        .I4(ir[4]),
        .I5(ir[10]),
        .O(\stat[0]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'h7777FF7F)) 
    \stat[0]_i_26 
       (.I0(ir[6]),
        .I1(ir[10]),
        .I2(ir[4]),
        .I3(ir[7]),
        .I4(ir[5]),
        .O(\stat[0]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hBBAABAAABBAAAAAA)) 
    \stat[0]_i_27 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\stat[0]_i_34_n_0 ),
        .I2(ir[8]),
        .I3(ir[11]),
        .I4(ir[7]),
        .I5(\sr_reg[13] [8]),
        .O(\stat[0]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'h08)) 
    \stat[0]_i_28 
       (.I0(brdy),
        .I1(ir[9]),
        .I2(ir[6]),
        .O(\stat[0]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h0007)) 
    \stat[0]_i_29 
       (.I0(ir[0]),
        .I1(\stat_reg[2]_12 [0]),
        .I2(\stat_reg[2]_12 [2]),
        .I3(ir[1]),
        .O(\stat[0]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hBAFBBAABFFFFFFFF)) 
    \stat[0]_i_30 
       (.I0(\stat[0]_i_35_n_0 ),
        .I1(ir[0]),
        .I2(ir[1]),
        .I3(ir[3]),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\stat[0]_i_10_n_0 ),
        .O(\stat[0]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFFF8CC88FFFFFFFF)) 
    \stat[0]_i_31 
       (.I0(\stat[0]_i_29_n_0 ),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[3]),
        .I3(ir[11]),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\stat[1]_i_14_n_0 ),
        .O(\stat[0]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h7)) 
    \stat[0]_i_32 
       (.I0(ir[4]),
        .I1(ir[5]),
        .O(\stat[0]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h0000000004440000)) 
    \stat[0]_i_33 
       (.I0(ir[11]),
        .I1(rst_n_fl_reg_17),
        .I2(ir[6]),
        .I3(\bcmd[1]_INST_0_i_5_n_0 ),
        .I4(ir[9]),
        .I5(brdy),
        .O(\stat[0]_i_33_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFDDDDDDDDDDDD)) 
    \stat[0]_i_34 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(crdy),
        .I3(div_crdy),
        .I4(ir[7]),
        .I5(ir[8]),
        .O(\stat[0]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h0000000055F5F575)) 
    \stat[0]_i_35 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(\mul_a_reg[15] [0]),
        .I2(ir[0]),
        .I3(ir[1]),
        .I4(ir[3]),
        .I5(\stat[0]_i_36_n_0 ),
        .O(\stat[0]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'h0DFFFF0D)) 
    \stat[0]_i_36 
       (.I0(ir[0]),
        .I1(\stat_reg[2]_12 [2]),
        .I2(ir[1]),
        .I3(brdy),
        .I4(\stat_reg[2]_12 [0]),
        .O(\stat[0]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'h8808880888088888)) 
    \stat[0]_i_4 
       (.I0(\stat[0]_i_11_n_0 ),
        .I1(\stat[0]_i_12_n_0 ),
        .I2(\stat[0]_i_13_n_0 ),
        .I3(\stat[0]_i_14_n_0 ),
        .I4(\stat[0]_i_15_n_0 ),
        .I5(\stat[0]_i_16_n_0 ),
        .O(\stat[0]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'h0000111130031111)) 
    \stat[0]_i_5 
       (.I0(\stat_reg[0]_11 ),
        .I1(\stat_reg[2]_12 [0]),
        .I2(\sr_reg[13] [7]),
        .I3(ir[11]),
        .I4(ir[13]),
        .I5(ir[14]),
        .O(\stat[0]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hAAA8AAA8AAA8A2A0)) 
    \stat[0]_i_6 
       (.I0(\stat[0]_i_18_n_0 ),
        .I1(ir[11]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(\stat[0]_i_2_0 ),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\stat[1]_i_13_n_0 ),
        .O(\stat[0]_i_6_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \stat[0]_i_7 
       (.I0(ir[14]),
        .I1(\stat_reg[2]_12 [2]),
        .O(\stat[0]_i_7_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[0]_i_8 
       (.I0(ir[3]),
        .I1(ir[0]),
        .O(\stat[0]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFFF)) 
    \stat[0]_i_9 
       (.I0(brdy),
        .I1(ir[1]),
        .I2(ir[13]),
        .I3(ir[11]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\stat[0]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hABAAABAAABAAAAAA)) 
    \stat[1]_i_1 
       (.I0(\stat[1]_i_2_n_0 ),
        .I1(\stat[1]_i_3_n_0 ),
        .I2(\bcmd[1]_INST_0_i_1_n_0 ),
        .I3(ir[12]),
        .I4(\stat_reg[1]_0 ),
        .I5(ir[13]),
        .O(\stat_reg[2]_5 [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4555)) 
    \stat[1]_i_10 
       (.I0(\stat[1]_i_17_n_0 ),
        .I1(\stat[1]_i_18_n_0 ),
        .I2(ir[7]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\stat[1]_i_19_n_0 ),
        .I5(\stat_reg[2]_12 [1]),
        .O(\stat[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF01010100)) 
    \stat[1]_i_11 
       (.I0(\stat[1]_i_20_n_0 ),
        .I1(\bcmd[3]_INST_0_i_16_n_0 ),
        .I2(\stat_reg[2]_12 [1]),
        .I3(\bcmd[0]_INST_0_i_3_n_0 ),
        .I4(\stat[1]_i_21_n_0 ),
        .I5(\stat[1]_i_22_n_0 ),
        .O(\stat[1]_i_11_n_0 ));
  LUT4 #(
    .INIT(16'hB0BB)) 
    \stat[1]_i_13 
       (.I0(ir[13]),
        .I1(\sr_reg[13] [5]),
        .I2(ir[14]),
        .I3(\sr_reg[13] [6]),
        .O(\stat[1]_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_14 
       (.I0(ir[13]),
        .I1(ir[14]),
        .O(\stat[1]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h004400F000440000)) 
    \stat[1]_i_15 
       (.I0(\sr_reg[13] [6]),
        .I1(\stat[1]_i_6_0 ),
        .I2(ctl_fetch_inferred_i_13_n_0),
        .I3(ir[11]),
        .I4(ir[13]),
        .I5(\iv_reg[0] ),
        .O(\stat[1]_i_15_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \stat[1]_i_16 
       (.I0(ir[4]),
        .I1(ir[5]),
        .I2(ir[6]),
        .O(\stat[1]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h2300000000000023)) 
    \stat[1]_i_17 
       (.I0(\stat_reg[2]_12 [0]),
        .I1(ir[7]),
        .I2(\sr_reg[13] [8]),
        .I3(ir[8]),
        .I4(ir[11]),
        .I5(\sr_reg[13] [10]),
        .O(\stat[1]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hF0FFDDFFFFFFDDF0)) 
    \stat[1]_i_18 
       (.I0(brdy),
        .I1(ir[6]),
        .I2(\stat[1]_i_10_0 ),
        .I3(ir[11]),
        .I4(ir[8]),
        .I5(\sr_reg[13] [9]),
        .O(\stat[1]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \stat[1]_i_19 
       (.I0(ir[9]),
        .I1(ir[10]),
        .O(\stat[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h88888888A8AA8888)) 
    \stat[1]_i_2 
       (.I0(\stat[1]_i_5_n_0 ),
        .I1(\stat[1]_i_6_n_0 ),
        .I2(\stat[1]_i_7_n_0 ),
        .I3(\stat[1]_i_8_n_0 ),
        .I4(\stat[1]_i_9_n_0 ),
        .I5(\ccmd[3]_INST_0_i_11_n_0 ),
        .O(\stat[1]_i_2_n_0 ));
  LUT5 #(
    .INIT(32'hC3FFF3DD)) 
    \stat[1]_i_20 
       (.I0(brdy),
        .I1(ir[6]),
        .I2(ir[7]),
        .I3(ir[11]),
        .I4(ir[8]),
        .O(\stat[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h0008800200020000)) 
    \stat[1]_i_21 
       (.I0(ir[8]),
        .I1(ir[3]),
        .I2(ir[4]),
        .I3(ir[5]),
        .I4(ir[7]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\stat[1]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFB000B000B000)) 
    \stat[1]_i_22 
       (.I0(\stat[1]_i_23_n_0 ),
        .I1(ir[11]),
        .I2(\iv_reg[0]_0 ),
        .I3(\stat[1]_i_24_n_0 ),
        .I4(\ccmd[3]_INST_0_i_24_n_0 ),
        .I5(\stat[1]_i_25_n_0 ),
        .O(\stat[1]_i_22_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000100000)) 
    \stat[1]_i_23 
       (.I0(ir[8]),
        .I1(brdy),
        .I2(ir[10]),
        .I3(ir[9]),
        .I4(ir[7]),
        .I5(ir[6]),
        .O(\stat[1]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hCFCCEEEECCCCEEEE)) 
    \stat[1]_i_24 
       (.I0(\stat[1]_i_10_0 ),
        .I1(ir[11]),
        .I2(\iv[15]_i_78_n_0 ),
        .I3(\stat[1]_i_26_n_0 ),
        .I4(rst_n_fl_reg_17),
        .I5(ir[7]),
        .O(\stat[1]_i_24_n_0 ));
  LUT4 #(
    .INIT(16'h0010)) 
    \stat[1]_i_25 
       (.I0(ir[6]),
        .I1(\stat_reg[2]_12 [0]),
        .I2(ir[7]),
        .I3(\stat_reg[2]_12 [1]),
        .O(\stat[1]_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h02)) 
    \stat[1]_i_26 
       (.I0(ir[10]),
        .I1(brdy),
        .I2(ir[8]),
        .O(\stat[1]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'h20F020F020F02000)) 
    \stat[1]_i_3 
       (.I0(\stat[1]_i_10_n_0 ),
        .I1(\stat[1]_i_11_n_0 ),
        .I2(ir[13]),
        .I3(ir[14]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\stat_reg[1]_1 ),
        .O(\stat[1]_i_3_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[1]_i_5 
       (.I0(ir[12]),
        .I1(ir[15]),
        .O(\stat[1]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF000D0000)) 
    \stat[1]_i_6 
       (.I0(\stat[1]_i_13_n_0 ),
        .I1(\stat[1]_i_14_n_0 ),
        .I2(\stat_reg[2]_12 [2]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\ccmd[3]_INST_0_i_19_n_0 ),
        .I5(\stat[1]_i_15_n_0 ),
        .O(\stat[1]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h080002022A200800)) 
    \stat[1]_i_7 
       (.I0(\iv_reg[0]_1 ),
        .I1(ir[1]),
        .I2(\stat_reg[2]_12 [2]),
        .I3(brdy),
        .I4(ir[0]),
        .I5(ir[3]),
        .O(\stat[1]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFAFFFAFFFFFFEFFF)) 
    \stat[1]_i_8 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(brdy),
        .I2(ir[3]),
        .I3(\iv_reg[0]_0 ),
        .I4(ir[1]),
        .I5(ir[0]),
        .O(\stat[1]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \stat[1]_i_9 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(ir[9]),
        .I3(ir[8]),
        .I4(ir[7]),
        .I5(\stat[1]_i_16_n_0 ),
        .O(\stat[1]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'h0101010101010155)) 
    \stat[2]_i_1 
       (.I0(ir[15]),
        .I1(ir[11]),
        .I2(\stat_reg[2]_14 ),
        .I3(\stat[2]_i_3_n_0 ),
        .I4(\stat_reg[2]_12 [2]),
        .I5(\stat_reg[2]_12 [1]),
        .O(\stat_reg[2]_5 [2]));
  LUT6 #(
    .INIT(64'hFFFFFFDFDFDFDFDF)) 
    \stat[2]_i_11 
       (.I0(\bcmd[3]_INST_0_i_2_n_0 ),
        .I1(\tr[31]_i_74_n_0 ),
        .I2(\bcmd[1]_INST_0_i_16_n_0 ),
        .I3(\stat_reg[2]_12 [2]),
        .I4(\stat[0]_i_8_n_0 ),
        .I5(\stat_reg[2]_12 [1]),
        .O(\stat[2]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hA8A8FFFFA8A8FFF0)) 
    \stat[2]_i_3 
       (.I0(\stat[2]_i_6_n_0 ),
        .I1(\stat_reg[2]_13 ),
        .I2(\stat_reg[2]_12 [0]),
        .I3(ir[13]),
        .I4(ir[11]),
        .I5(\mul_b_reg[15]_1 ),
        .O(\stat[2]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hDFFFFFFFFFFFFFFF)) 
    \stat[2]_i_6 
       (.I0(ir[10]),
        .I1(\ccmd[4]_INST_0_i_2_n_0 ),
        .I2(ir[14]),
        .I3(ir[13]),
        .I4(ir[12]),
        .I5(\stat[2]_i_9_n_0 ),
        .O(\stat[2]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF7A327A7A)) 
    \stat[2]_i_8 
       (.I0(\stat[0]_i_8_n_0 ),
        .I1(brdy),
        .I2(ir[1]),
        .I3(\stat_reg[2]_12 [0]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\stat[2]_i_11_n_0 ),
        .O(brdy_0));
  LUT6 #(
    .INIT(64'h0810000000000010)) 
    \stat[2]_i_9 
       (.I0(ir[5]),
        .I1(ir[4]),
        .I2(ir[7]),
        .I3(ir[6]),
        .I4(ir[3]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\stat[2]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF88F8)) 
    \tr[16]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[16]),
        .I2(bdatr[8]),
        .I3(\tr_reg[15]_3 ),
        .I4(\tr_reg[16]_0 ),
        .I5(\tr[16]_i_3_n_0 ),
        .O(cbus[16]));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[16]_i_18 
       (.I0(\tr[16]_i_7_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[16]),
        .I4(rst_n_fl_reg_14),
        .I5(\stat_reg[0] ),
        .O(\tr[16]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[16]_i_19 
       (.I0(rst_n_fl_reg_14),
        .I1(abus_0[16]),
        .I2(\tr[16]_i_7_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[16]_i_19_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[16]_i_21 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(rst_n_fl_reg_14),
        .I2(abus_0[16]),
        .O(\tr[16]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[16]_i_22 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[16]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[16]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hEEFE)) 
    \tr[16]_i_3 
       (.I0(\tr[16]_i_7_n_0 ),
        .I1(\tr[16]_i_8_n_0 ),
        .I2(niho_dsp_c[16]),
        .I3(\tr_reg[30]_1 ),
        .O(\tr[16]_i_3_n_0 ));
  LUT4 #(
    .INIT(16'h70FF)) 
    \tr[16]_i_30 
       (.I0(\stat_reg[0]_2 ),
        .I1(abus_0[15]),
        .I2(\bdatw[12]_INST_0_i_1_0 ),
        .I3(\sr_reg[13] [8]),
        .O(\sr_reg[8]_54 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF444F4F4)) 
    \tr[16]_i_7 
       (.I0(\tr[16]_i_18_n_0 ),
        .I1(\tr[16]_i_19_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I3(\tr[24]_i_5_0 ),
        .I4(\tr[16]_i_21_n_0 ),
        .I5(\tr[16]_i_22_n_0 ),
        .O(\tr[16]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[16]_i_8 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[16]_i_3_0 ),
        .I2(\tr[30]_i_2_0 [16]),
        .I3(div_crdy_reg),
        .I4(Q[16]),
        .I5(div_crdy_reg_0),
        .O(\tr[16]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[17]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[17]),
        .I2(bdatr[9]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[17]),
        .O(cbus[17]));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[17]_i_11 
       (.I0(\tr[17]_i_5_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(rst_n_fl_reg_13),
        .I3(abus_0[17]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\stat_reg[0] ),
        .O(\tr[17]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4C0C)) 
    \tr[17]_i_12 
       (.I0(rst_n_fl_reg_13),
        .I1(abus_0[17]),
        .I2(\stat_reg[2]_1 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[17]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[17]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[17]),
        .I2(rst_n_fl_reg_13),
        .O(\tr[17]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[17]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[17]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[17]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[17]_i_2 
       (.I0(\tr_reg[17]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[17]),
        .I3(\tr[17]_i_4_n_0 ),
        .I4(\tr[17]_i_5_n_0 ),
        .O(p_2_in[17]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[17]_i_4 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[17]_i_2_0 ),
        .I2(Q[17]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [17]),
        .I5(div_crdy_reg),
        .O(\tr[17]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4F4F444)) 
    \tr[17]_i_5 
       (.I0(\tr[17]_i_11_n_0 ),
        .I1(\tr[17]_i_12_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I3(\tr[17]_i_13_n_0 ),
        .I4(\tr[25]_i_5_0 ),
        .I5(\tr[17]_i_15_n_0 ),
        .O(\tr[17]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEBAAAAAAAAA)) 
    \tr[17]_i_8 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr_reg[8]_11 ),
        .I2(\tr[17]_i_3 ),
        .I3(\tr[17]_i_3_0 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(\sr_reg[8]_27 ),
        .O(\sr_reg[8]_31 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[18]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[18]),
        .I2(bdatr[10]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[18]),
        .O(cbus[18]));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[18]_i_11 
       (.I0(\tr[18]_i_5_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(rst_n_fl_reg_12),
        .I3(abus_0[18]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\stat_reg[0] ),
        .O(\tr[18]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[18]_i_12 
       (.I0(rst_n_fl_reg_12),
        .I1(abus_0[18]),
        .I2(\tr[18]_i_5_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[18]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[18]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[18]),
        .I2(rst_n_fl_reg_12),
        .O(\tr[18]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[18]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[18]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[18]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[18]_i_2 
       (.I0(\tr_reg[18]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[18]),
        .I3(\tr[18]_i_4_n_0 ),
        .I4(\tr[18]_i_5_n_0 ),
        .O(p_2_in[18]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[18]_i_4 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[18]_i_2_1 ),
        .I2(Q[18]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [18]),
        .I5(div_crdy_reg),
        .O(\tr[18]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF4F4F444)) 
    \tr[18]_i_5 
       (.I0(\tr[18]_i_11_n_0 ),
        .I1(\tr[18]_i_12_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I3(\tr[18]_i_13_n_0 ),
        .I4(\tr[18]_i_2_0 ),
        .I5(\tr[18]_i_15_n_0 ),
        .O(\tr[18]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h0000014555555555)) 
    \tr[18]_i_6 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr_reg[8]_11 ),
        .I2(\tr[18]_i_3 ),
        .I3(\tr[18]_i_3_0 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(\sr_reg[8]_27 ),
        .O(\sr_reg[8]_28 ));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[19]_i_10 
       (.I0(\tr[19]_i_5_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[19]),
        .I4(rst_n_fl_reg_11),
        .I5(\stat_reg[0] ),
        .O(\tr[19]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[19]_i_11 
       (.I0(rst_n_fl_reg_11),
        .I1(abus_0[19]),
        .I2(\tr[19]_i_5_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[19]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[19]_i_12 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[19]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[19]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[19]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(rst_n_fl_reg_11),
        .I2(abus_0[19]),
        .O(\tr[19]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4F4F4FFF4FFF4)) 
    \tr[19]_i_5 
       (.I0(\tr[19]_i_10_n_0 ),
        .I1(\tr[19]_i_11_n_0 ),
        .I2(\tr[19]_i_12_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I4(\tr[27]_i_5_0 ),
        .I5(\tr[19]_i_14_n_0 ),
        .O(\tr[19]_i_14_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEBAAAAAAAAA)) 
    \tr[19]_i_8 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr_reg[8]_11 ),
        .I2(\tr[19]_i_3 ),
        .I3(\tr[19]_i_3_0 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(\sr_reg[8]_27 ),
        .O(\sr_reg[8]_26 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[20]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[19]),
        .I2(bdatr[11]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[20]),
        .O(cbus[19]));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[20]_i_11 
       (.I0(\tr[20]_i_5_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[20]),
        .I4(rst_n_fl_reg_10),
        .I5(\stat_reg[0] ),
        .O(\tr[20]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[20]_i_12 
       (.I0(rst_n_fl_reg_10),
        .I1(abus_0[20]),
        .I2(\tr[20]_i_5_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[20]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[20]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(rst_n_fl_reg_10),
        .I2(abus_0[20]),
        .O(\tr[20]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[20]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[20]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[20]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hA8A8AA88)) 
    \tr[20]_i_17 
       (.I0(\sr_reg[8]_27 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\tr[20]_i_7 ),
        .I3(\iv[12]_i_26_n_0 ),
        .I4(\sr_reg[8]_19 ),
        .O(\sr_reg[8]_29 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[20]_i_2 
       (.I0(\tr_reg[20]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[19]),
        .I3(\tr[20]_i_4_n_0 ),
        .I4(\tr[20]_i_5_n_0 ),
        .O(p_2_in[20]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[20]_i_4 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[20]_i_2_0 ),
        .I2(\tr[30]_i_2_0 [19]),
        .I3(div_crdy_reg),
        .I4(Q[19]),
        .I5(div_crdy_reg_0),
        .O(\tr[20]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF444F4F4)) 
    \tr[20]_i_5 
       (.I0(\tr[20]_i_11_n_0 ),
        .I1(\tr[20]_i_12_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I3(\sr[4]_i_10_0 ),
        .I4(\tr[20]_i_14_n_0 ),
        .I5(\tr[20]_i_15_n_0 ),
        .O(\tr[20]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'h4544)) 
    \tr[20]_i_6 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr_reg[8]_4 ),
        .I2(\sr[4]_i_66_0 ),
        .I3(\tr[20]_i_3 ),
        .O(\sr_reg[8]_2 ));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[21]_i_10 
       (.I0(\tr[21]_i_5_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[21]),
        .I4(rst_n_fl_reg_9),
        .I5(\stat_reg[0] ),
        .O(\tr[21]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[21]_i_11 
       (.I0(rst_n_fl_reg_9),
        .I1(abus_0[21]),
        .I2(\tr[21]_i_5_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[21]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h5D)) 
    \tr[21]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(rst_n_fl_reg_9),
        .I2(abus_0[21]),
        .O(\tr[21]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[21]_i_14 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[21]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[21]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hA8A8AA88)) 
    \tr[21]_i_16 
       (.I0(\sr_reg[8]_27 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\tr[21]_i_7 ),
        .I3(\iv[13]_i_28_n_0 ),
        .I4(\sr_reg[8]_19 ),
        .O(\sr_reg[8]_30 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF444F4F4)) 
    \tr[21]_i_5 
       (.I0(\tr[21]_i_10_n_0 ),
        .I1(\tr[21]_i_11_n_0 ),
        .I2(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I3(\tr[21]_i_2 ),
        .I4(\tr[21]_i_13_n_0 ),
        .I5(\tr[21]_i_14_n_0 ),
        .O(\tr[21]_i_14_0 ));
  LUT4 #(
    .INIT(16'h4544)) 
    \tr[21]_i_6 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr_reg[8]_4 ),
        .I2(\sr[4]_i_66_0 ),
        .I3(\tr[21]_i_3 ),
        .O(\sr_reg[8]_6 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[22]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[20]),
        .I2(bdatr[12]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[22]),
        .O(cbus[20]));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[22]_i_11 
       (.I0(\tr[22]_i_5_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(rst_n_fl_reg_8),
        .I3(abus_0[22]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\stat_reg[0] ),
        .O(\tr[22]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[22]_i_12 
       (.I0(rst_n_fl_reg_8),
        .I1(abus_0[22]),
        .I2(\tr[22]_i_5_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[22]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[22]_i_13 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[22]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[22]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[22]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[22]),
        .I2(rst_n_fl_reg_8),
        .O(\tr[22]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hA8A8AA88)) 
    \tr[22]_i_16 
       (.I0(\sr_reg[8]_27 ),
        .I1(\sr[4]_i_66_0 ),
        .I2(\tr[22]_i_7_0 ),
        .I3(\iv[14]_i_28_n_0 ),
        .I4(\sr_reg[8]_19 ),
        .O(\tr[22]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[22]_i_2 
       (.I0(\tr_reg[22]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[20]),
        .I3(\tr[22]_i_4_n_0 ),
        .I4(\tr[22]_i_5_n_0 ),
        .O(p_2_in[22]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[22]_i_4 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[22]_i_2_0 ),
        .I2(Q[20]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [20]),
        .I5(div_crdy_reg),
        .O(\tr[22]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFF4FFF4FFF4F4F4)) 
    \tr[22]_i_5 
       (.I0(\tr[22]_i_11_n_0 ),
        .I1(\tr[22]_i_12_n_0 ),
        .I2(\tr[22]_i_13_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I4(\tr[22]_i_14_n_0 ),
        .I5(\sr[4]_i_10_1 ),
        .O(\tr[22]_i_5_n_0 ));
  LUT4 #(
    .INIT(16'hBABB)) 
    \tr[22]_i_7 
       (.I0(\tr[22]_i_16_n_0 ),
        .I1(\sr_reg[8]_4 ),
        .I2(\sr[4]_i_66_0 ),
        .I3(\tr[22]_i_3 ),
        .O(\sr_reg[8]_5 ));
  LUT6 #(
    .INIT(64'h888B8888888B888B)) 
    \tr[23]_i_12 
       (.I0(\tr[23]_i_24_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\tr[23]_i_5_0 ),
        .I3(\tr[25]_i_12_n_0 ),
        .I4(\tr[23]_i_25_n_0 ),
        .I5(\sr[6]_i_14_n_0 ),
        .O(\tr[23]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[23]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[23]),
        .I2(rst_n_fl_reg_7),
        .O(\tr[23]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h3530353F)) 
    \tr[23]_i_15 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\iv[15]_i_111_n_0 ),
        .I2(\stat_reg[0]_1 ),
        .I3(abus_0[23]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[23]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'h0DDDDD0D)) 
    \tr[23]_i_24 
       (.I0(abus_0[15]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[23]),
        .I4(rst_n_fl_reg_7),
        .O(\tr[23]_i_24_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[23]_i_25 
       (.I0(rst_n_fl_reg_7),
        .I1(abus_0[23]),
        .O(\tr[23]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'h888BBBBB888B8888)) 
    \tr[23]_i_5 
       (.I0(\tr[23]_i_12_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[23]_i_2 ),
        .I3(\tr[23]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[23]_i_15_n_0 ),
        .O(\tr[23]_i_15_0 ));
  LUT6 #(
    .INIT(64'hFFFFABFBAAAAAAAA)) 
    \tr[23]_i_8 
       (.I0(\sr_reg[8]_3 ),
        .I1(\tr[23]_i_3_0 ),
        .I2(\sr_reg[8]_11 ),
        .I3(\tr[23]_i_3 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(\sr_reg[8]_27 ),
        .O(\sr_reg[8]_32 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[24]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[21]),
        .I2(bdatr[13]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[24]),
        .O(cbus[21]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[24]_i_12 
       (.I0(\tr[24]_i_17_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\tr[24]_i_18_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[24]_i_5_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[24]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[24]_i_14 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[24]),
        .I2(rst_n_fl_reg_6),
        .O(\tr[24]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[24]_i_15 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[24]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[24]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h1)) 
    \tr[24]_i_16 
       (.I0(\stat_reg[0] ),
        .I1(\tr[24]_i_7 ),
        .O(\sr_reg[8]_27 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[24]_i_17 
       (.I0(abus_0[0]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[24]),
        .I4(rst_n_fl_reg_6),
        .O(\tr[24]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[24]_i_18 
       (.I0(rst_n_fl_reg_6),
        .I1(abus_0[24]),
        .O(\tr[24]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[24]_i_2 
       (.I0(\tr_reg[24]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[21]),
        .I3(\tr[24]_i_4_n_0 ),
        .I4(\tr[24]_i_5_n_0 ),
        .O(p_2_in[24]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[24]_i_4 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[24]_i_2_0 ),
        .I2(\tr[30]_i_2_0 [21]),
        .I3(div_crdy_reg),
        .I4(Q[21]),
        .I5(div_crdy_reg_0),
        .O(\tr[24]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[24]_i_5 
       (.I0(\tr[24]_i_12_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[16]_i_7_0 ),
        .I3(\tr[24]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[24]_i_15_n_0 ),
        .O(\tr[24]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'hEA)) 
    \tr[24]_i_8 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr[7]_i_20_0 ),
        .I2(\tr[24]_i_3 ),
        .O(\sr_reg[8]_36 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[25]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[22]),
        .I2(bdatr[14]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[25]),
        .O(cbus[22]));
  LUT4 #(
    .INIT(16'h0800)) 
    \tr[25]_i_12 
       (.I0(\stat_reg[0]_1 ),
        .I1(\stat_reg[0]_2 ),
        .I2(acmd),
        .I3(bbus_0[13]),
        .O(\tr[25]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'h04444404FFFFFFFF)) 
    \tr[25]_i_13 
       (.I0(\tr[25]_i_5_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[25]),
        .I4(rst_n_fl_reg_16),
        .I5(\stat_reg[0] ),
        .O(\tr[25]_i_13_n_0 ));
  LUT4 #(
    .INIT(16'hF4F0)) 
    \tr[25]_i_14 
       (.I0(rst_n_fl_reg_16),
        .I1(abus_0[25]),
        .I2(\tr[25]_i_5_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .O(\tr[25]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hF2F222F200000000)) 
    \tr[25]_i_15 
       (.I0(abus_0[17]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(rst_n_fl_reg_16),
        .I4(abus_0[25]),
        .I5(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .O(\tr[25]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[25]_i_16 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[25]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[25]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[25]_i_2 
       (.I0(\tr_reg[25]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[22]),
        .I3(\tr[25]_i_4_n_0 ),
        .I4(\tr[25]_i_5_n_0 ),
        .O(p_2_in[25]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[25]_i_4 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[25]_i_2_0 ),
        .I2(\tr[30]_i_2_0 [22]),
        .I3(div_crdy_reg),
        .I4(Q[22]),
        .I5(div_crdy_reg_0),
        .O(\tr[25]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF0F0E)) 
    \tr[25]_i_5 
       (.I0(\stat_reg[0]_0 ),
        .I1(\tr[25]_i_12_n_0 ),
        .I2(\tr[25]_i_13_n_0 ),
        .I3(\tr[25]_i_14_n_0 ),
        .I4(\tr[25]_i_15_n_0 ),
        .I5(\tr[25]_i_16_n_0 ),
        .O(\tr[25]_i_5_n_0 ));
  LUT3 #(
    .INIT(8'h7F)) 
    \tr[25]_i_8 
       (.I0(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I1(\stat_reg[0]_2 ),
        .I2(\sr_reg[13] [8]),
        .O(\sr_reg[8]_37 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[26]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[23]),
        .I2(bdatr[15]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[26]),
        .O(cbus[23]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[26]_i_11 
       (.I0(\tr[26]_i_16_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\tr[26]_i_17_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[18]_i_2_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[26]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[26]_i_12 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[26]),
        .I2(rst_n_fl_reg_5),
        .O(\tr[26]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[26]_i_14 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[26]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[26]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[26]_i_16 
       (.I0(abus_0[2]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[26]),
        .I4(rst_n_fl_reg_5),
        .O(\tr[26]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[26]_i_17 
       (.I0(rst_n_fl_reg_5),
        .I1(abus_0[26]),
        .O(\tr[26]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[26]_i_2 
       (.I0(\tr_reg[26]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[23]),
        .I3(\tr[26]_i_4_n_0 ),
        .I4(\tr[26]_i_5_n_0 ),
        .O(p_2_in[26]));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[26]_i_4 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[26]_i_2_0 ),
        .I2(Q[23]),
        .I3(div_crdy_reg_0),
        .I4(\tr[30]_i_2_0 [23]),
        .I5(div_crdy_reg),
        .O(\tr[26]_i_4_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[26]_i_5 
       (.I0(\tr[26]_i_11_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[26]_i_12_n_0 ),
        .I3(\tr[18]_i_5_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[26]_i_14_n_0 ),
        .O(\tr[26]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h04404444FFFFFFFF)) 
    \tr[27]_i_10 
       (.I0(\tr[27]_i_5_1 ),
        .I1(\stat_reg[0]_0 ),
        .I2(rst_n_fl_reg_4),
        .I3(abus_0[27]),
        .I4(\sr[6]_i_14_n_0 ),
        .I5(\stat_reg[0] ),
        .O(\tr[27]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF4F0)) 
    \tr[27]_i_11 
       (.I0(rst_n_fl_reg_4),
        .I1(abus_0[27]),
        .I2(\tr[27]_i_5_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[27]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hCCCC88C0000088C0)) 
    \tr[27]_i_12 
       (.I0(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I1(\niho_dsp_a[32]_INST_0_i_4_n_0 ),
        .I2(\iv[7]_i_14_n_0 ),
        .I3(abus_0[27]),
        .I4(\stat_reg[0]_1 ),
        .I5(\iv[15]_i_111_n_0 ),
        .O(\tr[27]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[27]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[27]),
        .I2(rst_n_fl_reg_4),
        .O(\tr[27]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFAAA7555)) 
    \tr[27]_i_15 
       (.I0(\stat_reg[0] ),
        .I1(abus_0[31]),
        .I2(\sr_reg[13] [8]),
        .I3(\bdatw[12]_INST_0_i_1_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\stat_reg[0]_2 ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'hFFF4FFF4FFF4F4F4)) 
    \tr[27]_i_5 
       (.I0(\tr[27]_i_10_n_0 ),
        .I1(\tr[27]_i_11_n_0 ),
        .I2(\tr[27]_i_12_n_0 ),
        .I3(\niho_dsp_a[15]_INST_0_i_2_0 ),
        .I4(\tr[27]_i_13_n_0 ),
        .I5(\tr[19]_i_5_0 ),
        .O(\tr[27]_i_14 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[28]_i_10 
       (.I0(\tr[28]_i_15_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\tr[28]_i_16_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\sr[4]_i_10_0 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[28]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[28]_i_12 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[28]),
        .I2(rst_n_fl_reg_3),
        .O(\tr[28]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[28]_i_13 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[28]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[28]_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \tr[28]_i_14 
       (.I0(\tr[28]_i_9_0 ),
        .I1(\sr_reg[8]_13 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(\sr_reg[8]_27 ),
        .O(\tr[28]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[28]_i_15 
       (.I0(abus_0[4]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[28]),
        .I4(rst_n_fl_reg_3),
        .O(\tr[28]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[28]_i_16 
       (.I0(rst_n_fl_reg_3),
        .I1(abus_0[28]),
        .O(\tr[28]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[28]_i_5 
       (.I0(\tr[28]_i_10_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[20]_i_5_0 ),
        .I3(\tr[28]_i_12_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[28]_i_13_n_0 ),
        .O(\tr[28]_i_13_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \tr[28]_i_9 
       (.I0(\sr_reg[8]_9 ),
        .I1(\tr[24]_i_3 ),
        .I2(\tr[28]_i_14_n_0 ),
        .I3(\tr[28]_i_3 ),
        .I4(\sr_reg[8]_10 ),
        .O(\sr_reg[8]_8 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[29]_i_11 
       (.I0(\tr[29]_i_16_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\tr[29]_i_17_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\tr[21]_i_2 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[29]_i_11_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[29]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[29]),
        .I2(rst_n_fl_reg_2),
        .O(\tr[29]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[29]_i_14 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[29]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[29]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \tr[29]_i_15 
       (.I0(\tr[29]_i_7 ),
        .I1(\sr_reg[8]_13 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(\sr_reg[8]_27 ),
        .O(\sr_reg[8]_68 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[29]_i_16 
       (.I0(abus_0[5]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[29]),
        .I4(rst_n_fl_reg_2),
        .O(\tr[29]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[29]_i_17 
       (.I0(rst_n_fl_reg_2),
        .I1(abus_0[29]),
        .O(\tr[29]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[29]_i_5 
       (.I0(\tr[29]_i_11_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[21]_i_5_0 ),
        .I3(\tr[29]_i_13_n_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[29]_i_14_n_0 ),
        .O(\tr[29]_i_14_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[30]_i_1 
       (.I0(\stat_reg[0]_3 ),
        .I1(cbus_i[24]),
        .I2(bdatr[16]),
        .I3(read_cyc[2]),
        .I4(read_cyc[1]),
        .I5(p_2_in[30]),
        .O(cbus[24]));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBB8B88)) 
    \tr[30]_i_12 
       (.I0(\tr[30]_i_19_n_0 ),
        .I1(\stat_reg[0]_0 ),
        .I2(\tr[30]_i_20_n_0 ),
        .I3(\sr[6]_i_14_n_0 ),
        .I4(\sr[4]_i_10_1 ),
        .I5(\tr[25]_i_12_n_0 ),
        .O(\tr[30]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[30]_i_13 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[30]),
        .I2(rst_n_fl_reg_1),
        .O(\tr[30]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[30]_i_15 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[30]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[30]_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hDDFFD0FF50FF50FF)) 
    \tr[30]_i_17 
       (.I0(\sr_reg[8]_7 ),
        .I1(abus_0[31]),
        .I2(\tr[30]_i_21_n_0 ),
        .I3(\stat_reg[0] ),
        .I4(\tr[19]_i_9 ),
        .I5(\sr[4]_i_66_0 ),
        .O(\sr_reg[8]_4 ));
  LUT6 #(
    .INIT(64'hFFFFFFEFFF00FF00)) 
    \tr[30]_i_18 
       (.I0(\tr[30]_i_8 ),
        .I1(\sr_reg[8]_13 ),
        .I2(\sr_reg[8]_19 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\sr[4]_i_66_0 ),
        .I5(\sr_reg[8]_27 ),
        .O(\sr_reg[8]_67 ));
  LUT5 #(
    .INIT(32'hF22222F2)) 
    \tr[30]_i_19 
       (.I0(abus_0[6]),
        .I1(\stat_reg[2]_1 ),
        .I2(\sr[6]_i_14_n_0 ),
        .I3(abus_0[30]),
        .I4(rst_n_fl_reg_1),
        .O(\tr[30]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[30]_i_2 
       (.I0(\tr_reg[30]_0 ),
        .I1(\tr_reg[30]_1 ),
        .I2(niho_dsp_c[24]),
        .I3(\tr[30]_i_5_n_0 ),
        .I4(\tr[30]_i_6_n_0 ),
        .O(p_2_in[30]));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[30]_i_20 
       (.I0(rst_n_fl_reg_1),
        .I1(abus_0[30]),
        .O(\tr[30]_i_20_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[30]_i_21 
       (.I0(\bdatw[12]_INST_0_i_1_0 ),
        .I1(\iv[15]_i_22 ),
        .O(\tr[30]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'h44F444F4FFFF44F4)) 
    \tr[30]_i_5 
       (.I0(\sr[6]_i_25_0 ),
        .I1(\tr[30]_i_2_1 ),
        .I2(\tr[30]_i_2_0 [24]),
        .I3(div_crdy_reg),
        .I4(Q[24]),
        .I5(div_crdy_reg_0),
        .O(\tr[30]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[30]_i_6 
       (.I0(\tr[30]_i_12_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[30]_i_13_n_0 ),
        .I3(\tr[22]_i_5_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[30]_i_15_n_0 ),
        .O(\tr[30]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'h00040000)) 
    \tr[31]_i_1 
       (.I0(ctl_selc[0]),
        .I1(ctl_selc[1]),
        .I2(ctl_selc_rn[1]),
        .I3(ctl_selc_rn[0]),
        .I4(\iv[15]_i_6_n_0 ),
        .O(\stat_reg[2]_0 [2]));
  LUT6 #(
    .INIT(64'hFF00FF10FFFFFF10)) 
    \tr[31]_i_10 
       (.I0(\tr[31]_i_24_n_0 ),
        .I1(\ccmd[4]_INST_0_i_4_n_0 ),
        .I2(\stat_reg[2]_12 [1]),
        .I3(\tr[31]_i_25_n_0 ),
        .I4(\stat_reg[2]_12 [0]),
        .I5(\tr[31]_i_26_n_0 ),
        .O(\tr[31]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hEAEE000000000000)) 
    \tr[31]_i_11 
       (.I0(\tr[31]_i_27_n_0 ),
        .I1(\tr[31]_i_28_n_0 ),
        .I2(\tr[31]_i_29_n_0 ),
        .I3(\stat[1]_i_10_0 ),
        .I4(\iv[15]_i_43_n_0 ),
        .I5(ir[3]),
        .O(\tr[31]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4500)) 
    \tr[31]_i_12 
       (.I0(\tr[31]_i_30_n_0 ),
        .I1(\tr[31]_i_6_n_0 ),
        .I2(ir[8]),
        .I3(\tr[31]_i_31_n_0 ),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\stat_reg[2]_12 [0]),
        .O(\tr[31]_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hBBB8BBBBBBB88888)) 
    \tr[31]_i_15 
       (.I0(\tr[31]_i_41_n_0 ),
        .I1(\stat_reg[0] ),
        .I2(\tr[31]_i_42_n_0 ),
        .I3(\tr[23]_i_5_0 ),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[31]_i_44_n_0 ),
        .O(\tr[31]_i_44_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00003070)) 
    \tr[31]_i_16 
       (.I0(ir[7]),
        .I1(ir[9]),
        .I2(ir[4]),
        .I3(ir[8]),
        .I4(ir[10]),
        .I5(\tr[31]_i_45_n_0 ),
        .O(\tr[31]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h00000000DFFF7F7F)) 
    \tr[31]_i_17 
       (.I0(\ccmd[3]_INST_0_i_23_n_0 ),
        .I1(ir[6]),
        .I2(ir[1]),
        .I3(ir[4]),
        .I4(ir[5]),
        .I5(\tr[31]_i_46_n_0 ),
        .O(\tr[31]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'h0000000080830000)) 
    \tr[31]_i_18 
       (.I0(ir[6]),
        .I1(ir[7]),
        .I2(ir[8]),
        .I3(\sr_reg[13] [8]),
        .I4(ir[4]),
        .I5(\stat[1]_i_19_n_0 ),
        .O(\tr[31]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hBBABAAAABBBBBBBB)) 
    \tr[31]_i_19 
       (.I0(\ccmd[1]_INST_0_i_1_0 ),
        .I1(\tr[31]_i_47_n_0 ),
        .I2(ir[4]),
        .I3(\iv[15]_i_44_n_0 ),
        .I4(\tr[31]_i_48_n_0 ),
        .I5(rst_n_fl_reg_20),
        .O(\tr[31]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hBFAABFFFBFFFBFFF)) 
    \tr[31]_i_20 
       (.I0(\tr[31]_i_49_n_0 ),
        .I1(\iv[15]_i_72_n_0 ),
        .I2(ir[1]),
        .I3(ir[8]),
        .I4(ir[4]),
        .I5(\iv[15]_i_75_n_0 ),
        .O(\tr[31]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h44F4444400000000)) 
    \tr[31]_i_21 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(\ccmd[3]_INST_0_i_10_n_0 ),
        .I2(\iv[15]_i_90_n_0 ),
        .I3(ir[3]),
        .I4(\bcmd[0]_INST_0_i_12_n_0 ),
        .I5(ir[1]),
        .O(\tr[31]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \tr[31]_i_22 
       (.I0(ir[6]),
        .I1(ir[5]),
        .I2(ir[4]),
        .I3(ir[9]),
        .I4(ir[8]),
        .I5(ir[7]),
        .O(\tr[31]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \tr[31]_i_23 
       (.I0(ir[2]),
        .I1(ir[3]),
        .I2(ir[1]),
        .I3(ir[0]),
        .O(\tr[31]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h0707070700070707)) 
    \tr[31]_i_24 
       (.I0(\tr[31]_i_50_n_0 ),
        .I1(\iv[15]_i_72_n_0 ),
        .I2(\tr[31]_i_51_n_0 ),
        .I3(\iv[15]_i_90_n_0 ),
        .I4(\bcmd[0]_INST_0_i_12_n_0 ),
        .I5(\stat[0]_i_8_n_0 ),
        .O(\tr[31]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF001100F1)) 
    \tr[31]_i_25 
       (.I0(\tr[31]_i_52_n_0 ),
        .I1(\ccmd[1]_INST_0_i_1_0 ),
        .I2(\tr[31]_i_53_n_0 ),
        .I3(\ccmd[2]_INST_0_i_8_n_0 ),
        .I4(\tr[31]_i_54_n_0 ),
        .I5(\stat_reg[2]_12 [2]),
        .O(\tr[31]_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    \tr[31]_i_26 
       (.I0(\tr[31]_i_22_n_0 ),
        .I1(\tr[31]_i_23_n_0 ),
        .I2(ir[10]),
        .I3(ir[15]),
        .I4(\stat_reg[2]_12 [1]),
        .I5(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\tr[31]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF00004100)) 
    \tr[31]_i_27 
       (.I0(\iv[15]_i_87_n_0 ),
        .I1(ir[8]),
        .I2(ir[11]),
        .I3(ir[10]),
        .I4(ir[9]),
        .I5(\tr[31]_i_55_n_0 ),
        .O(\tr[31]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hFEAAAAAAAAAAAAAA)) 
    \tr[31]_i_28 
       (.I0(\ccmd[4]_INST_0_i_1_n_0 ),
        .I1(\bcmd[0]_INST_0_i_12_n_0 ),
        .I2(ir[6]),
        .I3(ir[10]),
        .I4(\iv[15]_i_35_n_0 ),
        .I5(\tr[31]_i_56_n_0 ),
        .O(\tr[31]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \tr[31]_i_29 
       (.I0(ir[9]),
        .I1(ir[7]),
        .O(\tr[31]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hF200F200F200FFFF)) 
    \tr[31]_i_3 
       (.I0(ir[9]),
        .I1(\tr[31]_i_6_n_0 ),
        .I2(\tr[31]_i_7_n_0 ),
        .I3(\iv_reg[0] ),
        .I4(\tr[31]_i_8_n_0 ),
        .I5(\stat_reg[2]_12 [2]),
        .O(ctl_selc_rn[1]));
  LUT4 #(
    .INIT(16'h0305)) 
    \tr[31]_i_30 
       (.I0(\tr[31]_i_12_0 ),
        .I1(\tr[31]_i_58_n_0 ),
        .I2(ir[15]),
        .I3(ir[14]),
        .O(\tr[31]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hBABBAAAABABBBABB)) 
    \tr[31]_i_31 
       (.I0(\ccmd[4]_INST_0_i_4_n_0 ),
        .I1(\tr[31]_i_59_n_0 ),
        .I2(\tr[31]_i_60_n_0 ),
        .I3(ir[3]),
        .I4(\tr[31]_i_61_n_0 ),
        .I5(\ccmd[0]_INST_0_i_15_n_0 ),
        .O(\tr[31]_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hDDD0DDDD)) 
    \tr[31]_i_4 
       (.I0(\stat_reg[2]_12 [2]),
        .I1(\tr[31]_i_9_n_0 ),
        .I2(\tr[31]_i_10_n_0 ),
        .I3(\tr[31]_i_11_n_0 ),
        .I4(\tr[31]_i_12_n_0 ),
        .O(ctl_selc_rn[0]));
  LUT6 #(
    .INIT(64'hEAAEFFFFEAAE0000)) 
    \tr[31]_i_41 
       (.I0(\iv[15]_i_28_0 ),
        .I1(\sr[6]_i_14_n_0 ),
        .I2(abus_0[31]),
        .I3(rst_n_fl_reg_0),
        .I4(\stat_reg[0]_0 ),
        .I5(\tr[31]_i_70_n_0 ),
        .O(\tr[31]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \tr[31]_i_42 
       (.I0(\sr[6]_i_14_n_0 ),
        .I1(abus_0[31]),
        .I2(rst_n_fl_reg_0),
        .O(\tr[31]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[31]_i_44 
       (.I0(\iv[15]_i_111_n_0 ),
        .I1(\stat_reg[0]_1 ),
        .I2(\niho_dsp_a[32]_INST_0_i_3_n_0 ),
        .I3(abus_0[31]),
        .I4(\iv[7]_i_14_n_0 ),
        .O(\tr[31]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h00101010FFFFFFFF)) 
    \tr[31]_i_45 
       (.I0(\stat[1]_i_19_n_0 ),
        .I1(ir[7]),
        .I2(ir[4]),
        .I3(\sr_reg[13] [8]),
        .I4(ir[8]),
        .I5(ir[11]),
        .O(\tr[31]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h0000800000800008)) 
    \tr[31]_i_46 
       (.I0(\tr[31]_i_71_n_0 ),
        .I1(ir[1]),
        .I2(ir[6]),
        .I3(ir[5]),
        .I4(ir[3]),
        .I5(ir[4]),
        .O(\tr[31]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h00FF000100010001)) 
    \tr[31]_i_47 
       (.I0(ir[10]),
        .I1(\tr[31]_i_72_n_0 ),
        .I2(brdy),
        .I3(\ccmd[2]_INST_0_i_8_n_0 ),
        .I4(\bcmd[1]_INST_0_i_12_n_0 ),
        .I5(\fch_irq_lev[1]_i_5_n_0 ),
        .O(\tr[31]_i_47_n_0 ));
  LUT5 #(
    .INIT(32'h8AAAAAAA)) 
    \tr[31]_i_48 
       (.I0(\tr[31]_i_73_n_0 ),
        .I1(\iv[15]_i_88_n_0 ),
        .I2(\ccmd[0]_INST_0_i_15_n_0 ),
        .I3(ir[1]),
        .I4(ir[3]),
        .O(\tr[31]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'hB7)) 
    \tr[31]_i_49 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(ir[9]),
        .O(\tr[31]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF000040004000)) 
    \tr[31]_i_50 
       (.I0(ir[6]),
        .I1(brdy),
        .I2(ir[7]),
        .I3(ir[3]),
        .I4(ir[0]),
        .I5(ir[8]),
        .O(\tr[31]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000008F80)) 
    \tr[31]_i_51 
       (.I0(ir[3]),
        .I1(\iv[15]_i_75_n_0 ),
        .I2(ir[9]),
        .I3(ir[0]),
        .I4(\stat[0]_i_15_n_0 ),
        .I5(ir[8]),
        .O(\tr[31]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'hFFFBFFFFFFFFFFFB)) 
    \tr[31]_i_52 
       (.I0(\tr[31]_i_74_n_0 ),
        .I1(brdy),
        .I2(ir[2]),
        .I3(\tr[31]_i_75_n_0 ),
        .I4(ir[3]),
        .I5(ir[0]),
        .O(\tr[31]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \tr[31]_i_53 
       (.I0(ir[15]),
        .I1(\stat_reg[2]_12 [1]),
        .I2(\stat_reg[2]_12 [0]),
        .I3(\tr[31]_i_76_n_0 ),
        .I4(ir[2]),
        .I5(\stat[0]_i_8_n_0 ),
        .O(\tr[31]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \tr[31]_i_54 
       (.I0(ir[6]),
        .I1(ir[5]),
        .I2(ir[4]),
        .I3(ir[7]),
        .I4(ir[8]),
        .I5(\ccmd[1]_INST_0_i_17_n_0 ),
        .O(\tr[31]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0600060000000400)) 
    \tr[31]_i_55 
       (.I0(ir[11]),
        .I1(ir[10]),
        .I2(\iv[15]_i_78_n_0 ),
        .I3(brdy),
        .I4(ir[7]),
        .I5(ir[8]),
        .O(\tr[31]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h80F88080FFF8FF80)) 
    \tr[31]_i_56 
       (.I0(ir[0]),
        .I1(brdy),
        .I2(ir[5]),
        .I3(ir[7]),
        .I4(ir[4]),
        .I5(ir[6]),
        .O(\tr[31]_i_56_n_0 ));
  LUT5 #(
    .INIT(32'hEBBEBEBE)) 
    \tr[31]_i_58 
       (.I0(ir[13]),
        .I1(\sr_reg[13] [5]),
        .I2(ir[11]),
        .I3(ir[12]),
        .I4(\sr_reg[13] [7]),
        .O(\tr[31]_i_58_n_0 ));
  LUT6 #(
    .INIT(64'h0000011100000000)) 
    \tr[31]_i_59 
       (.I0(\ccmd[1]_INST_0_i_11_n_0 ),
        .I1(ir[7]),
        .I2(ir[8]),
        .I3(\sr_reg[13] [8]),
        .I4(ir[9]),
        .I5(ir[3]),
        .O(\tr[31]_i_59_n_0 ));
  LUT5 #(
    .INIT(32'hD5D55D55)) 
    \tr[31]_i_6 
       (.I0(ir[15]),
        .I1(ir[13]),
        .I2(ir[14]),
        .I3(ir[11]),
        .I4(ir[12]),
        .O(\tr[31]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFEEFFFF0F00FF)) 
    \tr[31]_i_60 
       (.I0(ir[8]),
        .I1(ir[7]),
        .I2(\tr[31]_i_77_n_0 ),
        .I3(ir[11]),
        .I4(ir[10]),
        .I5(ir[9]),
        .O(\tr[31]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hF3FFBFFF0EFEDEFF)) 
    \tr[31]_i_61 
       (.I0(ir[3]),
        .I1(ir[4]),
        .I2(ir[6]),
        .I3(ir[0]),
        .I4(ir[7]),
        .I5(ir[5]),
        .O(\tr[31]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h00000000ABABAB00)) 
    \tr[31]_i_7 
       (.I0(\tr[31]_i_16_n_0 ),
        .I1(\bcmd[3]_INST_0_i_16_n_0 ),
        .I2(\tr[31]_i_17_n_0 ),
        .I3(ir[11]),
        .I4(\tr[31]_i_18_n_0 ),
        .I5(\ccmd[4]_INST_0_i_4_n_0 ),
        .O(\tr[31]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hD5DFC0C055550000)) 
    \tr[31]_i_70 
       (.I0(\stat_reg[2]_1 ),
        .I1(bbus_0[13]),
        .I2(\stat_reg[0]_2 ),
        .I3(rst_n_fl_reg_0),
        .I4(abus_0[31]),
        .I5(\sr[6]_i_32_n_0 ),
        .O(\tr[31]_i_70_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[31]_i_71 
       (.I0(ir[8]),
        .I1(ir[7]),
        .O(\tr[31]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF7)) 
    \tr[31]_i_72 
       (.I0(\bcmd[3]_INST_0_i_13_n_0 ),
        .I1(ir[3]),
        .I2(ir[2]),
        .I3(ir[7]),
        .I4(\bdatw[31]_INST_0_i_78_n_0 ),
        .I5(\stat[1]_i_16_n_0 ),
        .O(\tr[31]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFD5FF)) 
    \tr[31]_i_73 
       (.I0(ir[8]),
        .I1(ir[7]),
        .I2(\stat[1]_i_10_0 ),
        .I3(ir[4]),
        .I4(ir[9]),
        .I5(\ccmd[1]_INST_0_i_11_n_0 ),
        .O(\tr[31]_i_73_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \tr[31]_i_74 
       (.I0(ir[10]),
        .I1(ir[9]),
        .I2(ir[8]),
        .I3(ir[7]),
        .O(\tr[31]_i_74_n_0 ));
  LUT4 #(
    .INIT(16'hFFFD)) 
    \tr[31]_i_75 
       (.I0(ir[1]),
        .I1(ir[6]),
        .I2(ir[5]),
        .I3(ir[4]),
        .O(\tr[31]_i_75_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[31]_i_76 
       (.I0(ir[1]),
        .I1(brdy),
        .O(\tr[31]_i_76_n_0 ));
  LUT4 #(
    .INIT(16'hC101)) 
    \tr[31]_i_77 
       (.I0(\sr_reg[13] [8]),
        .I1(ir[8]),
        .I2(ir[7]),
        .I3(ir[6]),
        .O(\tr[31]_i_77_n_0 ));
  LUT6 #(
    .INIT(64'hAAAA0008AAAAAAAA)) 
    \tr[31]_i_8 
       (.I0(\tr[31]_i_19_n_0 ),
        .I1(\tr[31]_i_20_n_0 ),
        .I2(\tr[31]_i_21_n_0 ),
        .I3(\ccmd[4]_INST_0_i_1_n_0 ),
        .I4(\ccmd[4]_INST_0_i_4_n_0 ),
        .I5(\iv_reg[0]_0 ),
        .O(\tr[31]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000040000)) 
    \tr[31]_i_9 
       (.I0(\tr[31]_i_22_n_0 ),
        .I1(\tr[31]_i_23_n_0 ),
        .I2(ir[10]),
        .I3(ir[15]),
        .I4(\iv_reg[0]_1 ),
        .I5(\ccmd[2]_INST_0_i_8_n_0 ),
        .O(\tr[31]_i_9_n_0 ));
endmodule

module niho_fsm
   (\stat_reg[2]_0 ,
    Q,
    \sr_reg[7] ,
    \stat_reg[1]_0 ,
    \stat_reg[0]_0 ,
    \stat_reg[1]_1 ,
    \stat_reg[1]_2 ,
    \stat_reg[0]_1 ,
    \stat_reg[0]_2 ,
    \stat_reg[1]_3 ,
    \stat_reg[0]_3 ,
    \stat_reg[2]_1 ,
    \stat_reg[0]_4 ,
    \stat_reg[1]_4 ,
    \stat_reg[2]_2 ,
    \stat_reg[1]_5 ,
    \stat_reg[1]_6 ,
    \stat_reg[0]_5 ,
    \stat_reg[1]_7 ,
    \stat_reg[1]_8 ,
    \stat_reg[0]_6 ,
    \stat_reg[2]_3 ,
    \stat_reg[1]_9 ,
    \stat_reg[2]_4 ,
    \stat_reg[1]_10 ,
    \stat_reg[1]_11 ,
    out,
    rgf_sr_flag,
    \stat[2]_i_2_0 ,
    ctl_fetch_fl_reg,
    \bcmd[2] ,
    \bcmd[2]_0 ,
    p_0_in,
    D,
    clk);
  output \stat_reg[2]_0 ;
  output [2:0]Q;
  output \sr_reg[7] ;
  output \stat_reg[1]_0 ;
  output \stat_reg[0]_0 ;
  output \stat_reg[1]_1 ;
  output \stat_reg[1]_2 ;
  output \stat_reg[0]_1 ;
  output \stat_reg[0]_2 ;
  output \stat_reg[1]_3 ;
  output \stat_reg[0]_3 ;
  output \stat_reg[2]_1 ;
  output \stat_reg[0]_4 ;
  output \stat_reg[1]_4 ;
  output \stat_reg[2]_2 ;
  output \stat_reg[1]_5 ;
  output \stat_reg[1]_6 ;
  output \stat_reg[0]_5 ;
  output \stat_reg[1]_7 ;
  output \stat_reg[1]_8 ;
  output \stat_reg[0]_6 ;
  output \stat_reg[2]_3 ;
  output \stat_reg[1]_9 ;
  output \stat_reg[2]_4 ;
  output \stat_reg[1]_10 ;
  output \stat_reg[1]_11 ;
  input [8:0]out;
  input [2:0]rgf_sr_flag;
  input \stat[2]_i_2_0 ;
  input ctl_fetch_fl_reg;
  input \bcmd[2] ;
  input \bcmd[2]_0 ;
  input p_0_in;
  input [2:0]D;
  input clk;

  wire \<const1> ;
  wire [2:0]D;
  wire [2:0]Q;
  wire \bcmd[2] ;
  wire \bcmd[2]_0 ;
  wire clk;
  wire ctl_fetch_fl_reg;
  wire [8:0]out;
  wire p_0_in;
  wire [2:0]rgf_sr_flag;
  wire \sr_reg[7] ;
  wire \stat[2]_i_2_0 ;
  wire \stat[2]_i_4_n_0 ;
  wire \stat_reg[0]_0 ;
  wire \stat_reg[0]_1 ;
  wire \stat_reg[0]_2 ;
  wire \stat_reg[0]_3 ;
  wire \stat_reg[0]_4 ;
  wire \stat_reg[0]_5 ;
  wire \stat_reg[0]_6 ;
  wire \stat_reg[1]_0 ;
  wire \stat_reg[1]_1 ;
  wire \stat_reg[1]_10 ;
  wire \stat_reg[1]_11 ;
  wire \stat_reg[1]_2 ;
  wire \stat_reg[1]_3 ;
  wire \stat_reg[1]_4 ;
  wire \stat_reg[1]_5 ;
  wire \stat_reg[1]_6 ;
  wire \stat_reg[1]_7 ;
  wire \stat_reg[1]_8 ;
  wire \stat_reg[1]_9 ;
  wire \stat_reg[2]_0 ;
  wire \stat_reg[2]_1 ;
  wire \stat_reg[2]_2 ;
  wire \stat_reg[2]_3 ;
  wire \stat_reg[2]_4 ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'h01)) 
    \badr[31]_INST_0_i_10 
       (.I0(Q[2]),
        .I1(Q[0]),
        .I2(Q[1]),
        .O(\stat_reg[2]_2 ));
  LUT3 #(
    .INIT(8'h01)) 
    \bcmd[0]_INST_0_i_10 
       (.I0(Q[2]),
        .I1(out[8]),
        .I2(Q[1]),
        .O(\stat_reg[2]_4 ));
  LUT2 #(
    .INIT(4'h2)) 
    \bcmd[1]_INST_0_i_6 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\stat_reg[0]_2 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \bcmd[2]_INST_0_i_1 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(out[8]),
        .I3(Q[2]),
        .I4(\bcmd[2] ),
        .I5(\bcmd[2]_0 ),
        .O(\stat_reg[1]_2 ));
  LUT2 #(
    .INIT(4'h1)) 
    \bcmd[3]_INST_0_i_3 
       (.I0(Q[0]),
        .I1(out[2]),
        .O(\stat_reg[0]_1 ));
  LUT2 #(
    .INIT(4'h6)) 
    \bdatw[31]_INST_0_i_62 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\stat_reg[0]_3 ));
  LUT4 #(
    .INIT(16'h1001)) 
    \ccmd[0]_INST_0_i_14 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(rgf_sr_flag[0]),
        .I3(out[4]),
        .O(\stat_reg[1]_5 ));
  LUT2 #(
    .INIT(4'h1)) 
    \ccmd[0]_INST_0_i_6 
       (.I0(Q[0]),
        .I1(Q[1]),
        .O(\stat_reg[0]_5 ));
  LUT2 #(
    .INIT(4'h2)) 
    \ccmd[1]_INST_0_i_10 
       (.I0(Q[1]),
        .I1(Q[0]),
        .O(\stat_reg[1]_7 ));
  LUT3 #(
    .INIT(8'hEF)) 
    \ccmd[1]_INST_0_i_12 
       (.I0(out[8]),
        .I1(Q[1]),
        .I2(Q[0]),
        .O(\stat_reg[1]_9 ));
  LUT2 #(
    .INIT(4'hE)) 
    \ccmd[2]_INST_0_i_13 
       (.I0(Q[1]),
        .I1(out[3]),
        .O(\stat_reg[1]_8 ));
  LUT3 #(
    .INIT(8'hDF)) 
    \ccmd[2]_INST_0_i_14 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[0]),
        .O(\stat_reg[2]_0 ));
  LUT4 #(
    .INIT(16'h0100)) 
    \ccmd[2]_INST_0_i_3 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(out[8]),
        .O(\stat_reg[1]_10 ));
  LUT6 #(
    .INIT(64'hFFFFFAFAFFFFF8FA)) 
    ctl_fetch_inferred_i_3
       (.I0(Q[0]),
        .I1(\stat_reg[1]_1 ),
        .I2(out[8]),
        .I3(out[7]),
        .I4(Q[2]),
        .I5(ctl_fetch_fl_reg),
        .O(\stat_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hAA8A)) 
    ctl_fetch_inferred_i_50
       (.I0(Q[1]),
        .I1(out[1]),
        .I2(out[0]),
        .I3(Q[2]),
        .O(\stat_reg[1]_3 ));
  LUT2 #(
    .INIT(4'hB)) 
    ctl_fetch_inferred_i_9
       (.I0(Q[1]),
        .I1(out[6]),
        .O(\stat_reg[1]_1 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \eir_fl[31]_i_3 
       (.I0(Q[2]),
        .I1(Q[1]),
        .I2(out[4]),
        .I3(Q[0]),
        .O(\stat_reg[2]_1 ));
  LUT2 #(
    .INIT(4'h1)) 
    \fch_irq_lev[1]_i_6 
       (.I0(Q[0]),
        .I1(out[4]),
        .O(\stat_reg[0]_4 ));
  LUT5 #(
    .INIT(32'h01101001)) 
    \iv[15]_i_119 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(out[4]),
        .I3(rgf_sr_flag[0]),
        .I4(rgf_sr_flag[2]),
        .O(\stat_reg[1]_6 ));
  LUT3 #(
    .INIT(8'h10)) 
    \niho_dsp_a[32]_INST_0_i_16 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(out[8]),
        .O(\stat_reg[1]_11 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sp[0]_i_17 
       (.I0(Q[2]),
        .I1(out[8]),
        .I2(Q[0]),
        .O(\stat_reg[2]_3 ));
  LUT2 #(
    .INIT(4'h1)) 
    \stat[0]_i_3 
       (.I0(Q[1]),
        .I1(Q[2]),
        .O(\stat_reg[1]_4 ));
  LUT3 #(
    .INIT(8'hBE)) 
    \stat[1]_i_12 
       (.I0(Q[0]),
        .I1(rgf_sr_flag[2]),
        .I2(out[4]),
        .O(\stat_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h88A0AAAAAAAAAAAA)) 
    \stat[2]_i_2 
       (.I0(\stat[2]_i_4_n_0 ),
        .I1(rgf_sr_flag[2]),
        .I2(rgf_sr_flag[1]),
        .I3(out[5]),
        .I4(out[6]),
        .I5(\stat_reg[1]_0 ),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFF51055551)) 
    \stat[2]_i_4 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(out[1]),
        .I4(out[0]),
        .I5(\stat[2]_i_2_0 ),
        .O(\stat[2]_i_4_n_0 ));
  LUT4 #(
    .INIT(16'h0001)) 
    \stat[2]_i_5 
       (.I0(Q[1]),
        .I1(Q[0]),
        .I2(Q[2]),
        .I3(out[7]),
        .O(\stat_reg[1]_0 ));
  FDRE \stat_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(Q[0]),
        .R(p_0_in));
  FDRE \stat_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(Q[1]),
        .R(p_0_in));
  FDRE \stat_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[2]),
        .Q(Q[2]),
        .R(p_0_in));
endmodule

module niho_mem
   (D,
    \cbus_i[31] ,
    read_cyc,
    .bdatr_0_sp_1(bdatr_0_sn_1),
    .bdatr_1_sp_1(bdatr_1_sn_1),
    .bdatr_2_sp_1(bdatr_2_sn_1),
    .bdatr_3_sp_1(bdatr_3_sn_1),
    .bdatr_4_sp_1(bdatr_4_sn_1),
    .bdatr_5_sp_1(bdatr_5_sn_1),
    .bdatr_6_sp_1(bdatr_6_sn_1),
    .bdatr_7_sp_1(bdatr_7_sn_1),
    \read_cyc_reg[1] ,
    .bdatr_8_sp_1(bdatr_8_sn_1),
    .bdatr_9_sp_1(bdatr_9_sn_1),
    .bdatr_10_sp_1(bdatr_10_sn_1),
    .bdatr_11_sp_1(bdatr_11_sn_1),
    .bdatr_12_sp_1(bdatr_12_sn_1),
    .bdatr_13_sp_1(bdatr_13_sn_1),
    .bdatr_14_sp_1(bdatr_14_sn_1),
    .bdatr_15_sp_1(bdatr_15_sn_1),
    \sr_reg[8] ,
    \sp_reg[27] ,
    \sp_reg[31] ,
    \sp_reg[23] ,
    \sp_reg[29] ,
    \sp_reg[28] ,
    \sp_reg[21] ,
    \sp_reg[19] ,
    \sp_reg[27]_0 ,
    \tr_reg[27] ,
    cbus_i,
    bdatr,
    p_2_in,
    out,
    \grn_reg[15] ,
    bcmd,
    brdy,
    p_0_in,
    clk,
    \read_cyc_reg[0] );
  output [6:0]D;
  output [6:0]\cbus_i[31] ;
  output [2:0]read_cyc;
  output \read_cyc_reg[1] ;
  output [6:0]\sr_reg[8] ;
  input [0:0]\sp_reg[27] ;
  input \sp_reg[31] ;
  input \sp_reg[23] ;
  input \sp_reg[29] ;
  input \sp_reg[28] ;
  input \sp_reg[21] ;
  input \sp_reg[19] ;
  input \sp_reg[27]_0 ;
  input \tr_reg[27] ;
  input [6:0]cbus_i;
  input [22:0]bdatr;
  input [6:0]p_2_in;
  input [0:0]out;
  input [6:0]\grn_reg[15] ;
  input [1:0]bcmd;
  input brdy;
  input p_0_in;
  input clk;
  input \read_cyc_reg[0] ;
  output bdatr_0_sn_1;
  output bdatr_1_sn_1;
  output bdatr_2_sn_1;
  output bdatr_3_sn_1;
  output bdatr_4_sn_1;
  output bdatr_5_sn_1;
  output bdatr_6_sn_1;
  output bdatr_7_sn_1;
  output bdatr_8_sn_1;
  output bdatr_9_sn_1;
  output bdatr_10_sn_1;
  output bdatr_11_sn_1;
  output bdatr_12_sn_1;
  output bdatr_13_sn_1;
  output bdatr_14_sn_1;
  output bdatr_15_sn_1;

  wire [6:0]D;
  wire [1:0]bcmd;
  wire [22:0]bdatr;
  wire bdatr_0_sn_1;
  wire bdatr_10_sn_1;
  wire bdatr_11_sn_1;
  wire bdatr_12_sn_1;
  wire bdatr_13_sn_1;
  wire bdatr_14_sn_1;
  wire bdatr_15_sn_1;
  wire bdatr_1_sn_1;
  wire bdatr_2_sn_1;
  wire bdatr_3_sn_1;
  wire bdatr_4_sn_1;
  wire bdatr_5_sn_1;
  wire bdatr_6_sn_1;
  wire bdatr_7_sn_1;
  wire bdatr_8_sn_1;
  wire bdatr_9_sn_1;
  wire brdy;
  wire [6:0]cbus_i;
  wire [6:0]\cbus_i[31] ;
  wire clk;
  wire [6:0]\grn_reg[15] ;
  wire [0:0]out;
  wire p_0_in;
  wire [6:0]p_2_in;
  wire [2:0]read_cyc;
  wire \read_cyc_reg[0] ;
  wire \read_cyc_reg[1] ;
  wire \sp_reg[19] ;
  wire \sp_reg[21] ;
  wire \sp_reg[23] ;
  wire [0:0]\sp_reg[27] ;
  wire \sp_reg[27]_0 ;
  wire \sp_reg[28] ;
  wire \sp_reg[29] ;
  wire \sp_reg[31] ;
  wire [6:0]\sr_reg[8] ;
  wire \tr_reg[27] ;

  niho_mem_bctl bctl
       (.D(D),
        .bcmd(bcmd),
        .bdatr(bdatr),
        .bdatr_0_sp_1(bdatr_0_sn_1),
        .bdatr_10_sp_1(bdatr_10_sn_1),
        .bdatr_11_sp_1(bdatr_11_sn_1),
        .bdatr_12_sp_1(bdatr_12_sn_1),
        .bdatr_13_sp_1(bdatr_13_sn_1),
        .bdatr_14_sp_1(bdatr_14_sn_1),
        .bdatr_15_sp_1(bdatr_15_sn_1),
        .bdatr_1_sp_1(bdatr_1_sn_1),
        .bdatr_2_sp_1(bdatr_2_sn_1),
        .bdatr_3_sp_1(bdatr_3_sn_1),
        .bdatr_4_sp_1(bdatr_4_sn_1),
        .bdatr_5_sp_1(bdatr_5_sn_1),
        .bdatr_6_sp_1(bdatr_6_sn_1),
        .bdatr_7_sp_1(bdatr_7_sn_1),
        .bdatr_8_sp_1(bdatr_8_sn_1),
        .bdatr_9_sp_1(bdatr_9_sn_1),
        .brdy(brdy),
        .cbus_i(cbus_i),
        .\cbus_i[31] (\cbus_i[31] ),
        .clk(clk),
        .\grn_reg[15] (\grn_reg[15] ),
        .out(out),
        .p_0_in(p_0_in),
        .p_2_in(p_2_in),
        .\read_cyc_reg[0]_0 (read_cyc[0]),
        .\read_cyc_reg[0]_1 (\read_cyc_reg[0] ),
        .\read_cyc_reg[1]_0 (read_cyc[1]),
        .\read_cyc_reg[1]_1 (\read_cyc_reg[1] ),
        .\read_cyc_reg[2]_0 (read_cyc[2]),
        .\sp_reg[19] (\sp_reg[19] ),
        .\sp_reg[21] (\sp_reg[21] ),
        .\sp_reg[23] (\sp_reg[23] ),
        .\sp_reg[27] (\sp_reg[27] ),
        .\sp_reg[27]_0 (\sp_reg[27]_0 ),
        .\sp_reg[28] (\sp_reg[28] ),
        .\sp_reg[29] (\sp_reg[29] ),
        .\sp_reg[31] (\sp_reg[31] ),
        .\sr_reg[8] (\sr_reg[8] ),
        .\tr_reg[27] (\tr_reg[27] ));
endmodule

module niho_mem_bctl
   (D,
    \cbus_i[31] ,
    \read_cyc_reg[2]_0 ,
    \read_cyc_reg[1]_0 ,
    .bdatr_0_sp_1(bdatr_0_sn_1),
    .bdatr_1_sp_1(bdatr_1_sn_1),
    .bdatr_2_sp_1(bdatr_2_sn_1),
    .bdatr_3_sp_1(bdatr_3_sn_1),
    .bdatr_4_sp_1(bdatr_4_sn_1),
    .bdatr_5_sp_1(bdatr_5_sn_1),
    .bdatr_6_sp_1(bdatr_6_sn_1),
    .bdatr_7_sp_1(bdatr_7_sn_1),
    \read_cyc_reg[1]_1 ,
    .bdatr_8_sp_1(bdatr_8_sn_1),
    \read_cyc_reg[0]_0 ,
    .bdatr_9_sp_1(bdatr_9_sn_1),
    .bdatr_10_sp_1(bdatr_10_sn_1),
    .bdatr_11_sp_1(bdatr_11_sn_1),
    .bdatr_12_sp_1(bdatr_12_sn_1),
    .bdatr_13_sp_1(bdatr_13_sn_1),
    .bdatr_14_sp_1(bdatr_14_sn_1),
    .bdatr_15_sp_1(bdatr_15_sn_1),
    \sr_reg[8] ,
    \sp_reg[27] ,
    \sp_reg[31] ,
    \sp_reg[23] ,
    \sp_reg[29] ,
    \sp_reg[28] ,
    \sp_reg[21] ,
    \sp_reg[19] ,
    \sp_reg[27]_0 ,
    \tr_reg[27] ,
    cbus_i,
    bdatr,
    p_2_in,
    out,
    \grn_reg[15] ,
    bcmd,
    brdy,
    p_0_in,
    clk,
    \read_cyc_reg[0]_1 );
  output [6:0]D;
  output [6:0]\cbus_i[31] ;
  output \read_cyc_reg[2]_0 ;
  output \read_cyc_reg[1]_0 ;
  output \read_cyc_reg[1]_1 ;
  output \read_cyc_reg[0]_0 ;
  output [6:0]\sr_reg[8] ;
  input [0:0]\sp_reg[27] ;
  input \sp_reg[31] ;
  input \sp_reg[23] ;
  input \sp_reg[29] ;
  input \sp_reg[28] ;
  input \sp_reg[21] ;
  input \sp_reg[19] ;
  input \sp_reg[27]_0 ;
  input \tr_reg[27] ;
  input [6:0]cbus_i;
  input [22:0]bdatr;
  input [6:0]p_2_in;
  input [0:0]out;
  input [6:0]\grn_reg[15] ;
  input [1:0]bcmd;
  input brdy;
  input p_0_in;
  input clk;
  input \read_cyc_reg[0]_1 ;
  output bdatr_0_sn_1;
  output bdatr_1_sn_1;
  output bdatr_2_sn_1;
  output bdatr_3_sn_1;
  output bdatr_4_sn_1;
  output bdatr_5_sn_1;
  output bdatr_6_sn_1;
  output bdatr_7_sn_1;
  output bdatr_8_sn_1;
  output bdatr_9_sn_1;
  output bdatr_10_sn_1;
  output bdatr_11_sn_1;
  output bdatr_12_sn_1;
  output bdatr_13_sn_1;
  output bdatr_14_sn_1;
  output bdatr_15_sn_1;

  wire \<const1> ;
  wire [6:0]D;
  wire [1:0]bcmd;
  wire [22:0]bdatr;
  wire bdatr_0_sn_1;
  wire bdatr_10_sn_1;
  wire bdatr_11_sn_1;
  wire bdatr_12_sn_1;
  wire bdatr_13_sn_1;
  wire bdatr_14_sn_1;
  wire bdatr_15_sn_1;
  wire bdatr_1_sn_1;
  wire bdatr_2_sn_1;
  wire bdatr_3_sn_1;
  wire bdatr_4_sn_1;
  wire bdatr_5_sn_1;
  wire bdatr_6_sn_1;
  wire bdatr_7_sn_1;
  wire bdatr_8_sn_1;
  wire bdatr_9_sn_1;
  wire brdy;
  wire [6:0]cbus_i;
  wire [6:0]\cbus_i[31] ;
  wire clk;
  wire [6:0]\grn_reg[15] ;
  wire [0:0]out;
  wire p_0_in;
  wire [6:0]p_2_in;
  wire \read_cyc[1]_i_1_n_0 ;
  wire \read_cyc[2]_i_1_n_0 ;
  wire \read_cyc_reg[0]_0 ;
  wire \read_cyc_reg[0]_1 ;
  wire \read_cyc_reg[1]_0 ;
  wire \read_cyc_reg[1]_1 ;
  wire \read_cyc_reg[2]_0 ;
  wire \sp_reg[19] ;
  wire \sp_reg[21] ;
  wire \sp_reg[23] ;
  wire [0:0]\sp_reg[27] ;
  wire \sp_reg[27]_0 ;
  wire \sp_reg[28] ;
  wire \sp_reg[29] ;
  wire \sp_reg[31] ;
  wire [6:0]\sr_reg[8] ;
  wire \tr_reg[27] ;

  VCC VCC
       (.P(\<const1> ));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[11]_i_1 
       (.I0(\cbus_i[31] [3]),
        .I1(out),
        .I2(\grn_reg[15] [3]),
        .O(\sr_reg[8] [3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[12]_i_1 
       (.I0(\cbus_i[31] [4]),
        .I1(out),
        .I2(\grn_reg[15] [4]),
        .O(\sr_reg[8] [4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[13]_i_1 
       (.I0(\cbus_i[31] [5]),
        .I1(out),
        .I2(\grn_reg[15] [5]),
        .O(\sr_reg[8] [5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[15]_i_2 
       (.I0(\cbus_i[31] [6]),
        .I1(out),
        .I2(\grn_reg[15] [6]),
        .O(\sr_reg[8] [6]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[3]_i_1 
       (.I0(\cbus_i[31] [0]),
        .I1(out),
        .I2(\grn_reg[15] [0]),
        .O(\sr_reg[8] [0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[5]_i_1 
       (.I0(\cbus_i[31] [1]),
        .I1(out),
        .I2(\grn_reg[15] [1]),
        .O(\sr_reg[8] [1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \bank02/grn[7]_i_1 
       (.I0(\cbus_i[31] [2]),
        .I1(out),
        .I2(\grn_reg[15] [2]),
        .O(\sr_reg[8] [2]));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[0]_i_4 
       (.I0(bdatr[0]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_0_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[0]_i_5 
       (.I0(bdatr[8]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[0]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_8_sn_1));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[15]_i_7 
       (.I0(\read_cyc_reg[1]_0 ),
        .I1(\read_cyc_reg[2]_0 ),
        .O(\read_cyc_reg[1]_1 ));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[1]_i_4 
       (.I0(bdatr[1]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_1_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[1]_i_5 
       (.I0(bdatr[9]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[1]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_9_sn_1));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[2]_i_4 
       (.I0(bdatr[2]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_2_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[2]_i_5 
       (.I0(bdatr[10]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[2]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_10_sn_1));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[3]_i_4 
       (.I0(bdatr[3]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_3_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[3]_i_5 
       (.I0(bdatr[11]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[3]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_11_sn_1));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[4]_i_4 
       (.I0(bdatr[4]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_4_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[4]_i_5 
       (.I0(bdatr[12]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[4]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_12_sn_1));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[5]_i_4 
       (.I0(bdatr[5]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_5_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[5]_i_5 
       (.I0(bdatr[13]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[5]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_13_sn_1));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[6]_i_4 
       (.I0(bdatr[6]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_6_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[6]_i_5 
       (.I0(bdatr[14]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[6]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_14_sn_1));
  LUT3 #(
    .INIT(8'h08)) 
    \iv[7]_i_4 
       (.I0(bdatr[7]),
        .I1(\read_cyc_reg[2]_0 ),
        .I2(\read_cyc_reg[1]_0 ),
        .O(bdatr_7_sn_1));
  LUT5 #(
    .INIT(32'hE2000000)) 
    \iv[7]_i_5 
       (.I0(bdatr[15]),
        .I1(\read_cyc_reg[0]_0 ),
        .I2(bdatr[7]),
        .I3(\read_cyc_reg[1]_0 ),
        .I4(\read_cyc_reg[2]_0 ),
        .O(bdatr_15_sn_1));
  LUT3 #(
    .INIT(8'hB8)) 
    \read_cyc[1]_i_1 
       (.I0(bcmd[1]),
        .I1(brdy),
        .I2(\read_cyc_reg[1]_0 ),
        .O(\read_cyc[1]_i_1_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \read_cyc[2]_i_1 
       (.I0(bcmd[0]),
        .I1(brdy),
        .I2(\read_cyc_reg[2]_0 ),
        .O(\read_cyc[2]_i_1_n_0 ));
  FDRE \read_cyc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\read_cyc_reg[0]_1 ),
        .Q(\read_cyc_reg[0]_0 ),
        .R(p_0_in));
  FDRE \read_cyc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\read_cyc[1]_i_1_n_0 ),
        .Q(\read_cyc_reg[1]_0 ),
        .R(p_0_in));
  FDRE \read_cyc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\read_cyc[2]_i_1_n_0 ),
        .Q(\read_cyc_reg[2]_0 ),
        .R(p_0_in));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[19]_i_1 
       (.I0(\cbus_i[31] [0]),
        .I1(\sp_reg[27] ),
        .I2(\sp_reg[19] ),
        .O(D[0]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[21]_i_1 
       (.I0(\cbus_i[31] [1]),
        .I1(\sp_reg[27] ),
        .I2(\sp_reg[21] ),
        .O(D[1]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[23]_i_1 
       (.I0(\cbus_i[31] [2]),
        .I1(\sp_reg[27] ),
        .I2(\sp_reg[23] ),
        .O(D[2]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[27]_i_1 
       (.I0(\cbus_i[31] [3]),
        .I1(\sp_reg[27] ),
        .I2(\sp_reg[27]_0 ),
        .O(D[3]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[28]_i_1 
       (.I0(\cbus_i[31] [4]),
        .I1(\sp_reg[27] ),
        .I2(\sp_reg[28] ),
        .O(D[4]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[29]_i_1 
       (.I0(\cbus_i[31] [5]),
        .I1(\sp_reg[27] ),
        .I2(\sp_reg[29] ),
        .O(D[5]));
  LUT3 #(
    .INIT(8'hB8)) 
    \sp[31]_i_1 
       (.I0(\cbus_i[31] [6]),
        .I1(\sp_reg[27] ),
        .I2(\sp_reg[31] ),
        .O(D[6]));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[19]_i_1 
       (.I0(\tr_reg[27] ),
        .I1(cbus_i[0]),
        .I2(bdatr[16]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(p_2_in[0]),
        .O(\cbus_i[31] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[21]_i_1 
       (.I0(\tr_reg[27] ),
        .I1(cbus_i[1]),
        .I2(bdatr[17]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(p_2_in[1]),
        .O(\cbus_i[31] [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[23]_i_1 
       (.I0(\tr_reg[27] ),
        .I1(cbus_i[2]),
        .I2(bdatr[18]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(p_2_in[2]),
        .O(\cbus_i[31] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[27]_i_1 
       (.I0(\tr_reg[27] ),
        .I1(cbus_i[3]),
        .I2(bdatr[19]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(p_2_in[3]),
        .O(\cbus_i[31] [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[28]_i_1 
       (.I0(\tr_reg[27] ),
        .I1(cbus_i[4]),
        .I2(bdatr[20]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(p_2_in[4]),
        .O(\cbus_i[31] [4]));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[29]_i_1 
       (.I0(\tr_reg[27] ),
        .I1(cbus_i[5]),
        .I2(bdatr[21]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(p_2_in[5]),
        .O(\cbus_i[31] [5]));
  LUT6 #(
    .INIT(64'hFFFFFFFF8888F888)) 
    \tr[31]_i_2 
       (.I0(\tr_reg[27] ),
        .I1(cbus_i[6]),
        .I2(bdatr[22]),
        .I3(\read_cyc_reg[2]_0 ),
        .I4(\read_cyc_reg[1]_0 ),
        .I5(p_2_in[6]),
        .O(\cbus_i[31] [6]));
endmodule

module niho_rgf
   (out,
    \sp_reg[0] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \sp_reg[5] ,
    \sp_reg[6] ,
    \sp_reg[7] ,
    \sp_reg[8] ,
    \sp_reg[9] ,
    \sp_reg[10] ,
    \sp_reg[11] ,
    \sp_reg[12] ,
    \sp_reg[13] ,
    \sp_reg[14] ,
    \sp_reg[15] ,
    \sp_reg[16] ,
    \sp_reg[17] ,
    \sp_reg[18] ,
    \sp_reg[19] ,
    \sp_reg[20] ,
    \sp_reg[21] ,
    \sp_reg[22] ,
    \sp_reg[23] ,
    \sp_reg[24] ,
    \sp_reg[25] ,
    \sp_reg[26] ,
    \sp_reg[27] ,
    \sp_reg[28] ,
    \sp_reg[29] ,
    \sp_reg[30] ,
    \sp_reg[31] ,
    O,
    \sr_reg[8] ,
    \art/add/sr[5]_i_14 ,
    p_2_in,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \badr[21]_INST_0_i_1 ,
    \tr_reg[5] ,
    abus_0,
    \bdatw[8]_INST_0_i_2 ,
    \iv[7]_i_33 ,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr[4]_i_21 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr[4]_i_147 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \iv[13]_i_10 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr[4]_i_65 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \iv[13]_i_27 ,
    \sr_reg[8]_26 ,
    \iv[8]_i_20 ,
    \sr_reg[8]_27 ,
    \iv[14]_i_35 ,
    \sr_reg[8]_28 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr[4]_i_116 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \sr_reg[8]_33 ,
    \tr[17]_i_9 ,
    \tr[24]_i_10 ,
    \tr[30]_i_10 ,
    \tr[20]_i_9 ,
    \tr[22]_i_9 ,
    \tr[18]_i_9 ,
    \tr[26]_i_9 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \sr_reg[8]_36 ,
    \sr_reg[8]_37 ,
    alu_sr_flag,
    \sr_reg[8]_38 ,
    \sr_reg[8]_39 ,
    \iv[7]_i_17 ,
    \sr_reg[8]_40 ,
    \iv[11]_i_11 ,
    \sr_reg[8]_41 ,
    \sr_reg[8]_42 ,
    \sr_reg[8]_43 ,
    \iv[10]_i_10 ,
    \iv[10]_i_9 ,
    \sr_reg[8]_44 ,
    \sr_reg[8]_45 ,
    \sr_reg[8]_46 ,
    \iv[14]_i_11 ,
    \sr_reg[8]_47 ,
    \iv[9]_i_11 ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    \iv[14]_i_49 ,
    \sr_reg[8]_50 ,
    \sr_reg[8]_51 ,
    \iv[0]_i_25 ,
    \iv[4]_i_35 ,
    \sr_reg[8]_52 ,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    \sr_reg[8]_57 ,
    \sr_reg[8]_58 ,
    \sr_reg[8]_59 ,
    \sr_reg[8]_60 ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    \sr_reg[8]_63 ,
    \sr_reg[8]_64 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    \sr_reg[8]_67 ,
    \sr_reg[8]_68 ,
    \sr_reg[8]_69 ,
    \sr_reg[8]_70 ,
    \sr_reg[8]_71 ,
    \sr_reg[8]_72 ,
    \sr_reg[8]_73 ,
    \sr_reg[8]_74 ,
    \sr_reg[8]_75 ,
    \sr_reg[8]_76 ,
    \sr_reg[8]_77 ,
    \sr_reg[8]_78 ,
    \sr_reg[8]_79 ,
    \iv[8]_i_34 ,
    \sr_reg[8]_80 ,
    \sr_reg[8]_81 ,
    \sr_reg[8]_82 ,
    \sr_reg[8]_83 ,
    \sr_reg[8]_84 ,
    \sr_reg[8]_85 ,
    \sr_reg[8]_86 ,
    \sr_reg[8]_87 ,
    \sr_reg[8]_88 ,
    \sr_reg[8]_89 ,
    \sr_reg[8]_90 ,
    \sr_reg[8]_91 ,
    \sr_reg[8]_92 ,
    \sr_reg[8]_93 ,
    \sr_reg[8]_94 ,
    \sr_reg[8]_95 ,
    \sr_reg[8]_96 ,
    \sr_reg[8]_97 ,
    \sr_reg[8]_98 ,
    \sr_reg[8]_99 ,
    \sr_reg[8]_100 ,
    \sr_reg[8]_101 ,
    \sr_reg[8]_102 ,
    \sr_reg[8]_103 ,
    \iv[7]_i_25 ,
    \sr_reg[8]_104 ,
    \sr_reg[8]_105 ,
    \sr_reg[8]_106 ,
    \sr_reg[6] ,
    \sr_reg[8]_107 ,
    \badr[0]_INST_0_i_1 ,
    \sr_reg[8]_108 ,
    \sr_reg[8]_109 ,
    \sr_reg[8]_110 ,
    \sr_reg[8]_111 ,
    \sr_reg[6]_0 ,
    \sr_reg[8]_112 ,
    \sr_reg[8]_113 ,
    \sr_reg[8]_114 ,
    \sr_reg[6]_1 ,
    \sr_reg[8]_115 ,
    \sr_reg[8]_116 ,
    \sr_reg[8]_117 ,
    \sr_reg[8]_118 ,
    \sr_reg[8]_119 ,
    \sr_reg[8]_120 ,
    \sr_reg[8]_121 ,
    \sr_reg[8]_122 ,
    \sr_reg[8]_123 ,
    \sr_reg[8]_124 ,
    \sr_reg[8]_125 ,
    \sr_reg[8]_126 ,
    \sr_reg[6]_2 ,
    \sr_reg[8]_127 ,
    \sr_reg[6]_3 ,
    \sr_reg[8]_128 ,
    \sr_reg[8]_129 ,
    \badr[5]_INST_0_i_1 ,
    \sp_reg[4]_0 ,
    \sr_reg[4] ,
    \grn_reg[4] ,
    \niho_dsp_a[15]_INST_0_i_3 ,
    niho_dsp_a,
    \iv[15]_i_108 ,
    \sr_reg[8]_130 ,
    \iv[15]_i_108_0 ,
    \iv[15]_i_108_1 ,
    \iv[15]_i_108_2 ,
    \iv[15]_i_108_3 ,
    \sr_reg[8]_131 ,
    \iv[15]_i_108_4 ,
    \sr_reg[8]_132 ,
    \iv[15]_i_108_5 ,
    \sr_reg[8]_133 ,
    \iv[15]_i_108_6 ,
    \sr_reg[8]_134 ,
    \sr_reg[8]_135 ,
    \badr[5]_INST_0_i_1_0 ,
    \sr_reg[8]_136 ,
    \iv[15]_i_108_7 ,
    \sr_reg[8]_137 ,
    \sr_reg[8]_138 ,
    \iv[15]_i_108_8 ,
    \badr[1]_INST_0_i_1 ,
    \sr_reg[8]_139 ,
    \badr[0]_INST_0_i_1_0 ,
    \iv[15]_i_108_9 ,
    mul_a_i,
    \iv[15]_i_108_10 ,
    \iv[15]_i_108_11 ,
    \iv[15]_i_108_12 ,
    \iv[15]_i_108_13 ,
    \iv[15]_i_108_14 ,
    \iv[15]_i_108_15 ,
    \iv[15]_i_108_16 ,
    \iv[15]_i_108_17 ,
    \iv[15]_i_108_18 ,
    \iv[15]_i_108_19 ,
    \iv[15]_i_108_20 ,
    \iv[15]_i_108_21 ,
    \iv[15]_i_108_22 ,
    \sr_reg[8]_140 ,
    \iv[15]_i_108_23 ,
    mul_rslt0,
    \sr_reg[8]_141 ,
    \art/add/iv[7]_i_32 ,
    \sr_reg[6]_4 ,
    \art/add/sr[5]_i_18 ,
    \sr_reg[8]_142 ,
    \sr_reg[8]_143 ,
    \sr_reg[8]_144 ,
    \sr_reg[8]_145 ,
    \sr_reg[8]_146 ,
    \sr_reg[8]_147 ,
    \sr_reg[8]_148 ,
    \sr_reg[8]_149 ,
    \sr_reg[8]_150 ,
    fch_pc,
    rgf_pc,
    abus_o,
    fch_irq_req,
    .irq_lev_0_sp_1(irq_lev_0_sn_1),
    \sr_reg[7] ,
    \sr_reg[5] ,
    \sr_reg[7]_0 ,
    \sr_reg[4]_0 ,
    \sr_reg[7]_1 ,
    \sr_reg[4]_1 ,
    \sr_reg[6]_5 ,
    \sr_reg[7]_2 ,
    \sr_reg[8]_151 ,
    bbus_o,
    \sr_reg[8]_152 ,
    \sr_reg[8]_153 ,
    \sr_reg[8]_154 ,
    \sr_reg[8]_155 ,
    \sr_reg[8]_156 ,
    \sr_reg[8]_157 ,
    \stat_reg[0] ,
    .irq_lev_1_sp_1(irq_lev_1_sn_1),
    \sr_reg[5]_0 ,
    \sr_reg[6]_6 ,
    \sr_reg[6]_7 ,
    \sr_reg[6]_8 ,
    \sr_reg[8]_158 ,
    \sr_reg[8]_159 ,
    \sr_reg[8]_160 ,
    \badr[6]_INST_0_i_1 ,
    \sr_reg[8]_161 ,
    \badr[4]_INST_0_i_1 ,
    \sr[6]_i_13 ,
    \sr_reg[8]_162 ,
    \sr_reg[8]_163 ,
    \badr[2]_INST_0_i_1 ,
    niho_dsp_b,
    \sr_reg[8]_164 ,
    \sr_reg[8]_165 ,
    \sr_reg[8]_166 ,
    \sr_reg[8]_167 ,
    p_0_in,
    \iv_reg[15] ,
    \iv_reg[15]_0 ,
    \tr_reg[31] ,
    \iv_reg[14] ,
    \iv_reg[13] ,
    \iv_reg[12] ,
    \iv_reg[11] ,
    \iv_reg[10] ,
    \iv_reg[9] ,
    \iv_reg[8] ,
    \iv_reg[7] ,
    \iv_reg[6] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \sr_reg[15] ,
    \sr_reg[14] ,
    \sr_reg[13] ,
    \sr_reg[12] ,
    \sr_reg[11] ,
    \sr_reg[10] ,
    \sr_reg[9] ,
    \sr_reg[8]_168 ,
    \sr_reg[7]_3 ,
    \sr_reg[6]_9 ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sp_reg[31]_0 ,
    \sp_reg[30]_0 ,
    \sp_reg[29]_0 ,
    \sp_reg[28]_0 ,
    \sp_reg[27]_0 ,
    \sp_reg[26]_0 ,
    \sp_reg[25]_0 ,
    \sp_reg[24]_0 ,
    \sp_reg[23]_0 ,
    \sp_reg[22]_0 ,
    \sp_reg[21]_0 ,
    \sp_reg[20]_0 ,
    \sp_reg[19]_0 ,
    \sp_reg[18]_0 ,
    \sp_reg[17]_0 ,
    \sp_reg[16]_0 ,
    \tr_reg[31]_0 ,
    \tr_reg[30] ,
    \tr_reg[29] ,
    \tr_reg[28] ,
    \tr_reg[27] ,
    \tr_reg[26] ,
    \tr_reg[25] ,
    \tr_reg[24] ,
    \tr_reg[23] ,
    \tr_reg[22] ,
    \tr_reg[21] ,
    \tr_reg[20] ,
    \tr_reg[19] ,
    \tr_reg[18] ,
    \tr_reg[17] ,
    \tr_reg[16] ,
    \sp_reg[1]_0 ,
    \sp_reg[2]_0 ,
    \sp_reg[3]_0 ,
    D,
    rst_n,
    \sr_reg[15]_0 ,
    abus_sel_cr,
    ctl_sp_id4,
    ctl_sp_inc,
    ctl_sp_dec,
    cbus_sel_0,
    \sr_reg[5]_1 ,
    \sr_reg[6]_10 ,
    \tr_reg[31]_1 ,
    \tr_reg[31]_2 ,
    \tr_reg[27]_0 ,
    niho_dsp_c,
    \tr_reg[23]_0 ,
    \tr_reg[29]_0 ,
    \tr_reg[28]_0 ,
    \tr_reg[21]_0 ,
    \tr_reg[19]_0 ,
    \tr_reg[27]_1 ,
    bbus_0,
    \iv[13]_i_17 ,
    \iv[13]_i_17_0 ,
    \iv[7]_i_7 ,
    \iv[7]_i_7_0 ,
    \iv[7]_i_7_1 ,
    \tr_reg[1] ,
    \tr_reg[1]_0 ,
    \sr_reg[4]_2 ,
    \sr_reg[4]_3 ,
    \sr[4]_i_5 ,
    \sr[4]_i_5_0 ,
    \sr[4]_i_16 ,
    \sr[4]_i_89 ,
    \sr[4]_i_5_1 ,
    \sr[4]_i_21_0 ,
    \sr[4]_i_21_1 ,
    \tr[19]_i_3 ,
    \sr[4]_i_5_2 ,
    \sr[4]_i_20 ,
    \sr[4]_i_20_0 ,
    \iv[13]_i_2 ,
    \sr[4]_i_20_1 ,
    \sr[4]_i_20_2 ,
    \iv[12]_i_2 ,
    \sr[4]_i_44 ,
    \iv[0]_i_3 ,
    \iv[10]_i_2 ,
    \sr[4]_i_16_0 ,
    \sr[4]_i_33 ,
    \sr[4]_i_39 ,
    \iv[8]_i_2 ,
    \sr[4]_i_40 ,
    \tr[22]_i_3 ,
    \tr[24]_i_2 ,
    \tr[24]_i_3 ,
    \tr[23]_i_2 ,
    \tr[17]_i_2 ,
    \tr[21]_i_2 ,
    \tr[22]_i_2 ,
    \tr[20]_i_2 ,
    \tr[18]_i_2 ,
    \tr[28]_i_2 ,
    \tr[25]_i_2 ,
    \tr[19]_i_2 ,
    \iv[15]_i_8 ,
    \iv[15]_i_8_0 ,
    \iv[15]_i_8_1 ,
    \tr[19]_i_3_0 ,
    \sr_reg[6]_11 ,
    \sr[4]_i_36 ,
    \sr[5]_i_3 ,
    \tr[30]_i_3 ,
    \tr[30]_i_3_0 ,
    \tr[26]_i_3 ,
    \tr[29]_i_3 ,
    \sr[4]_i_42 ,
    \sr[4]_i_43 ,
    \iv[0]_i_3_0 ,
    \iv[5]_i_3 ,
    \iv[4]_i_3 ,
    \sr[4]_i_39_0 ,
    \sr[4]_i_40_0 ,
    \sr[4]_i_37 ,
    \sr[6]_i_4 ,
    \iv[0]_i_3_1 ,
    \iv[0]_i_10 ,
    \iv[15]_i_8_2 ,
    \iv[1]_i_10 ,
    \iv[1]_i_10_0 ,
    \iv[1]_i_10_1 ,
    \iv[3]_i_10 ,
    \iv[3]_i_10_0 ,
    \iv[3]_i_10_1 ,
    \sr[4]_i_45 ,
    \sr[4]_i_44_0 ,
    \sr[4]_i_35 ,
    \iv[6]_i_10 ,
    \iv[6]_i_10_0 ,
    \iv[6]_i_10_1 ,
    \iv[0]_i_10_0 ,
    \sr[6]_i_12 ,
    \sr[6]_i_12_0 ,
    \tr[16]_i_6 ,
    \tr[16]_i_6_0 ,
    \iv[7]_i_9 ,
    \sr[4]_i_43_0 ,
    \iv[1]_i_9 ,
    \iv[2]_i_9 ,
    \iv[3]_i_9 ,
    \sr[4]_i_45_0 ,
    \sr[4]_i_44_1 ,
    \iv[10]_i_5 ,
    \iv[5]_i_9 ,
    \iv[4]_i_9 ,
    \iv[8]_i_5 ,
    \iv[14]_i_5 ,
    \iv[9]_i_5 ,
    \sr[4]_i_38 ,
    \tr[21]_i_3 ,
    \tr[20]_i_3 ,
    \tr[24]_i_3_0 ,
    \iv[0]_i_10_1 ,
    \sr[4]_i_87 ,
    \sr[6]_i_11 ,
    \sr[4]_i_41 ,
    \iv[0]_i_19 ,
    \iv[7]_i_3 ,
    \sr[4]_i_61 ,
    \sr[4]_i_139 ,
    \mul_b_reg[5] ,
    \mul_b_reg[5]_0 ,
    \iv[0]_i_7 ,
    \iv[15]_i_96 ,
    \iv[15]_i_96_0 ,
    \mul_b_reg[0] ,
    \mul_b_reg[0]_0 ,
    mul_rslt,
    mul_a,
    \niho_dsp_b[5] ,
    \mul_a_reg[15] ,
    \tr[22]_i_11 ,
    \remden_reg[26] ,
    \remden_reg[29] ,
    \remden_reg[25] ,
    \remden_reg[24] ,
    \remden_reg[23] ,
    \remden_reg[22] ,
    \remden_reg[21] ,
    \remden_reg[20] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] ,
    Q,
    \tr[19]_i_2_0 ,
    \tr[29]_i_2 ,
    \tr[19]_i_2_1 ,
    \sr[4]_i_3 ,
    \iv[0]_i_6 ,
    \iv[0]_i_6_0 ,
    \iv[4]_i_6 ,
    \iv[8]_i_8 ,
    S,
    .abus_o_16_sp_1(abus_o_16_sn_1),
    irq,
    irq_lev,
    \badr[31]_INST_0_i_69 ,
    \stat_reg[1] ,
    \stat[0]_i_6 ,
    \sr[4]_i_19 ,
    \sr[4]_i_18 ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    bbus_sel_0,
    abus_sel_0,
    \mul_a_reg[32] ,
    \remden_reg[19] ,
    \sr[5]_i_2 ,
    \tr_reg[31]_i_13 ,
    \remden_reg[30] ,
    \tr_reg[31]_i_13_0 ,
    \tr_reg[31]_i_13_1 ,
    \remden_reg[28] ,
    \tr_reg[31]_i_32 ,
    \remden_reg[27] ,
    \tr_reg[31]_i_32_0 ,
    \remden_reg[26]_0 ,
    \tr_reg[31]_i_32_1 ,
    \tr_reg[31]_i_32_2 ,
    \tr_reg[23]_i_11 ,
    \tr_reg[23]_i_11_0 ,
    \tr_reg[23]_i_11_1 ,
    \tr_reg[23]_i_11_2 ,
    \sr_reg[6]_i_6 ,
    \sr_reg[6]_i_6_0 ,
    \sr_reg[6]_i_6_1 ,
    .niho_dsp_b_0_sp_1(niho_dsp_b_0_sn_1),
    \niho_dsp_b[5]_0 ,
    \i_/bdatw[15]_INST_0_i_65 ,
    ctl_selb_rn,
    \i_/bdatw[15]_INST_0_i_65_0 ,
    \i_/bdatw[15]_INST_0_i_65_1 ,
    ctl_selb_0,
    \i_/bdatw[15]_INST_0_i_65_2 ,
    \i_/bdatw[15]_INST_0_i_67 ,
    \i_/bdatw[15]_INST_0_i_27 ,
    \i_/bdatw[15]_INST_0_i_67_0 ,
    \i_/bdatw[15]_INST_0_i_27_0 ,
    clk,
    \sr_reg[11]_0 ,
    \sr_reg[10]_0 ,
    \sr_reg[8]_169 ,
    \sr_reg[7]_4 ,
    \sr_reg[6]_12 ,
    \sr_reg[5]_2 ,
    \sr_reg[4]_4 ,
    \sr_reg[3]_0 ,
    \sr_reg[2]_0 ,
    \sr_reg[1]_0 ,
    \sr_reg[0] ,
    \sp_reg[31]_1 ,
    \mul_a_reg[14] ,
    \mul_a_reg[13] ,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \mul_a_reg[4] ,
    \mul_a_reg[3] ,
    \mul_a_reg[2] ,
    \mul_a_reg[1] ,
    \mul_a_reg[0] ,
    \mul_a_reg[32]_0 ,
    \mul_a_reg[30] ,
    \mul_a_reg[29] ,
    \mul_a_reg[28] ,
    \mul_a_reg[27] ,
    \mul_a_reg[26] ,
    \mul_a_reg[25] ,
    \mul_a_reg[24] ,
    \mul_a_reg[23] ,
    \mul_a_reg[22] ,
    \mul_a_reg[21] ,
    \mul_a_reg[20] ,
    \mul_a_reg[19] ,
    \mul_a_reg[18] ,
    \mul_a_reg[17] ,
    \mul_a_reg[16] ,
    bbus_sel_cr,
    bbus_sr,
    E,
    cbus,
    \grn_reg[15] ,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    \grn_reg[15]_2 ,
    \grn_reg[15]_3 ,
    \grn_reg[15]_4 ,
    \grn_reg[15]_5 ,
    \grn_reg[15]_6 ,
    \grn_reg[15]_7 ,
    \grn_reg[15]_8 ,
    \grn_reg[15]_9 ,
    \grn_reg[15]_10 ,
    \grn_reg[15]_11 ,
    \grn_reg[15]_12 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[15]_22 ,
    \pc_reg[15] ,
    \tr_reg[0] );
  output [12:0]out;
  output [0:0]\sp_reg[0] ;
  output \sp_reg[1] ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  output \sp_reg[5] ;
  output \sp_reg[6] ;
  output \sp_reg[7] ;
  output \sp_reg[8] ;
  output \sp_reg[9] ;
  output \sp_reg[10] ;
  output \sp_reg[11] ;
  output \sp_reg[12] ;
  output \sp_reg[13] ;
  output \sp_reg[14] ;
  output \sp_reg[15] ;
  output \sp_reg[16] ;
  output \sp_reg[17] ;
  output \sp_reg[18] ;
  output \sp_reg[19] ;
  output \sp_reg[20] ;
  output \sp_reg[21] ;
  output \sp_reg[22] ;
  output \sp_reg[23] ;
  output \sp_reg[24] ;
  output \sp_reg[25] ;
  output \sp_reg[26] ;
  output \sp_reg[27] ;
  output \sp_reg[28] ;
  output \sp_reg[29] ;
  output \sp_reg[30] ;
  output \sp_reg[31] ;
  output [0:0]O;
  output \sr_reg[8] ;
  output [3:0]\art/add/sr[5]_i_14 ;
  output [6:0]p_2_in;
  output \sr_reg[8]_0 ;
  output [0:0]\sr_reg[8]_1 ;
  output \badr[21]_INST_0_i_1 ;
  output [1:0]\tr_reg[5] ;
  output [31:0]abus_0;
  output \bdatw[8]_INST_0_i_2 ;
  output \iv[7]_i_33 ;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr[4]_i_21 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr[4]_i_147 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \iv[13]_i_10 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr[4]_i_65 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \iv[13]_i_27 ;
  output \sr_reg[8]_26 ;
  output \iv[8]_i_20 ;
  output \sr_reg[8]_27 ;
  output \iv[14]_i_35 ;
  output \sr_reg[8]_28 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr[4]_i_116 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \sr_reg[8]_33 ;
  output \tr[17]_i_9 ;
  output \tr[24]_i_10 ;
  output \tr[30]_i_10 ;
  output \tr[20]_i_9 ;
  output \tr[22]_i_9 ;
  output \tr[18]_i_9 ;
  output \tr[26]_i_9 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \sr_reg[8]_36 ;
  output \sr_reg[8]_37 ;
  output [0:0]alu_sr_flag;
  output \sr_reg[8]_38 ;
  output \sr_reg[8]_39 ;
  output \iv[7]_i_17 ;
  output \sr_reg[8]_40 ;
  output \iv[11]_i_11 ;
  output \sr_reg[8]_41 ;
  output \sr_reg[8]_42 ;
  output \sr_reg[8]_43 ;
  output \iv[10]_i_10 ;
  output \iv[10]_i_9 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[8]_45 ;
  output \sr_reg[8]_46 ;
  output \iv[14]_i_11 ;
  output \sr_reg[8]_47 ;
  output \iv[9]_i_11 ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output \iv[14]_i_49 ;
  output \sr_reg[8]_50 ;
  output \sr_reg[8]_51 ;
  output \iv[0]_i_25 ;
  output \iv[4]_i_35 ;
  output \sr_reg[8]_52 ;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output \sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output \sr_reg[8]_57 ;
  output \sr_reg[8]_58 ;
  output \sr_reg[8]_59 ;
  output \sr_reg[8]_60 ;
  output \sr_reg[8]_61 ;
  output \sr_reg[8]_62 ;
  output \sr_reg[8]_63 ;
  output \sr_reg[8]_64 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output \sr_reg[8]_67 ;
  output \sr_reg[8]_68 ;
  output \sr_reg[8]_69 ;
  output \sr_reg[8]_70 ;
  output \sr_reg[8]_71 ;
  output \sr_reg[8]_72 ;
  output \sr_reg[8]_73 ;
  output \sr_reg[8]_74 ;
  output \sr_reg[8]_75 ;
  output \sr_reg[8]_76 ;
  output \sr_reg[8]_77 ;
  output \sr_reg[8]_78 ;
  output \sr_reg[8]_79 ;
  output \iv[8]_i_34 ;
  output \sr_reg[8]_80 ;
  output \sr_reg[8]_81 ;
  output \sr_reg[8]_82 ;
  output \sr_reg[8]_83 ;
  output \sr_reg[8]_84 ;
  output \sr_reg[8]_85 ;
  output \sr_reg[8]_86 ;
  output \sr_reg[8]_87 ;
  output \sr_reg[8]_88 ;
  output \sr_reg[8]_89 ;
  output \sr_reg[8]_90 ;
  output \sr_reg[8]_91 ;
  output \sr_reg[8]_92 ;
  output \sr_reg[8]_93 ;
  output \sr_reg[8]_94 ;
  output \sr_reg[8]_95 ;
  output \sr_reg[8]_96 ;
  output \sr_reg[8]_97 ;
  output \sr_reg[8]_98 ;
  output \sr_reg[8]_99 ;
  output \sr_reg[8]_100 ;
  output \sr_reg[8]_101 ;
  output \sr_reg[8]_102 ;
  output \sr_reg[8]_103 ;
  output \iv[7]_i_25 ;
  output \sr_reg[8]_104 ;
  output \sr_reg[8]_105 ;
  output \sr_reg[8]_106 ;
  output \sr_reg[6] ;
  output \sr_reg[8]_107 ;
  output \badr[0]_INST_0_i_1 ;
  output \sr_reg[8]_108 ;
  output \sr_reg[8]_109 ;
  output \sr_reg[8]_110 ;
  output \sr_reg[8]_111 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[8]_112 ;
  output \sr_reg[8]_113 ;
  output \sr_reg[8]_114 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[8]_115 ;
  output \sr_reg[8]_116 ;
  output \sr_reg[8]_117 ;
  output \sr_reg[8]_118 ;
  output \sr_reg[8]_119 ;
  output \sr_reg[8]_120 ;
  output \sr_reg[8]_121 ;
  output \sr_reg[8]_122 ;
  output \sr_reg[8]_123 ;
  output \sr_reg[8]_124 ;
  output \sr_reg[8]_125 ;
  output \sr_reg[8]_126 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[8]_127 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[8]_128 ;
  output \sr_reg[8]_129 ;
  output \badr[5]_INST_0_i_1 ;
  output \sp_reg[4]_0 ;
  output \sr_reg[4] ;
  output \grn_reg[4] ;
  output \niho_dsp_a[15]_INST_0_i_3 ;
  output [32:0]niho_dsp_a;
  output \iv[15]_i_108 ;
  output \sr_reg[8]_130 ;
  output \iv[15]_i_108_0 ;
  output \iv[15]_i_108_1 ;
  output \iv[15]_i_108_2 ;
  output \iv[15]_i_108_3 ;
  output \sr_reg[8]_131 ;
  output \iv[15]_i_108_4 ;
  output \sr_reg[8]_132 ;
  output \iv[15]_i_108_5 ;
  output \sr_reg[8]_133 ;
  output \iv[15]_i_108_6 ;
  output \sr_reg[8]_134 ;
  output \sr_reg[8]_135 ;
  output \badr[5]_INST_0_i_1_0 ;
  output \sr_reg[8]_136 ;
  output \iv[15]_i_108_7 ;
  output \sr_reg[8]_137 ;
  output \sr_reg[8]_138 ;
  output \iv[15]_i_108_8 ;
  output \badr[1]_INST_0_i_1 ;
  output \sr_reg[8]_139 ;
  output \badr[0]_INST_0_i_1_0 ;
  output \iv[15]_i_108_9 ;
  output [13:0]mul_a_i;
  output \iv[15]_i_108_10 ;
  output \iv[15]_i_108_11 ;
  output \iv[15]_i_108_12 ;
  output \iv[15]_i_108_13 ;
  output \iv[15]_i_108_14 ;
  output \iv[15]_i_108_15 ;
  output \iv[15]_i_108_16 ;
  output \iv[15]_i_108_17 ;
  output \iv[15]_i_108_18 ;
  output \iv[15]_i_108_19 ;
  output \iv[15]_i_108_20 ;
  output \iv[15]_i_108_21 ;
  output \iv[15]_i_108_22 ;
  output \sr_reg[8]_140 ;
  output \iv[15]_i_108_23 ;
  output mul_rslt0;
  output \sr_reg[8]_141 ;
  output [3:0]\art/add/iv[7]_i_32 ;
  output [3:0]\sr_reg[6]_4 ;
  output [3:0]\art/add/sr[5]_i_18 ;
  output \sr_reg[8]_142 ;
  output \sr_reg[8]_143 ;
  output \sr_reg[8]_144 ;
  output \sr_reg[8]_145 ;
  output \sr_reg[8]_146 ;
  output \sr_reg[8]_147 ;
  output \sr_reg[8]_148 ;
  output \sr_reg[8]_149 ;
  output \sr_reg[8]_150 ;
  output [15:0]fch_pc;
  output [15:0]rgf_pc;
  output [31:0]abus_o;
  output fch_irq_req;
  output \sr_reg[7] ;
  output \sr_reg[5] ;
  output \sr_reg[7]_0 ;
  output \sr_reg[4]_0 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[6]_5 ;
  output \sr_reg[7]_2 ;
  output \sr_reg[8]_151 ;
  output [1:0]bbus_o;
  output \sr_reg[8]_152 ;
  output \sr_reg[8]_153 ;
  output \sr_reg[8]_154 ;
  output \sr_reg[8]_155 ;
  output \sr_reg[8]_156 ;
  output \sr_reg[8]_157 ;
  output \stat_reg[0] ;
  output \sr_reg[5]_0 ;
  output \sr_reg[6]_6 ;
  output \sr_reg[6]_7 ;
  output \sr_reg[6]_8 ;
  output \sr_reg[8]_158 ;
  output [1:0]\sr_reg[8]_159 ;
  output \sr_reg[8]_160 ;
  output \badr[6]_INST_0_i_1 ;
  output \sr_reg[8]_161 ;
  output \badr[4]_INST_0_i_1 ;
  output \sr[6]_i_13 ;
  output \sr_reg[8]_162 ;
  output \sr_reg[8]_163 ;
  output \badr[2]_INST_0_i_1 ;
  output [1:0]niho_dsp_b;
  output \sr_reg[8]_164 ;
  output \sr_reg[8]_165 ;
  output \sr_reg[8]_166 ;
  output \sr_reg[8]_167 ;
  output p_0_in;
  output \iv_reg[15] ;
  output [15:0]\iv_reg[15]_0 ;
  output [31:0]\tr_reg[31] ;
  output \iv_reg[14] ;
  output \iv_reg[13] ;
  output \iv_reg[12] ;
  output \iv_reg[11] ;
  output \iv_reg[10] ;
  output \iv_reg[9] ;
  output \iv_reg[8] ;
  output \iv_reg[7] ;
  output \iv_reg[6] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \sr_reg[15] ;
  output \sr_reg[14] ;
  output \sr_reg[13] ;
  output \sr_reg[12] ;
  output \sr_reg[11] ;
  output \sr_reg[10] ;
  output \sr_reg[9] ;
  output \sr_reg[8]_168 ;
  output \sr_reg[7]_3 ;
  output \sr_reg[6]_9 ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sp_reg[31]_0 ;
  output \sp_reg[30]_0 ;
  output \sp_reg[29]_0 ;
  output \sp_reg[28]_0 ;
  output \sp_reg[27]_0 ;
  output \sp_reg[26]_0 ;
  output \sp_reg[25]_0 ;
  output \sp_reg[24]_0 ;
  output \sp_reg[23]_0 ;
  output \sp_reg[22]_0 ;
  output \sp_reg[21]_0 ;
  output \sp_reg[20]_0 ;
  output \sp_reg[19]_0 ;
  output \sp_reg[18]_0 ;
  output \sp_reg[17]_0 ;
  output \sp_reg[16]_0 ;
  output \tr_reg[31]_0 ;
  output \tr_reg[30] ;
  output \tr_reg[29] ;
  output \tr_reg[28] ;
  output \tr_reg[27] ;
  output \tr_reg[26] ;
  output \tr_reg[25] ;
  output \tr_reg[24] ;
  output \tr_reg[23] ;
  output \tr_reg[22] ;
  output \tr_reg[21] ;
  output \tr_reg[20] ;
  output \tr_reg[19] ;
  output \tr_reg[18] ;
  output \tr_reg[17] ;
  output \tr_reg[16] ;
  output \sp_reg[1]_0 ;
  output \sp_reg[2]_0 ;
  output \sp_reg[3]_0 ;
  input [1:0]D;
  input rst_n;
  input \sr_reg[15]_0 ;
  input [3:0]abus_sel_cr;
  input ctl_sp_id4;
  input ctl_sp_inc;
  input ctl_sp_dec;
  input [0:0]cbus_sel_0;
  input \sr_reg[5]_1 ;
  input \sr_reg[6]_10 ;
  input \tr_reg[31]_1 ;
  input \tr_reg[31]_2 ;
  input \tr_reg[27]_0 ;
  input [5:0]niho_dsp_c;
  input \tr_reg[23]_0 ;
  input \tr_reg[29]_0 ;
  input \tr_reg[28]_0 ;
  input \tr_reg[21]_0 ;
  input \tr_reg[19]_0 ;
  input \tr_reg[27]_1 ;
  input [4:0]bbus_0;
  input \iv[13]_i_17 ;
  input \iv[13]_i_17_0 ;
  input \iv[7]_i_7 ;
  input \iv[7]_i_7_0 ;
  input \iv[7]_i_7_1 ;
  input \tr_reg[1] ;
  input \tr_reg[1]_0 ;
  input \sr_reg[4]_2 ;
  input \sr_reg[4]_3 ;
  input \sr[4]_i_5 ;
  input \sr[4]_i_5_0 ;
  input \sr[4]_i_16 ;
  input \sr[4]_i_89 ;
  input \sr[4]_i_5_1 ;
  input \sr[4]_i_21_0 ;
  input \sr[4]_i_21_1 ;
  input \tr[19]_i_3 ;
  input \sr[4]_i_5_2 ;
  input \sr[4]_i_20 ;
  input \sr[4]_i_20_0 ;
  input \iv[13]_i_2 ;
  input \sr[4]_i_20_1 ;
  input \sr[4]_i_20_2 ;
  input \iv[12]_i_2 ;
  input \sr[4]_i_44 ;
  input \iv[0]_i_3 ;
  input \iv[10]_i_2 ;
  input \sr[4]_i_16_0 ;
  input \sr[4]_i_33 ;
  input \sr[4]_i_39 ;
  input \iv[8]_i_2 ;
  input \sr[4]_i_40 ;
  input \tr[22]_i_3 ;
  input \tr[24]_i_2 ;
  input \tr[24]_i_3 ;
  input \tr[23]_i_2 ;
  input \tr[17]_i_2 ;
  input \tr[21]_i_2 ;
  input \tr[22]_i_2 ;
  input \tr[20]_i_2 ;
  input \tr[18]_i_2 ;
  input \tr[28]_i_2 ;
  input \tr[25]_i_2 ;
  input \tr[19]_i_2 ;
  input \iv[15]_i_8 ;
  input \iv[15]_i_8_0 ;
  input \iv[15]_i_8_1 ;
  input \tr[19]_i_3_0 ;
  input \sr_reg[6]_11 ;
  input \sr[4]_i_36 ;
  input \sr[5]_i_3 ;
  input \tr[30]_i_3 ;
  input \tr[30]_i_3_0 ;
  input \tr[26]_i_3 ;
  input \tr[29]_i_3 ;
  input \sr[4]_i_42 ;
  input \sr[4]_i_43 ;
  input \iv[0]_i_3_0 ;
  input \iv[5]_i_3 ;
  input \iv[4]_i_3 ;
  input \sr[4]_i_39_0 ;
  input \sr[4]_i_40_0 ;
  input \sr[4]_i_37 ;
  input \sr[6]_i_4 ;
  input \iv[0]_i_3_1 ;
  input \iv[0]_i_10 ;
  input \iv[15]_i_8_2 ;
  input \iv[1]_i_10 ;
  input \iv[1]_i_10_0 ;
  input \iv[1]_i_10_1 ;
  input \iv[3]_i_10 ;
  input \iv[3]_i_10_0 ;
  input \iv[3]_i_10_1 ;
  input \sr[4]_i_45 ;
  input \sr[4]_i_44_0 ;
  input \sr[4]_i_35 ;
  input \iv[6]_i_10 ;
  input \iv[6]_i_10_0 ;
  input \iv[6]_i_10_1 ;
  input \iv[0]_i_10_0 ;
  input \sr[6]_i_12 ;
  input \sr[6]_i_12_0 ;
  input \tr[16]_i_6 ;
  input \tr[16]_i_6_0 ;
  input \iv[7]_i_9 ;
  input \sr[4]_i_43_0 ;
  input \iv[1]_i_9 ;
  input \iv[2]_i_9 ;
  input \iv[3]_i_9 ;
  input \sr[4]_i_45_0 ;
  input \sr[4]_i_44_1 ;
  input \iv[10]_i_5 ;
  input \iv[5]_i_9 ;
  input \iv[4]_i_9 ;
  input \iv[8]_i_5 ;
  input \iv[14]_i_5 ;
  input \iv[9]_i_5 ;
  input \sr[4]_i_38 ;
  input \tr[21]_i_3 ;
  input \tr[20]_i_3 ;
  input \tr[24]_i_3_0 ;
  input \iv[0]_i_10_1 ;
  input \sr[4]_i_87 ;
  input \sr[6]_i_11 ;
  input \sr[4]_i_41 ;
  input \iv[0]_i_19 ;
  input \iv[7]_i_3 ;
  input \sr[4]_i_61 ;
  input \sr[4]_i_139 ;
  input \mul_b_reg[5] ;
  input \mul_b_reg[5]_0 ;
  input \iv[0]_i_7 ;
  input \iv[15]_i_96 ;
  input \iv[15]_i_96_0 ;
  input \mul_b_reg[0] ;
  input \mul_b_reg[0]_0 ;
  input mul_rslt;
  input [32:0]mul_a;
  input \niho_dsp_b[5] ;
  input \mul_a_reg[15] ;
  input \tr[22]_i_11 ;
  input \remden_reg[26] ;
  input \remden_reg[29] ;
  input \remden_reg[25] ;
  input \remden_reg[24] ;
  input \remden_reg[23] ;
  input \remden_reg[22] ;
  input \remden_reg[21] ;
  input \remden_reg[20] ;
  input \remden_reg[18] ;
  input \remden_reg[17] ;
  input \remden_reg[16] ;
  input [5:0]Q;
  input \tr[19]_i_2_0 ;
  input [5:0]\tr[29]_i_2 ;
  input \tr[19]_i_2_1 ;
  input \sr[4]_i_3 ;
  input \iv[0]_i_6 ;
  input [2:0]\iv[0]_i_6_0 ;
  input [2:0]\iv[4]_i_6 ;
  input [3:0]\iv[8]_i_8 ;
  input [3:0]S;
  input irq;
  input [1:0]irq_lev;
  input [5:0]\badr[31]_INST_0_i_69 ;
  input \stat_reg[1] ;
  input [1:0]\stat[0]_i_6 ;
  input \sr[4]_i_19 ;
  input \sr[4]_i_18 ;
  input \grn_reg[0] ;
  input \grn_reg[0]_0 ;
  input [7:0]bbus_sel_0;
  input [7:0]abus_sel_0;
  input \mul_a_reg[32] ;
  input \remden_reg[19] ;
  input \sr[5]_i_2 ;
  input \tr_reg[31]_i_13 ;
  input \remden_reg[30] ;
  input \tr_reg[31]_i_13_0 ;
  input \tr_reg[31]_i_13_1 ;
  input \remden_reg[28] ;
  input \tr_reg[31]_i_32 ;
  input \remden_reg[27] ;
  input \tr_reg[31]_i_32_0 ;
  input \remden_reg[26]_0 ;
  input \tr_reg[31]_i_32_1 ;
  input \tr_reg[31]_i_32_2 ;
  input \tr_reg[23]_i_11 ;
  input \tr_reg[23]_i_11_0 ;
  input \tr_reg[23]_i_11_1 ;
  input \tr_reg[23]_i_11_2 ;
  input \sr_reg[6]_i_6 ;
  input \sr_reg[6]_i_6_0 ;
  input \sr_reg[6]_i_6_1 ;
  input \niho_dsp_b[5]_0 ;
  input \i_/bdatw[15]_INST_0_i_65 ;
  input [1:0]ctl_selb_rn;
  input \i_/bdatw[15]_INST_0_i_65_0 ;
  input \i_/bdatw[15]_INST_0_i_65_1 ;
  input [0:0]ctl_selb_0;
  input \i_/bdatw[15]_INST_0_i_65_2 ;
  input \i_/bdatw[15]_INST_0_i_67 ;
  input \i_/bdatw[15]_INST_0_i_27 ;
  input \i_/bdatw[15]_INST_0_i_67_0 ;
  input \i_/bdatw[15]_INST_0_i_27_0 ;
  input clk;
  input \sr_reg[11]_0 ;
  input \sr_reg[10]_0 ;
  input \sr_reg[8]_169 ;
  input \sr_reg[7]_4 ;
  input \sr_reg[6]_12 ;
  input \sr_reg[5]_2 ;
  input \sr_reg[4]_4 ;
  input \sr_reg[3]_0 ;
  input \sr_reg[2]_0 ;
  input \sr_reg[1]_0 ;
  input \sr_reg[0] ;
  input [31:0]\sp_reg[31]_1 ;
  input \mul_a_reg[14] ;
  input \mul_a_reg[13] ;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input \mul_a_reg[4] ;
  input \mul_a_reg[3] ;
  input \mul_a_reg[2] ;
  input \mul_a_reg[1] ;
  input \mul_a_reg[0] ;
  input \mul_a_reg[32]_0 ;
  input \mul_a_reg[30] ;
  input \mul_a_reg[29] ;
  input \mul_a_reg[28] ;
  input \mul_a_reg[27] ;
  input \mul_a_reg[26] ;
  input \mul_a_reg[25] ;
  input \mul_a_reg[24] ;
  input \mul_a_reg[23] ;
  input \mul_a_reg[22] ;
  input \mul_a_reg[21] ;
  input \mul_a_reg[20] ;
  input \mul_a_reg[19] ;
  input \mul_a_reg[18] ;
  input \mul_a_reg[17] ;
  input \mul_a_reg[16] ;
  input [5:0]bbus_sel_cr;
  input [1:0]bbus_sr;
  input [0:0]E;
  input [31:0]cbus;
  input [0:0]\grn_reg[15] ;
  input [0:0]\grn_reg[15]_0 ;
  input [0:0]\grn_reg[15]_1 ;
  input [0:0]\grn_reg[15]_2 ;
  input [0:0]\grn_reg[15]_3 ;
  input [0:0]\grn_reg[15]_4 ;
  input [15:0]\grn_reg[15]_5 ;
  input [0:0]\grn_reg[15]_6 ;
  input [0:0]\grn_reg[15]_7 ;
  input [0:0]\grn_reg[15]_8 ;
  input [0:0]\grn_reg[15]_9 ;
  input [0:0]\grn_reg[15]_10 ;
  input [0:0]\grn_reg[15]_11 ;
  input [0:0]\grn_reg[15]_12 ;
  input [0:0]\grn_reg[15]_13 ;
  input [0:0]\grn_reg[15]_14 ;
  input [0:0]\grn_reg[15]_15 ;
  input [0:0]\grn_reg[15]_16 ;
  input [0:0]\grn_reg[15]_17 ;
  input [0:0]\grn_reg[15]_18 ;
  input [0:0]\grn_reg[15]_19 ;
  input [0:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
  input [0:0]\grn_reg[15]_22 ;
  input [15:0]\pc_reg[15] ;
  input [1:0]\tr_reg[0] ;
  output irq_lev_0_sn_1;
  output irq_lev_1_sn_1;
  input abus_o_16_sn_1;
  input niho_dsp_b_0_sn_1;

  wire [1:0]D;
  wire [0:0]E;
  wire [0:0]O;
  wire [5:0]Q;
  wire [3:0]S;
  wire [31:0]abus_0;
  wire [31:0]abus_o;
  wire abus_o_16_sn_1;
  wire abus_out_n_4;
  wire abus_out_n_5;
  wire [7:0]abus_sel_0;
  wire [3:0]abus_sel_cr;
  wire [31:16]abus_sp;
  wire [0:0]alu_sr_flag;
  wire [3:0]\art/add/iv[7]_i_32 ;
  wire [3:0]\art/add/sr[5]_i_14 ;
  wire [3:0]\art/add/sr[5]_i_18 ;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[0]_INST_0_i_1_0 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1 ;
  wire [5:0]\badr[31]_INST_0_i_69 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1_0 ;
  wire \badr[6]_INST_0_i_1 ;
  wire bank02_n_0;
  wire bank02_n_1;
  wire bank02_n_10;
  wire bank02_n_100;
  wire bank02_n_101;
  wire bank02_n_102;
  wire bank02_n_103;
  wire bank02_n_104;
  wire bank02_n_105;
  wire bank02_n_106;
  wire bank02_n_107;
  wire bank02_n_108;
  wire bank02_n_109;
  wire bank02_n_11;
  wire bank02_n_110;
  wire bank02_n_111;
  wire bank02_n_112;
  wire bank02_n_113;
  wire bank02_n_114;
  wire bank02_n_115;
  wire bank02_n_116;
  wire bank02_n_117;
  wire bank02_n_118;
  wire bank02_n_119;
  wire bank02_n_12;
  wire bank02_n_120;
  wire bank02_n_121;
  wire bank02_n_122;
  wire bank02_n_123;
  wire bank02_n_124;
  wire bank02_n_125;
  wire bank02_n_126;
  wire bank02_n_127;
  wire bank02_n_13;
  wire bank02_n_14;
  wire bank02_n_140;
  wire bank02_n_144;
  wire bank02_n_15;
  wire bank02_n_150;
  wire bank02_n_16;
  wire bank02_n_17;
  wire bank02_n_177;
  wire bank02_n_178;
  wire bank02_n_18;
  wire bank02_n_181;
  wire bank02_n_182;
  wire bank02_n_183;
  wire bank02_n_186;
  wire bank02_n_187;
  wire bank02_n_189;
  wire bank02_n_19;
  wire bank02_n_190;
  wire bank02_n_191;
  wire bank02_n_196;
  wire bank02_n_197;
  wire bank02_n_198;
  wire bank02_n_2;
  wire bank02_n_20;
  wire bank02_n_200;
  wire bank02_n_202;
  wire bank02_n_203;
  wire bank02_n_204;
  wire bank02_n_206;
  wire bank02_n_207;
  wire bank02_n_21;
  wire bank02_n_214;
  wire bank02_n_216;
  wire bank02_n_217;
  wire bank02_n_218;
  wire bank02_n_22;
  wire bank02_n_23;
  wire bank02_n_231;
  wire bank02_n_234;
  wire bank02_n_235;
  wire bank02_n_24;
  wire bank02_n_243;
  wire bank02_n_245;
  wire bank02_n_247;
  wire bank02_n_25;
  wire bank02_n_251;
  wire bank02_n_252;
  wire bank02_n_253;
  wire bank02_n_259;
  wire bank02_n_26;
  wire bank02_n_260;
  wire bank02_n_261;
  wire bank02_n_264;
  wire bank02_n_265;
  wire bank02_n_266;
  wire bank02_n_267;
  wire bank02_n_27;
  wire bank02_n_272;
  wire bank02_n_274;
  wire bank02_n_279;
  wire bank02_n_28;
  wire bank02_n_280;
  wire bank02_n_282;
  wire bank02_n_283;
  wire bank02_n_284;
  wire bank02_n_286;
  wire bank02_n_289;
  wire bank02_n_29;
  wire bank02_n_291;
  wire bank02_n_295;
  wire bank02_n_298;
  wire bank02_n_3;
  wire bank02_n_30;
  wire bank02_n_300;
  wire bank02_n_301;
  wire bank02_n_304;
  wire bank02_n_31;
  wire bank02_n_32;
  wire bank02_n_33;
  wire bank02_n_34;
  wire bank02_n_347;
  wire bank02_n_35;
  wire bank02_n_36;
  wire bank02_n_364;
  wire bank02_n_37;
  wire bank02_n_38;
  wire bank02_n_385;
  wire bank02_n_387;
  wire bank02_n_388;
  wire bank02_n_39;
  wire bank02_n_390;
  wire bank02_n_4;
  wire bank02_n_40;
  wire bank02_n_41;
  wire bank02_n_415;
  wire bank02_n_416;
  wire bank02_n_417;
  wire bank02_n_418;
  wire bank02_n_419;
  wire bank02_n_42;
  wire bank02_n_420;
  wire bank02_n_421;
  wire bank02_n_422;
  wire bank02_n_423;
  wire bank02_n_424;
  wire bank02_n_425;
  wire bank02_n_426;
  wire bank02_n_427;
  wire bank02_n_428;
  wire bank02_n_429;
  wire bank02_n_43;
  wire bank02_n_430;
  wire bank02_n_431;
  wire bank02_n_432;
  wire bank02_n_433;
  wire bank02_n_434;
  wire bank02_n_435;
  wire bank02_n_436;
  wire bank02_n_437;
  wire bank02_n_438;
  wire bank02_n_439;
  wire bank02_n_44;
  wire bank02_n_440;
  wire bank02_n_441;
  wire bank02_n_442;
  wire bank02_n_443;
  wire bank02_n_444;
  wire bank02_n_445;
  wire bank02_n_446;
  wire bank02_n_447;
  wire bank02_n_448;
  wire bank02_n_449;
  wire bank02_n_45;
  wire bank02_n_450;
  wire bank02_n_451;
  wire bank02_n_452;
  wire bank02_n_453;
  wire bank02_n_454;
  wire bank02_n_455;
  wire bank02_n_456;
  wire bank02_n_457;
  wire bank02_n_458;
  wire bank02_n_459;
  wire bank02_n_46;
  wire bank02_n_460;
  wire bank02_n_461;
  wire bank02_n_462;
  wire bank02_n_463;
  wire bank02_n_464;
  wire bank02_n_465;
  wire bank02_n_466;
  wire bank02_n_467;
  wire bank02_n_468;
  wire bank02_n_469;
  wire bank02_n_47;
  wire bank02_n_470;
  wire bank02_n_471;
  wire bank02_n_472;
  wire bank02_n_473;
  wire bank02_n_474;
  wire bank02_n_475;
  wire bank02_n_476;
  wire bank02_n_477;
  wire bank02_n_478;
  wire bank02_n_479;
  wire bank02_n_48;
  wire bank02_n_480;
  wire bank02_n_481;
  wire bank02_n_482;
  wire bank02_n_483;
  wire bank02_n_484;
  wire bank02_n_485;
  wire bank02_n_486;
  wire bank02_n_487;
  wire bank02_n_488;
  wire bank02_n_489;
  wire bank02_n_49;
  wire bank02_n_490;
  wire bank02_n_5;
  wire bank02_n_50;
  wire bank02_n_51;
  wire bank02_n_52;
  wire bank02_n_53;
  wire bank02_n_54;
  wire bank02_n_55;
  wire bank02_n_56;
  wire bank02_n_57;
  wire bank02_n_58;
  wire bank02_n_59;
  wire bank02_n_6;
  wire bank02_n_60;
  wire bank02_n_61;
  wire bank02_n_62;
  wire bank02_n_63;
  wire bank02_n_64;
  wire bank02_n_65;
  wire bank02_n_66;
  wire bank02_n_67;
  wire bank02_n_68;
  wire bank02_n_69;
  wire bank02_n_7;
  wire bank02_n_70;
  wire bank02_n_71;
  wire bank02_n_72;
  wire bank02_n_73;
  wire bank02_n_74;
  wire bank02_n_75;
  wire bank02_n_76;
  wire bank02_n_77;
  wire bank02_n_78;
  wire bank02_n_79;
  wire bank02_n_8;
  wire bank02_n_80;
  wire bank02_n_81;
  wire bank02_n_82;
  wire bank02_n_83;
  wire bank02_n_84;
  wire bank02_n_85;
  wire bank02_n_86;
  wire bank02_n_87;
  wire bank02_n_88;
  wire bank02_n_89;
  wire bank02_n_9;
  wire bank02_n_90;
  wire bank02_n_91;
  wire bank02_n_92;
  wire bank02_n_93;
  wire bank02_n_94;
  wire bank02_n_95;
  wire bank02_n_96;
  wire bank02_n_97;
  wire bank02_n_98;
  wire bank02_n_99;
  wire bank13_n_0;
  wire bank13_n_1;
  wire bank13_n_10;
  wire bank13_n_100;
  wire bank13_n_101;
  wire bank13_n_102;
  wire bank13_n_103;
  wire bank13_n_104;
  wire bank13_n_105;
  wire bank13_n_106;
  wire bank13_n_107;
  wire bank13_n_108;
  wire bank13_n_109;
  wire bank13_n_11;
  wire bank13_n_110;
  wire bank13_n_111;
  wire bank13_n_112;
  wire bank13_n_113;
  wire bank13_n_114;
  wire bank13_n_115;
  wire bank13_n_116;
  wire bank13_n_117;
  wire bank13_n_118;
  wire bank13_n_119;
  wire bank13_n_12;
  wire bank13_n_120;
  wire bank13_n_121;
  wire bank13_n_122;
  wire bank13_n_123;
  wire bank13_n_124;
  wire bank13_n_125;
  wire bank13_n_126;
  wire bank13_n_127;
  wire bank13_n_128;
  wire bank13_n_129;
  wire bank13_n_13;
  wire bank13_n_130;
  wire bank13_n_131;
  wire bank13_n_132;
  wire bank13_n_133;
  wire bank13_n_134;
  wire bank13_n_135;
  wire bank13_n_136;
  wire bank13_n_137;
  wire bank13_n_138;
  wire bank13_n_139;
  wire bank13_n_14;
  wire bank13_n_140;
  wire bank13_n_141;
  wire bank13_n_142;
  wire bank13_n_143;
  wire bank13_n_144;
  wire bank13_n_145;
  wire bank13_n_146;
  wire bank13_n_147;
  wire bank13_n_148;
  wire bank13_n_149;
  wire bank13_n_15;
  wire bank13_n_150;
  wire bank13_n_151;
  wire bank13_n_152;
  wire bank13_n_153;
  wire bank13_n_154;
  wire bank13_n_155;
  wire bank13_n_156;
  wire bank13_n_157;
  wire bank13_n_158;
  wire bank13_n_159;
  wire bank13_n_16;
  wire bank13_n_160;
  wire bank13_n_161;
  wire bank13_n_162;
  wire bank13_n_163;
  wire bank13_n_164;
  wire bank13_n_165;
  wire bank13_n_166;
  wire bank13_n_167;
  wire bank13_n_168;
  wire bank13_n_169;
  wire bank13_n_17;
  wire bank13_n_170;
  wire bank13_n_171;
  wire bank13_n_172;
  wire bank13_n_173;
  wire bank13_n_174;
  wire bank13_n_175;
  wire bank13_n_176;
  wire bank13_n_177;
  wire bank13_n_178;
  wire bank13_n_179;
  wire bank13_n_18;
  wire bank13_n_180;
  wire bank13_n_181;
  wire bank13_n_182;
  wire bank13_n_183;
  wire bank13_n_184;
  wire bank13_n_185;
  wire bank13_n_186;
  wire bank13_n_187;
  wire bank13_n_188;
  wire bank13_n_189;
  wire bank13_n_19;
  wire bank13_n_190;
  wire bank13_n_191;
  wire bank13_n_192;
  wire bank13_n_193;
  wire bank13_n_194;
  wire bank13_n_195;
  wire bank13_n_196;
  wire bank13_n_197;
  wire bank13_n_198;
  wire bank13_n_199;
  wire bank13_n_2;
  wire bank13_n_20;
  wire bank13_n_200;
  wire bank13_n_201;
  wire bank13_n_202;
  wire bank13_n_203;
  wire bank13_n_204;
  wire bank13_n_205;
  wire bank13_n_206;
  wire bank13_n_207;
  wire bank13_n_208;
  wire bank13_n_209;
  wire bank13_n_21;
  wire bank13_n_210;
  wire bank13_n_211;
  wire bank13_n_212;
  wire bank13_n_213;
  wire bank13_n_214;
  wire bank13_n_215;
  wire bank13_n_216;
  wire bank13_n_217;
  wire bank13_n_218;
  wire bank13_n_219;
  wire bank13_n_22;
  wire bank13_n_220;
  wire bank13_n_221;
  wire bank13_n_222;
  wire bank13_n_223;
  wire bank13_n_224;
  wire bank13_n_225;
  wire bank13_n_226;
  wire bank13_n_227;
  wire bank13_n_228;
  wire bank13_n_229;
  wire bank13_n_23;
  wire bank13_n_230;
  wire bank13_n_231;
  wire bank13_n_232;
  wire bank13_n_233;
  wire bank13_n_234;
  wire bank13_n_235;
  wire bank13_n_236;
  wire bank13_n_24;
  wire bank13_n_25;
  wire bank13_n_26;
  wire bank13_n_27;
  wire bank13_n_28;
  wire bank13_n_29;
  wire bank13_n_3;
  wire bank13_n_30;
  wire bank13_n_31;
  wire bank13_n_32;
  wire bank13_n_33;
  wire bank13_n_34;
  wire bank13_n_35;
  wire bank13_n_36;
  wire bank13_n_37;
  wire bank13_n_38;
  wire bank13_n_39;
  wire bank13_n_4;
  wire bank13_n_40;
  wire bank13_n_41;
  wire bank13_n_42;
  wire bank13_n_43;
  wire bank13_n_44;
  wire bank13_n_45;
  wire bank13_n_46;
  wire bank13_n_47;
  wire bank13_n_48;
  wire bank13_n_49;
  wire bank13_n_5;
  wire bank13_n_50;
  wire bank13_n_51;
  wire bank13_n_52;
  wire bank13_n_53;
  wire bank13_n_54;
  wire bank13_n_55;
  wire bank13_n_56;
  wire bank13_n_57;
  wire bank13_n_58;
  wire bank13_n_59;
  wire bank13_n_6;
  wire bank13_n_60;
  wire bank13_n_61;
  wire bank13_n_62;
  wire bank13_n_63;
  wire bank13_n_65;
  wire bank13_n_66;
  wire bank13_n_67;
  wire bank13_n_68;
  wire bank13_n_69;
  wire bank13_n_7;
  wire bank13_n_70;
  wire bank13_n_71;
  wire bank13_n_72;
  wire bank13_n_73;
  wire bank13_n_74;
  wire bank13_n_75;
  wire bank13_n_76;
  wire bank13_n_77;
  wire bank13_n_78;
  wire bank13_n_79;
  wire bank13_n_8;
  wire bank13_n_80;
  wire bank13_n_81;
  wire bank13_n_82;
  wire bank13_n_83;
  wire bank13_n_84;
  wire bank13_n_85;
  wire bank13_n_86;
  wire bank13_n_87;
  wire bank13_n_88;
  wire bank13_n_89;
  wire bank13_n_9;
  wire bank13_n_90;
  wire bank13_n_91;
  wire bank13_n_92;
  wire bank13_n_93;
  wire bank13_n_94;
  wire bank13_n_95;
  wire bank13_n_96;
  wire bank13_n_97;
  wire bank13_n_98;
  wire bank13_n_99;
  wire [0:0]bank_sel;
  wire [4:0]bbus_0;
  wire [1:0]bbus_o;
  wire bbus_out_n_10;
  wire bbus_out_n_11;
  wire bbus_out_n_16;
  wire bbus_out_n_17;
  wire bbus_out_n_28;
  wire bbus_out_n_29;
  wire bbus_out_n_30;
  wire bbus_out_n_35;
  wire [7:0]bbus_sel_0;
  wire [5:0]bbus_sel_cr;
  wire [1:0]bbus_sr;
  wire \bdatw[8]_INST_0_i_2 ;
  wire [31:0]cbus;
  wire [0:0]cbus_sel_0;
  wire clk;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire ctl_sp_dec;
  wire ctl_sp_id4;
  wire ctl_sp_inc;
  wire fch_irq_req;
  wire [15:0]fch_pc;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [0:0]\grn_reg[15] ;
  wire [0:0]\grn_reg[15]_0 ;
  wire [0:0]\grn_reg[15]_1 ;
  wire [0:0]\grn_reg[15]_10 ;
  wire [0:0]\grn_reg[15]_11 ;
  wire [0:0]\grn_reg[15]_12 ;
  wire [0:0]\grn_reg[15]_13 ;
  wire [0:0]\grn_reg[15]_14 ;
  wire [0:0]\grn_reg[15]_15 ;
  wire [0:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [0:0]\grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [0:0]\grn_reg[15]_2 ;
  wire [0:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [0:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_3 ;
  wire [0:0]\grn_reg[15]_4 ;
  wire [15:0]\grn_reg[15]_5 ;
  wire [0:0]\grn_reg[15]_6 ;
  wire [0:0]\grn_reg[15]_7 ;
  wire [0:0]\grn_reg[15]_8 ;
  wire [0:0]\grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \i_/bdatw[15]_INST_0_i_27 ;
  wire \i_/bdatw[15]_INST_0_i_27_0 ;
  wire \i_/bdatw[15]_INST_0_i_65 ;
  wire \i_/bdatw[15]_INST_0_i_65_0 ;
  wire \i_/bdatw[15]_INST_0_i_65_1 ;
  wire \i_/bdatw[15]_INST_0_i_65_2 ;
  wire \i_/bdatw[15]_INST_0_i_67 ;
  wire \i_/bdatw[15]_INST_0_i_67_0 ;
  wire irq;
  wire [1:0]irq_lev;
  wire irq_lev_0_sn_1;
  wire irq_lev_1_sn_1;
  wire \iv[0]_i_10 ;
  wire \iv[0]_i_10_0 ;
  wire \iv[0]_i_10_1 ;
  wire \iv[0]_i_19 ;
  wire \iv[0]_i_25 ;
  wire \iv[0]_i_3 ;
  wire \iv[0]_i_3_0 ;
  wire \iv[0]_i_3_1 ;
  wire \iv[0]_i_6 ;
  wire [2:0]\iv[0]_i_6_0 ;
  wire \iv[0]_i_7 ;
  wire \iv[10]_i_10 ;
  wire \iv[10]_i_2 ;
  wire \iv[10]_i_5 ;
  wire \iv[10]_i_9 ;
  wire \iv[11]_i_11 ;
  wire \iv[12]_i_2 ;
  wire \iv[13]_i_10 ;
  wire \iv[13]_i_17 ;
  wire \iv[13]_i_17_0 ;
  wire \iv[13]_i_2 ;
  wire \iv[13]_i_27 ;
  wire \iv[14]_i_11 ;
  wire \iv[14]_i_35 ;
  wire \iv[14]_i_49 ;
  wire \iv[14]_i_5 ;
  wire \iv[15]_i_108 ;
  wire \iv[15]_i_108_0 ;
  wire \iv[15]_i_108_1 ;
  wire \iv[15]_i_108_10 ;
  wire \iv[15]_i_108_11 ;
  wire \iv[15]_i_108_12 ;
  wire \iv[15]_i_108_13 ;
  wire \iv[15]_i_108_14 ;
  wire \iv[15]_i_108_15 ;
  wire \iv[15]_i_108_16 ;
  wire \iv[15]_i_108_17 ;
  wire \iv[15]_i_108_18 ;
  wire \iv[15]_i_108_19 ;
  wire \iv[15]_i_108_2 ;
  wire \iv[15]_i_108_20 ;
  wire \iv[15]_i_108_21 ;
  wire \iv[15]_i_108_22 ;
  wire \iv[15]_i_108_23 ;
  wire \iv[15]_i_108_3 ;
  wire \iv[15]_i_108_4 ;
  wire \iv[15]_i_108_5 ;
  wire \iv[15]_i_108_6 ;
  wire \iv[15]_i_108_7 ;
  wire \iv[15]_i_108_8 ;
  wire \iv[15]_i_108_9 ;
  wire \iv[15]_i_8 ;
  wire \iv[15]_i_8_0 ;
  wire \iv[15]_i_8_1 ;
  wire \iv[15]_i_8_2 ;
  wire \iv[15]_i_96 ;
  wire \iv[15]_i_96_0 ;
  wire \iv[1]_i_10 ;
  wire \iv[1]_i_10_0 ;
  wire \iv[1]_i_10_1 ;
  wire \iv[1]_i_9 ;
  wire \iv[2]_i_9 ;
  wire \iv[3]_i_10 ;
  wire \iv[3]_i_10_0 ;
  wire \iv[3]_i_10_1 ;
  wire \iv[3]_i_9 ;
  wire \iv[4]_i_3 ;
  wire \iv[4]_i_35 ;
  wire [2:0]\iv[4]_i_6 ;
  wire \iv[4]_i_9 ;
  wire \iv[5]_i_3 ;
  wire \iv[5]_i_9 ;
  wire \iv[6]_i_10 ;
  wire \iv[6]_i_10_0 ;
  wire \iv[6]_i_10_1 ;
  wire \iv[7]_i_17 ;
  wire \iv[7]_i_25 ;
  wire \iv[7]_i_3 ;
  wire \iv[7]_i_33 ;
  wire \iv[7]_i_7 ;
  wire \iv[7]_i_7_0 ;
  wire \iv[7]_i_7_1 ;
  wire \iv[7]_i_9 ;
  wire \iv[8]_i_2 ;
  wire \iv[8]_i_20 ;
  wire \iv[8]_i_34 ;
  wire \iv[8]_i_5 ;
  wire [3:0]\iv[8]_i_8 ;
  wire \iv[9]_i_11 ;
  wire \iv[9]_i_5 ;
  wire \iv_reg[10] ;
  wire \iv_reg[11] ;
  wire \iv_reg[12] ;
  wire \iv_reg[13] ;
  wire \iv_reg[14] ;
  wire \iv_reg[15] ;
  wire [15:0]\iv_reg[15]_0 ;
  wire \iv_reg[6] ;
  wire \iv_reg[7] ;
  wire \iv_reg[8] ;
  wire \iv_reg[9] ;
  wire [32:0]mul_a;
  wire [13:0]mul_a_i;
  wire \mul_a_reg[0] ;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[13] ;
  wire \mul_a_reg[14] ;
  wire \mul_a_reg[15] ;
  wire \mul_a_reg[16] ;
  wire \mul_a_reg[17] ;
  wire \mul_a_reg[18] ;
  wire \mul_a_reg[19] ;
  wire \mul_a_reg[1] ;
  wire \mul_a_reg[20] ;
  wire \mul_a_reg[21] ;
  wire \mul_a_reg[22] ;
  wire \mul_a_reg[23] ;
  wire \mul_a_reg[24] ;
  wire \mul_a_reg[25] ;
  wire \mul_a_reg[26] ;
  wire \mul_a_reg[27] ;
  wire \mul_a_reg[28] ;
  wire \mul_a_reg[29] ;
  wire \mul_a_reg[2] ;
  wire \mul_a_reg[30] ;
  wire \mul_a_reg[32] ;
  wire \mul_a_reg[32]_0 ;
  wire \mul_a_reg[3] ;
  wire \mul_a_reg[4] ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[9] ;
  wire \mul_b_reg[0] ;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[5] ;
  wire \mul_b_reg[5]_0 ;
  wire mul_rslt;
  wire mul_rslt0;
  wire [32:0]niho_dsp_a;
  wire \niho_dsp_a[15]_INST_0_i_3 ;
  wire [1:0]niho_dsp_b;
  wire \niho_dsp_b[5] ;
  wire \niho_dsp_b[5]_0 ;
  wire niho_dsp_b_0_sn_1;
  wire [5:0]niho_dsp_c;
  wire [12:0]out;
  wire p_0_in;
  wire [15:0]p_0_in_0;
  wire [31:1]p_0_in_1;
  wire [15:9]p_0_in_2;
  wire [15:0]p_1_in;
  wire [6:0]p_2_in;
  wire [15:0]\pc_reg[15] ;
  wire \remden_reg[16] ;
  wire \remden_reg[17] ;
  wire \remden_reg[18] ;
  wire \remden_reg[19] ;
  wire \remden_reg[20] ;
  wire \remden_reg[21] ;
  wire \remden_reg[22] ;
  wire \remden_reg[23] ;
  wire \remden_reg[24] ;
  wire \remden_reg[25] ;
  wire \remden_reg[26] ;
  wire \remden_reg[26]_0 ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire [15:0]rgf_pc;
  wire rst_n;
  wire [31:1]sp_dec_0;
  wire [0:0]\sp_reg[0] ;
  wire \sp_reg[10] ;
  wire \sp_reg[11] ;
  wire \sp_reg[12] ;
  wire \sp_reg[13] ;
  wire \sp_reg[14] ;
  wire \sp_reg[15] ;
  wire \sp_reg[16] ;
  wire \sp_reg[16]_0 ;
  wire \sp_reg[17] ;
  wire \sp_reg[17]_0 ;
  wire \sp_reg[18] ;
  wire \sp_reg[18]_0 ;
  wire \sp_reg[19] ;
  wire \sp_reg[19]_0 ;
  wire \sp_reg[1] ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[20] ;
  wire \sp_reg[20]_0 ;
  wire \sp_reg[21] ;
  wire \sp_reg[21]_0 ;
  wire \sp_reg[22] ;
  wire \sp_reg[22]_0 ;
  wire \sp_reg[23] ;
  wire \sp_reg[23]_0 ;
  wire \sp_reg[24] ;
  wire \sp_reg[24]_0 ;
  wire \sp_reg[25] ;
  wire \sp_reg[25]_0 ;
  wire \sp_reg[26] ;
  wire \sp_reg[26]_0 ;
  wire \sp_reg[27] ;
  wire \sp_reg[27]_0 ;
  wire \sp_reg[28] ;
  wire \sp_reg[28]_0 ;
  wire \sp_reg[29] ;
  wire \sp_reg[29]_0 ;
  wire \sp_reg[2] ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[30] ;
  wire \sp_reg[30]_0 ;
  wire \sp_reg[31] ;
  wire \sp_reg[31]_0 ;
  wire [31:0]\sp_reg[31]_1 ;
  wire \sp_reg[3] ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[4] ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[5] ;
  wire \sp_reg[6] ;
  wire \sp_reg[7] ;
  wire \sp_reg[8] ;
  wire \sp_reg[9] ;
  wire \sr[4]_i_116 ;
  wire \sr[4]_i_139 ;
  wire \sr[4]_i_147 ;
  wire \sr[4]_i_16 ;
  wire \sr[4]_i_16_0 ;
  wire \sr[4]_i_18 ;
  wire \sr[4]_i_19 ;
  wire \sr[4]_i_20 ;
  wire \sr[4]_i_20_0 ;
  wire \sr[4]_i_20_1 ;
  wire \sr[4]_i_20_2 ;
  wire \sr[4]_i_21 ;
  wire \sr[4]_i_21_0 ;
  wire \sr[4]_i_21_1 ;
  wire \sr[4]_i_3 ;
  wire \sr[4]_i_33 ;
  wire \sr[4]_i_35 ;
  wire \sr[4]_i_36 ;
  wire \sr[4]_i_37 ;
  wire \sr[4]_i_38 ;
  wire \sr[4]_i_39 ;
  wire \sr[4]_i_39_0 ;
  wire \sr[4]_i_40 ;
  wire \sr[4]_i_40_0 ;
  wire \sr[4]_i_41 ;
  wire \sr[4]_i_42 ;
  wire \sr[4]_i_43 ;
  wire \sr[4]_i_43_0 ;
  wire \sr[4]_i_44 ;
  wire \sr[4]_i_44_0 ;
  wire \sr[4]_i_44_1 ;
  wire \sr[4]_i_45 ;
  wire \sr[4]_i_45_0 ;
  wire \sr[4]_i_5 ;
  wire \sr[4]_i_5_0 ;
  wire \sr[4]_i_5_1 ;
  wire \sr[4]_i_5_2 ;
  wire \sr[4]_i_61 ;
  wire \sr[4]_i_65 ;
  wire \sr[4]_i_87 ;
  wire \sr[4]_i_89 ;
  wire \sr[5]_i_2 ;
  wire \sr[5]_i_3 ;
  wire \sr[6]_i_11 ;
  wire \sr[6]_i_12 ;
  wire \sr[6]_i_12_0 ;
  wire \sr[6]_i_13 ;
  wire \sr[6]_i_4 ;
  wire \sr_reg[0] ;
  wire \sr_reg[10] ;
  wire \sr_reg[10]_0 ;
  wire \sr_reg[11] ;
  wire \sr_reg[11]_0 ;
  wire \sr_reg[12] ;
  wire \sr_reg[13] ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[15]_0 ;
  wire \sr_reg[1] ;
  wire \sr_reg[1]_0 ;
  wire \sr_reg[2] ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[3] ;
  wire \sr_reg[3]_0 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[4]_3 ;
  wire \sr_reg[4]_4 ;
  wire \sr_reg[5] ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_11 ;
  wire \sr_reg[6]_12 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire [3:0]\sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_7 ;
  wire \sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;
  wire \sr_reg[6]_i_6 ;
  wire \sr_reg[6]_i_6_0 ;
  wire \sr_reg[6]_i_6_1 ;
  wire \sr_reg[7] ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[7]_3 ;
  wire \sr_reg[7]_4 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire [0:0]\sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_100 ;
  wire \sr_reg[8]_101 ;
  wire \sr_reg[8]_102 ;
  wire \sr_reg[8]_103 ;
  wire \sr_reg[8]_104 ;
  wire \sr_reg[8]_105 ;
  wire \sr_reg[8]_106 ;
  wire \sr_reg[8]_107 ;
  wire \sr_reg[8]_108 ;
  wire \sr_reg[8]_109 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_110 ;
  wire \sr_reg[8]_111 ;
  wire \sr_reg[8]_112 ;
  wire \sr_reg[8]_113 ;
  wire \sr_reg[8]_114 ;
  wire \sr_reg[8]_115 ;
  wire \sr_reg[8]_116 ;
  wire \sr_reg[8]_117 ;
  wire \sr_reg[8]_118 ;
  wire \sr_reg[8]_119 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_120 ;
  wire \sr_reg[8]_121 ;
  wire \sr_reg[8]_122 ;
  wire \sr_reg[8]_123 ;
  wire \sr_reg[8]_124 ;
  wire \sr_reg[8]_125 ;
  wire \sr_reg[8]_126 ;
  wire \sr_reg[8]_127 ;
  wire \sr_reg[8]_128 ;
  wire \sr_reg[8]_129 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_130 ;
  wire \sr_reg[8]_131 ;
  wire \sr_reg[8]_132 ;
  wire \sr_reg[8]_133 ;
  wire \sr_reg[8]_134 ;
  wire \sr_reg[8]_135 ;
  wire \sr_reg[8]_136 ;
  wire \sr_reg[8]_137 ;
  wire \sr_reg[8]_138 ;
  wire \sr_reg[8]_139 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_140 ;
  wire \sr_reg[8]_141 ;
  wire \sr_reg[8]_142 ;
  wire \sr_reg[8]_143 ;
  wire \sr_reg[8]_144 ;
  wire \sr_reg[8]_145 ;
  wire \sr_reg[8]_146 ;
  wire \sr_reg[8]_147 ;
  wire \sr_reg[8]_148 ;
  wire \sr_reg[8]_149 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_150 ;
  wire \sr_reg[8]_151 ;
  wire \sr_reg[8]_152 ;
  wire \sr_reg[8]_153 ;
  wire \sr_reg[8]_154 ;
  wire \sr_reg[8]_155 ;
  wire \sr_reg[8]_156 ;
  wire \sr_reg[8]_157 ;
  wire \sr_reg[8]_158 ;
  wire [1:0]\sr_reg[8]_159 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_160 ;
  wire \sr_reg[8]_161 ;
  wire \sr_reg[8]_162 ;
  wire \sr_reg[8]_163 ;
  wire \sr_reg[8]_164 ;
  wire \sr_reg[8]_165 ;
  wire \sr_reg[8]_166 ;
  wire \sr_reg[8]_167 ;
  wire \sr_reg[8]_168 ;
  wire \sr_reg[8]_169 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_51 ;
  wire \sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire \sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire \sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_60 ;
  wire \sr_reg[8]_61 ;
  wire \sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire \sr_reg[8]_71 ;
  wire \sr_reg[8]_72 ;
  wire \sr_reg[8]_73 ;
  wire \sr_reg[8]_74 ;
  wire \sr_reg[8]_75 ;
  wire \sr_reg[8]_76 ;
  wire \sr_reg[8]_77 ;
  wire \sr_reg[8]_78 ;
  wire \sr_reg[8]_79 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_80 ;
  wire \sr_reg[8]_81 ;
  wire \sr_reg[8]_82 ;
  wire \sr_reg[8]_83 ;
  wire \sr_reg[8]_84 ;
  wire \sr_reg[8]_85 ;
  wire \sr_reg[8]_86 ;
  wire \sr_reg[8]_87 ;
  wire \sr_reg[8]_88 ;
  wire \sr_reg[8]_89 ;
  wire \sr_reg[8]_9 ;
  wire \sr_reg[8]_90 ;
  wire \sr_reg[8]_91 ;
  wire \sr_reg[8]_92 ;
  wire \sr_reg[8]_93 ;
  wire \sr_reg[8]_94 ;
  wire \sr_reg[8]_95 ;
  wire \sr_reg[8]_96 ;
  wire \sr_reg[8]_97 ;
  wire \sr_reg[8]_98 ;
  wire \sr_reg[8]_99 ;
  wire \sr_reg[9] ;
  wire sreg_n_101;
  wire sreg_n_102;
  wire sreg_n_103;
  wire sreg_n_107;
  wire sreg_n_108;
  wire sreg_n_109;
  wire sreg_n_110;
  wire sreg_n_113;
  wire sreg_n_116;
  wire sreg_n_117;
  wire sreg_n_118;
  wire sreg_n_119;
  wire sreg_n_120;
  wire sreg_n_122;
  wire sreg_n_123;
  wire sreg_n_124;
  wire sreg_n_125;
  wire sreg_n_126;
  wire sreg_n_127;
  wire sreg_n_128;
  wire sreg_n_129;
  wire sreg_n_130;
  wire sreg_n_131;
  wire sreg_n_132;
  wire sreg_n_133;
  wire sreg_n_134;
  wire sreg_n_135;
  wire sreg_n_136;
  wire sreg_n_137;
  wire sreg_n_138;
  wire sreg_n_140;
  wire sreg_n_142;
  wire sreg_n_143;
  wire sreg_n_144;
  wire sreg_n_145;
  wire sreg_n_146;
  wire sreg_n_147;
  wire sreg_n_148;
  wire sreg_n_149;
  wire sreg_n_150;
  wire sreg_n_151;
  wire sreg_n_152;
  wire sreg_n_153;
  wire sreg_n_154;
  wire sreg_n_156;
  wire sreg_n_157;
  wire sreg_n_16;
  wire sreg_n_17;
  wire sreg_n_18;
  wire sreg_n_19;
  wire sreg_n_218;
  wire sreg_n_219;
  wire sreg_n_220;
  wire sreg_n_221;
  wire sreg_n_222;
  wire sreg_n_223;
  wire sreg_n_24;
  wire sreg_n_26;
  wire sreg_n_261;
  wire sreg_n_262;
  wire sreg_n_263;
  wire sreg_n_264;
  wire sreg_n_265;
  wire sreg_n_266;
  wire sreg_n_267;
  wire sreg_n_268;
  wire sreg_n_269;
  wire sreg_n_270;
  wire sreg_n_274;
  wire sreg_n_275;
  wire sreg_n_276;
  wire sreg_n_28;
  wire sreg_n_280;
  wire sreg_n_281;
  wire sreg_n_282;
  wire sreg_n_283;
  wire sreg_n_284;
  wire sreg_n_285;
  wire sreg_n_286;
  wire sreg_n_287;
  wire sreg_n_288;
  wire sreg_n_289;
  wire sreg_n_29;
  wire sreg_n_290;
  wire sreg_n_291;
  wire sreg_n_292;
  wire sreg_n_293;
  wire sreg_n_294;
  wire sreg_n_295;
  wire sreg_n_296;
  wire sreg_n_297;
  wire sreg_n_298;
  wire sreg_n_299;
  wire sreg_n_30;
  wire sreg_n_300;
  wire sreg_n_301;
  wire sreg_n_302;
  wire sreg_n_303;
  wire sreg_n_304;
  wire sreg_n_305;
  wire sreg_n_306;
  wire sreg_n_307;
  wire sreg_n_308;
  wire sreg_n_309;
  wire sreg_n_31;
  wire sreg_n_310;
  wire sreg_n_311;
  wire sreg_n_312;
  wire sreg_n_313;
  wire sreg_n_314;
  wire sreg_n_315;
  wire sreg_n_316;
  wire sreg_n_317;
  wire sreg_n_318;
  wire sreg_n_319;
  wire sreg_n_32;
  wire sreg_n_320;
  wire sreg_n_321;
  wire sreg_n_322;
  wire sreg_n_323;
  wire sreg_n_324;
  wire sreg_n_325;
  wire sreg_n_326;
  wire sreg_n_327;
  wire sreg_n_328;
  wire sreg_n_329;
  wire sreg_n_33;
  wire sreg_n_330;
  wire sreg_n_331;
  wire sreg_n_332;
  wire sreg_n_333;
  wire sreg_n_334;
  wire sreg_n_335;
  wire sreg_n_336;
  wire sreg_n_337;
  wire sreg_n_338;
  wire sreg_n_339;
  wire sreg_n_340;
  wire sreg_n_341;
  wire sreg_n_342;
  wire sreg_n_343;
  wire sreg_n_344;
  wire sreg_n_345;
  wire sreg_n_346;
  wire sreg_n_347;
  wire sreg_n_348;
  wire sreg_n_349;
  wire sreg_n_350;
  wire sreg_n_351;
  wire sreg_n_352;
  wire sreg_n_353;
  wire sreg_n_354;
  wire sreg_n_355;
  wire sreg_n_356;
  wire sreg_n_357;
  wire sreg_n_358;
  wire sreg_n_359;
  wire sreg_n_36;
  wire sreg_n_360;
  wire sreg_n_361;
  wire sreg_n_362;
  wire sreg_n_363;
  wire sreg_n_364;
  wire sreg_n_365;
  wire sreg_n_366;
  wire sreg_n_367;
  wire sreg_n_368;
  wire sreg_n_369;
  wire sreg_n_370;
  wire sreg_n_371;
  wire sreg_n_372;
  wire sreg_n_373;
  wire sreg_n_374;
  wire sreg_n_375;
  wire sreg_n_376;
  wire sreg_n_377;
  wire sreg_n_378;
  wire sreg_n_379;
  wire sreg_n_380;
  wire sreg_n_381;
  wire sreg_n_382;
  wire sreg_n_383;
  wire sreg_n_384;
  wire sreg_n_385;
  wire sreg_n_386;
  wire sreg_n_387;
  wire sreg_n_388;
  wire sreg_n_389;
  wire sreg_n_390;
  wire sreg_n_391;
  wire sreg_n_392;
  wire sreg_n_393;
  wire sreg_n_394;
  wire sreg_n_395;
  wire sreg_n_396;
  wire sreg_n_397;
  wire sreg_n_398;
  wire sreg_n_399;
  wire sreg_n_400;
  wire sreg_n_401;
  wire sreg_n_402;
  wire sreg_n_403;
  wire sreg_n_404;
  wire sreg_n_405;
  wire sreg_n_406;
  wire sreg_n_407;
  wire sreg_n_408;
  wire sreg_n_409;
  wire sreg_n_410;
  wire sreg_n_411;
  wire sreg_n_412;
  wire sreg_n_413;
  wire sreg_n_414;
  wire sreg_n_415;
  wire sreg_n_416;
  wire sreg_n_417;
  wire sreg_n_418;
  wire sreg_n_419;
  wire sreg_n_420;
  wire sreg_n_421;
  wire sreg_n_422;
  wire sreg_n_423;
  wire sreg_n_424;
  wire sreg_n_425;
  wire sreg_n_426;
  wire sreg_n_427;
  wire sreg_n_428;
  wire sreg_n_429;
  wire sreg_n_43;
  wire sreg_n_430;
  wire sreg_n_431;
  wire sreg_n_432;
  wire sreg_n_433;
  wire sreg_n_434;
  wire sreg_n_435;
  wire sreg_n_436;
  wire sreg_n_437;
  wire sreg_n_438;
  wire sreg_n_439;
  wire sreg_n_440;
  wire sreg_n_441;
  wire sreg_n_442;
  wire sreg_n_443;
  wire sreg_n_444;
  wire sreg_n_445;
  wire sreg_n_446;
  wire sreg_n_447;
  wire sreg_n_448;
  wire sreg_n_449;
  wire sreg_n_45;
  wire sreg_n_451;
  wire sreg_n_452;
  wire sreg_n_466;
  wire sreg_n_467;
  wire sreg_n_468;
  wire sreg_n_469;
  wire sreg_n_47;
  wire sreg_n_54;
  wire sreg_n_55;
  wire sreg_n_57;
  wire sreg_n_62;
  wire sreg_n_64;
  wire sreg_n_65;
  wire sreg_n_66;
  wire sreg_n_67;
  wire sreg_n_68;
  wire sreg_n_69;
  wire sreg_n_70;
  wire sreg_n_73;
  wire sreg_n_74;
  wire sreg_n_75;
  wire sreg_n_76;
  wire sreg_n_77;
  wire sreg_n_79;
  wire sreg_n_80;
  wire sreg_n_84;
  wire sreg_n_85;
  wire sreg_n_86;
  wire sreg_n_94;
  wire sreg_n_95;
  wire sreg_n_99;
  wire [1:0]\stat[0]_i_6 ;
  wire \stat_reg[0] ;
  wire \stat_reg[1] ;
  wire \tr[16]_i_6 ;
  wire \tr[16]_i_6_0 ;
  wire \tr[17]_i_2 ;
  wire \tr[17]_i_9 ;
  wire \tr[18]_i_2 ;
  wire \tr[18]_i_9 ;
  wire \tr[19]_i_2 ;
  wire \tr[19]_i_2_0 ;
  wire \tr[19]_i_2_1 ;
  wire \tr[19]_i_3 ;
  wire \tr[19]_i_3_0 ;
  wire \tr[20]_i_2 ;
  wire \tr[20]_i_3 ;
  wire \tr[20]_i_9 ;
  wire \tr[21]_i_2 ;
  wire \tr[21]_i_3 ;
  wire \tr[22]_i_11 ;
  wire \tr[22]_i_2 ;
  wire \tr[22]_i_3 ;
  wire \tr[22]_i_9 ;
  wire \tr[23]_i_2 ;
  wire \tr[24]_i_10 ;
  wire \tr[24]_i_2 ;
  wire \tr[24]_i_3 ;
  wire \tr[24]_i_3_0 ;
  wire \tr[25]_i_2 ;
  wire \tr[26]_i_3 ;
  wire \tr[26]_i_9 ;
  wire \tr[28]_i_2 ;
  wire [5:0]\tr[29]_i_2 ;
  wire \tr[29]_i_3 ;
  wire \tr[30]_i_10 ;
  wire \tr[30]_i_3 ;
  wire \tr[30]_i_3_0 ;
  wire [1:0]\tr_reg[0] ;
  wire \tr_reg[16] ;
  wire \tr_reg[17] ;
  wire \tr_reg[18] ;
  wire \tr_reg[19] ;
  wire \tr_reg[19]_0 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[20] ;
  wire \tr_reg[21] ;
  wire \tr_reg[21]_0 ;
  wire \tr_reg[22] ;
  wire \tr_reg[23] ;
  wire \tr_reg[23]_0 ;
  wire \tr_reg[23]_i_11 ;
  wire \tr_reg[23]_i_11_0 ;
  wire \tr_reg[23]_i_11_1 ;
  wire \tr_reg[23]_i_11_2 ;
  wire \tr_reg[24] ;
  wire \tr_reg[25] ;
  wire \tr_reg[26] ;
  wire \tr_reg[27] ;
  wire \tr_reg[27]_0 ;
  wire \tr_reg[27]_1 ;
  wire \tr_reg[28] ;
  wire \tr_reg[28]_0 ;
  wire \tr_reg[29] ;
  wire \tr_reg[29]_0 ;
  wire \tr_reg[30] ;
  wire [31:0]\tr_reg[31] ;
  wire \tr_reg[31]_0 ;
  wire \tr_reg[31]_1 ;
  wire \tr_reg[31]_2 ;
  wire \tr_reg[31]_i_13 ;
  wire \tr_reg[31]_i_13_0 ;
  wire \tr_reg[31]_i_13_1 ;
  wire \tr_reg[31]_i_32 ;
  wire \tr_reg[31]_i_32_0 ;
  wire \tr_reg[31]_i_32_1 ;
  wire \tr_reg[31]_i_32_2 ;
  wire [1:0]\tr_reg[5] ;

  niho_rgf_bus abus_out
       (.DI(abus_0[15:12]),
        .abus_sel_cr(abus_sel_cr),
        .abus_sp(abus_sp),
        .\mul_a_reg[0] (\mul_a_reg[0] ),
        .\mul_a_reg[0]_0 (bank13_n_134),
        .\mul_a_reg[0]_1 (bank13_n_150),
        .\mul_a_reg[0]_2 (bank13_n_96),
        .\mul_a_reg[0]_3 (bank13_n_80),
        .\mul_a_reg[10] (\mul_a_reg[10] ),
        .\mul_a_reg[10]_0 (bank13_n_124),
        .\mul_a_reg[10]_1 (bank13_n_140),
        .\mul_a_reg[10]_2 (bank13_n_86),
        .\mul_a_reg[10]_3 (bank13_n_70),
        .\mul_a_reg[11] (\mul_a_reg[11] ),
        .\mul_a_reg[11]_0 (bank13_n_123),
        .\mul_a_reg[11]_1 (bank13_n_139),
        .\mul_a_reg[11]_2 (bank13_n_85),
        .\mul_a_reg[11]_3 (bank13_n_69),
        .\mul_a_reg[12] (\mul_a_reg[12] ),
        .\mul_a_reg[12]_0 (bank13_n_122),
        .\mul_a_reg[12]_1 (bank13_n_138),
        .\mul_a_reg[12]_2 (bank13_n_84),
        .\mul_a_reg[12]_3 (bank13_n_68),
        .\mul_a_reg[13] (\mul_a_reg[13] ),
        .\mul_a_reg[13]_0 (bank13_n_121),
        .\mul_a_reg[13]_1 (bank13_n_137),
        .\mul_a_reg[13]_2 (bank13_n_83),
        .\mul_a_reg[13]_3 (bank13_n_67),
        .\mul_a_reg[14] (\mul_a_reg[14] ),
        .\mul_a_reg[14]_0 (bank13_n_120),
        .\mul_a_reg[14]_1 (bank13_n_136),
        .\mul_a_reg[14]_2 (bank13_n_82),
        .\mul_a_reg[14]_3 (bank13_n_66),
        .\mul_a_reg[15] (\mul_a_reg[15] ),
        .\mul_a_reg[15]_0 (bank13_n_119),
        .\mul_a_reg[15]_1 (bank13_n_135),
        .\mul_a_reg[15]_2 (bank13_n_81),
        .\mul_a_reg[15]_3 (bank13_n_65),
        .\mul_a_reg[15]_4 ({p_0_in_1[15:1],\sp_reg[0] }),
        .\mul_a_reg[16] (\mul_a_reg[16] ),
        .\mul_a_reg[16]_0 (bank02_n_474),
        .\mul_a_reg[16]_1 (bank02_n_490),
        .\mul_a_reg[16]_2 (bank13_n_188),
        .\mul_a_reg[16]_3 (bank13_n_204),
        .\mul_a_reg[17] (\mul_a_reg[17] ),
        .\mul_a_reg[17]_0 (bank02_n_473),
        .\mul_a_reg[17]_1 (bank02_n_489),
        .\mul_a_reg[17]_2 (bank13_n_187),
        .\mul_a_reg[17]_3 (bank13_n_203),
        .\mul_a_reg[18] (\mul_a_reg[18] ),
        .\mul_a_reg[18]_0 (bank02_n_472),
        .\mul_a_reg[18]_1 (bank02_n_488),
        .\mul_a_reg[18]_2 (bank13_n_186),
        .\mul_a_reg[18]_3 (bank13_n_202),
        .\mul_a_reg[19] (\mul_a_reg[19] ),
        .\mul_a_reg[19]_0 (bank02_n_471),
        .\mul_a_reg[19]_1 (bank02_n_487),
        .\mul_a_reg[19]_2 (bank13_n_185),
        .\mul_a_reg[19]_3 (bank13_n_201),
        .\mul_a_reg[1] (\mul_a_reg[1] ),
        .\mul_a_reg[1]_0 (bank13_n_133),
        .\mul_a_reg[1]_1 (bank13_n_149),
        .\mul_a_reg[1]_2 (bank13_n_95),
        .\mul_a_reg[1]_3 (bank13_n_79),
        .\mul_a_reg[20] (\mul_a_reg[20] ),
        .\mul_a_reg[20]_0 (bank02_n_470),
        .\mul_a_reg[20]_1 (bank02_n_486),
        .\mul_a_reg[20]_2 (bank13_n_184),
        .\mul_a_reg[20]_3 (bank13_n_200),
        .\mul_a_reg[21] (\mul_a_reg[21] ),
        .\mul_a_reg[21]_0 (bank02_n_469),
        .\mul_a_reg[21]_1 (bank02_n_485),
        .\mul_a_reg[21]_2 (bank13_n_183),
        .\mul_a_reg[21]_3 (bank13_n_199),
        .\mul_a_reg[22] (\mul_a_reg[22] ),
        .\mul_a_reg[22]_0 (bank02_n_468),
        .\mul_a_reg[22]_1 (bank02_n_484),
        .\mul_a_reg[22]_2 (bank13_n_182),
        .\mul_a_reg[22]_3 (bank13_n_198),
        .\mul_a_reg[23] (\mul_a_reg[23] ),
        .\mul_a_reg[23]_0 (bank02_n_467),
        .\mul_a_reg[23]_1 (bank02_n_483),
        .\mul_a_reg[23]_2 (bank13_n_181),
        .\mul_a_reg[23]_3 (bank13_n_197),
        .\mul_a_reg[24] (\mul_a_reg[24] ),
        .\mul_a_reg[24]_0 (bank02_n_466),
        .\mul_a_reg[24]_1 (bank02_n_482),
        .\mul_a_reg[24]_2 (bank13_n_180),
        .\mul_a_reg[24]_3 (bank13_n_196),
        .\mul_a_reg[25] (\mul_a_reg[25] ),
        .\mul_a_reg[25]_0 (bank02_n_465),
        .\mul_a_reg[25]_1 (bank02_n_481),
        .\mul_a_reg[25]_2 (bank13_n_179),
        .\mul_a_reg[25]_3 (bank13_n_195),
        .\mul_a_reg[26] (\mul_a_reg[26] ),
        .\mul_a_reg[26]_0 (bank02_n_464),
        .\mul_a_reg[26]_1 (bank02_n_480),
        .\mul_a_reg[26]_2 (bank13_n_178),
        .\mul_a_reg[26]_3 (bank13_n_194),
        .\mul_a_reg[27] (\mul_a_reg[27] ),
        .\mul_a_reg[27]_0 (bank02_n_463),
        .\mul_a_reg[27]_1 (bank02_n_479),
        .\mul_a_reg[27]_2 (bank13_n_177),
        .\mul_a_reg[27]_3 (bank13_n_193),
        .\mul_a_reg[28] (\mul_a_reg[28] ),
        .\mul_a_reg[28]_0 (bank02_n_462),
        .\mul_a_reg[28]_1 (bank02_n_478),
        .\mul_a_reg[28]_2 (bank13_n_176),
        .\mul_a_reg[28]_3 (bank13_n_192),
        .\mul_a_reg[29] (\mul_a_reg[29] ),
        .\mul_a_reg[29]_0 (bank02_n_461),
        .\mul_a_reg[29]_1 (bank02_n_477),
        .\mul_a_reg[29]_2 (bank13_n_175),
        .\mul_a_reg[29]_3 (bank13_n_191),
        .\mul_a_reg[2] (\mul_a_reg[2] ),
        .\mul_a_reg[2]_0 (bank13_n_132),
        .\mul_a_reg[2]_1 (bank13_n_148),
        .\mul_a_reg[2]_2 (bank13_n_94),
        .\mul_a_reg[2]_3 (bank13_n_78),
        .\mul_a_reg[30] (\mul_a_reg[30] ),
        .\mul_a_reg[30]_0 (bank02_n_460),
        .\mul_a_reg[30]_1 (bank02_n_476),
        .\mul_a_reg[30]_2 (bank13_n_174),
        .\mul_a_reg[30]_3 (bank13_n_190),
        .\mul_a_reg[32] (\mul_a_reg[32]_0 ),
        .\mul_a_reg[32]_0 (bank02_n_459),
        .\mul_a_reg[32]_1 (bank02_n_475),
        .\mul_a_reg[32]_2 (bank13_n_173),
        .\mul_a_reg[32]_3 (bank13_n_189),
        .\mul_a_reg[3] (\mul_a_reg[3] ),
        .\mul_a_reg[3]_0 (bank13_n_131),
        .\mul_a_reg[3]_1 (bank13_n_147),
        .\mul_a_reg[3]_2 (bank13_n_93),
        .\mul_a_reg[3]_3 (bank13_n_77),
        .\mul_a_reg[4] (\mul_a_reg[4] ),
        .\mul_a_reg[4]_0 (bank13_n_130),
        .\mul_a_reg[4]_1 (bank13_n_146),
        .\mul_a_reg[4]_2 (bank13_n_92),
        .\mul_a_reg[4]_3 (bank13_n_76),
        .\mul_a_reg[5] (\mul_a_reg[5] ),
        .\mul_a_reg[5]_0 (bank13_n_129),
        .\mul_a_reg[5]_1 (bank13_n_145),
        .\mul_a_reg[5]_2 (bank13_n_91),
        .\mul_a_reg[5]_3 (bank13_n_75),
        .\mul_a_reg[6] (\mul_a_reg[6] ),
        .\mul_a_reg[6]_0 (bank13_n_128),
        .\mul_a_reg[6]_1 (bank13_n_144),
        .\mul_a_reg[6]_2 (bank13_n_90),
        .\mul_a_reg[6]_3 (bank13_n_74),
        .\mul_a_reg[7] (\mul_a_reg[7] ),
        .\mul_a_reg[7]_0 (bank13_n_127),
        .\mul_a_reg[7]_1 (bank13_n_143),
        .\mul_a_reg[7]_2 (bank13_n_89),
        .\mul_a_reg[7]_3 (bank13_n_73),
        .\mul_a_reg[8] (\mul_a_reg[8] ),
        .\mul_a_reg[8]_0 (bank13_n_126),
        .\mul_a_reg[8]_1 (bank13_n_142),
        .\mul_a_reg[8]_2 (bank13_n_88),
        .\mul_a_reg[8]_3 (bank13_n_72),
        .\mul_a_reg[9] (\mul_a_reg[9] ),
        .\mul_a_reg[9]_0 (bank13_n_125),
        .\mul_a_reg[9]_1 (bank13_n_141),
        .\mul_a_reg[9]_2 (bank13_n_87),
        .\mul_a_reg[9]_3 (bank13_n_71),
        .out({p_0_in_2[15:14],out[12:9],p_0_in_2[9],out[8:0]}),
        .p_0_in(p_0_in_0),
        .p_1_in(p_1_in),
        .rgf_pc(rgf_pc),
        .sp_dec_0(sp_dec_0[15:1]),
        .\sp_reg[15] (abus_out_n_5),
        .\sr_reg[15] (abus_out_n_4),
        .\tr_reg[11] (abus_0[11:8]),
        .\tr_reg[16] (abus_0[16]),
        .\tr_reg[17] (abus_0[17]),
        .\tr_reg[18] (abus_0[18]),
        .\tr_reg[19] (abus_0[19]),
        .\tr_reg[20] (abus_0[20]),
        .\tr_reg[21] (abus_0[21]),
        .\tr_reg[22] (abus_0[22]),
        .\tr_reg[23] (abus_0[23]),
        .\tr_reg[24] (abus_0[24]),
        .\tr_reg[25] (abus_0[25]),
        .\tr_reg[26] (abus_0[26]),
        .\tr_reg[27] (abus_0[27]),
        .\tr_reg[28] (abus_0[28]),
        .\tr_reg[29] (abus_0[29]),
        .\tr_reg[30] (abus_0[30]),
        .\tr_reg[31] (abus_0[31]),
        .\tr_reg[3] (abus_0[3:0]),
        .\tr_reg[7] (abus_0[7:4]));
  niho_rgf_bank bank02
       (.CO(bank02_n_364),
        .DI(abus_0[15:12]),
        .E(E),
        .S(S),
        .SR(p_0_in),
        .abus_o(abus_o[15:0]),
        .\abus_o[11] (abus_0[11:8]),
        .\abus_o[3] (abus_0[3:0]),
        .\abus_o[7] (abus_0[7:4]),
        .abus_o_0_sp_1(abus_o_16_sn_1),
        .abus_sel_0(abus_sel_0),
        .\art/add/iv[7]_i_32 (\art/add/iv[7]_i_32 ),
        .\art/add/sr[5]_i_14 (\art/add/sr[5]_i_14 ),
        .\art/add/sr[5]_i_18 (\art/add/sr[5]_i_18 ),
        .\badr[0]_INST_0_i_1 (\badr[0]_INST_0_i_1 ),
        .\badr[0]_INST_0_i_1_0 (bank02_n_283),
        .\badr[14]_INST_0_i_1 (bank02_n_259),
        .\badr[14]_INST_0_i_1_0 (bank02_n_279),
        .\badr[15]_INST_0_i_1 (bank02_n_264),
        .\badr[16]_INST_0_i_1 (bank02_n_284),
        .\badr[16]_INST_0_i_1_0 (sreg_n_397),
        .\badr[16]_INST_0_i_1_1 (sreg_n_381),
        .\badr[17]_INST_0_i_1 (sreg_n_398),
        .\badr[17]_INST_0_i_1_0 (sreg_n_382),
        .\badr[18]_INST_0_i_1 (sreg_n_399),
        .\badr[18]_INST_0_i_1_0 (sreg_n_383),
        .\badr[19]_INST_0_i_1 (sreg_n_400),
        .\badr[19]_INST_0_i_1_0 (sreg_n_384),
        .\badr[20]_INST_0_i_1 (sreg_n_401),
        .\badr[20]_INST_0_i_1_0 (sreg_n_385),
        .\badr[21]_INST_0_i_1 (\badr[21]_INST_0_i_1 ),
        .\badr[21]_INST_0_i_1_0 (sreg_n_402),
        .\badr[21]_INST_0_i_1_1 (sreg_n_386),
        .\badr[22]_INST_0_i_1 (sreg_n_403),
        .\badr[22]_INST_0_i_1_0 (sreg_n_387),
        .\badr[23]_INST_0_i_1 (sreg_n_404),
        .\badr[23]_INST_0_i_1_0 (sreg_n_388),
        .\badr[24]_INST_0_i_1 (sreg_n_405),
        .\badr[24]_INST_0_i_1_0 (sreg_n_389),
        .\badr[25]_INST_0_i_1 (sreg_n_406),
        .\badr[25]_INST_0_i_1_0 (sreg_n_390),
        .\badr[26]_INST_0_i_1 (sreg_n_407),
        .\badr[26]_INST_0_i_1_0 (sreg_n_391),
        .\badr[27]_INST_0_i_1 (sreg_n_408),
        .\badr[27]_INST_0_i_1_0 (sreg_n_392),
        .\badr[28]_INST_0_i_1 (sreg_n_409),
        .\badr[28]_INST_0_i_1_0 (sreg_n_393),
        .\badr[29]_INST_0_i_1 (sreg_n_410),
        .\badr[29]_INST_0_i_1_0 (sreg_n_394),
        .\badr[30]_INST_0_i_1 (sreg_n_411),
        .\badr[30]_INST_0_i_1_0 (sreg_n_395),
        .\badr[31]_INST_0_i_1 (sreg_n_412),
        .\badr[31]_INST_0_i_1_0 (sreg_n_396),
        .\badr[5]_INST_0_i_1 (\badr[5]_INST_0_i_1 ),
        .bank_sel(bank_sel),
        .bbus_0({bbus_0[4:2],bbus_0[0]}),
        .bbus_o(bbus_o),
        .bbus_sel_0({bbus_sel_0[7],bbus_sel_0[4:0]}),
        .\bdatw[8]_INST_0_i_2 (\bdatw[8]_INST_0_i_2 ),
        .cbus(cbus[15:0]),
        .clk(clk),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .\grn_reg[0] (bank02_n_430),
        .\grn_reg[0]_0 (bank02_n_436),
        .\grn_reg[0]_1 (bank02_n_452),
        .\grn_reg[0]_2 (bank02_n_458),
        .\grn_reg[0]_3 (bank02_n_474),
        .\grn_reg[0]_4 (bank02_n_490),
        .\grn_reg[0]_5 (sreg_n_284),
        .\grn_reg[0]_6 (sreg_n_16),
        .\grn_reg[0]_7 (sreg_n_282),
        .\grn_reg[0]_8 (sreg_n_18),
        .\grn_reg[10] (bank02_n_420),
        .\grn_reg[10]_0 (bank02_n_442),
        .\grn_reg[10]_1 (bank02_n_464),
        .\grn_reg[10]_2 (bank02_n_480),
        .\grn_reg[11] (bank02_n_419),
        .\grn_reg[11]_0 (bank02_n_441),
        .\grn_reg[11]_1 (bank02_n_463),
        .\grn_reg[11]_2 (bank02_n_479),
        .\grn_reg[12] (bank02_n_418),
        .\grn_reg[12]_0 (bank02_n_440),
        .\grn_reg[12]_1 (bank02_n_462),
        .\grn_reg[12]_2 (bank02_n_478),
        .\grn_reg[13] (bank02_n_417),
        .\grn_reg[13]_0 (bank02_n_439),
        .\grn_reg[13]_1 (bank02_n_461),
        .\grn_reg[13]_2 (bank02_n_477),
        .\grn_reg[14] (bank02_n_416),
        .\grn_reg[14]_0 (bank02_n_438),
        .\grn_reg[14]_1 (bank02_n_460),
        .\grn_reg[14]_2 (bank02_n_476),
        .\grn_reg[15] ({bank02_n_16,bank02_n_17,bank02_n_18,bank02_n_19,bank02_n_20,bank02_n_21,bank02_n_22,bank02_n_23,bank02_n_24,bank02_n_25,bank02_n_26,bank02_n_27,bank02_n_28,bank02_n_29,bank02_n_30,bank02_n_31}),
        .\grn_reg[15]_0 ({bank02_n_32,bank02_n_33,bank02_n_34,bank02_n_35,bank02_n_36,bank02_n_37,bank02_n_38,bank02_n_39,bank02_n_40,bank02_n_41,bank02_n_42,bank02_n_43,bank02_n_44,bank02_n_45,bank02_n_46,bank02_n_47}),
        .\grn_reg[15]_1 ({bank02_n_48,bank02_n_49,bank02_n_50,bank02_n_51,bank02_n_52,bank02_n_53,bank02_n_54,bank02_n_55,bank02_n_56,bank02_n_57,bank02_n_58,bank02_n_59,bank02_n_60,bank02_n_61,bank02_n_62,bank02_n_63}),
        .\grn_reg[15]_10 (\grn_reg[15] ),
        .\grn_reg[15]_11 (\grn_reg[15]_0 ),
        .\grn_reg[15]_12 (\grn_reg[15]_1 ),
        .\grn_reg[15]_13 (\grn_reg[15]_2 ),
        .\grn_reg[15]_14 (\grn_reg[15]_3 ),
        .\grn_reg[15]_15 (\grn_reg[15]_4 ),
        .\grn_reg[15]_16 (\grn_reg[15]_5 ),
        .\grn_reg[15]_17 (\grn_reg[15]_6 ),
        .\grn_reg[15]_18 (\grn_reg[15]_7 ),
        .\grn_reg[15]_19 (\grn_reg[15]_8 ),
        .\grn_reg[15]_2 ({bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72,bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78,bank02_n_79}),
        .\grn_reg[15]_20 (\grn_reg[15]_9 ),
        .\grn_reg[15]_21 (\grn_reg[15]_10 ),
        .\grn_reg[15]_3 ({bank02_n_80,bank02_n_81,bank02_n_82,bank02_n_83,bank02_n_84,bank02_n_85,bank02_n_86,bank02_n_87,bank02_n_88,bank02_n_89,bank02_n_90,bank02_n_91,bank02_n_92,bank02_n_93,bank02_n_94,bank02_n_95}),
        .\grn_reg[15]_4 ({bank02_n_96,bank02_n_97,bank02_n_98,bank02_n_99,bank02_n_100,bank02_n_101,bank02_n_102,bank02_n_103,bank02_n_104,bank02_n_105,bank02_n_106,bank02_n_107,bank02_n_108,bank02_n_109,bank02_n_110,bank02_n_111}),
        .\grn_reg[15]_5 ({bank02_n_112,bank02_n_113,bank02_n_114,bank02_n_115,bank02_n_116,bank02_n_117,bank02_n_118,bank02_n_119,bank02_n_120,bank02_n_121,bank02_n_122,bank02_n_123,bank02_n_124,bank02_n_125,bank02_n_126,bank02_n_127}),
        .\grn_reg[15]_6 (bank02_n_415),
        .\grn_reg[15]_7 (bank02_n_437),
        .\grn_reg[15]_8 (bank02_n_459),
        .\grn_reg[15]_9 (bank02_n_475),
        .\grn_reg[1] (bank02_n_429),
        .\grn_reg[1]_0 (bank02_n_435),
        .\grn_reg[1]_1 (bank02_n_451),
        .\grn_reg[1]_2 (bank02_n_457),
        .\grn_reg[1]_3 (bank02_n_473),
        .\grn_reg[1]_4 (bank02_n_489),
        .\grn_reg[2] (bank02_n_428),
        .\grn_reg[2]_0 (bank02_n_434),
        .\grn_reg[2]_1 (bank02_n_450),
        .\grn_reg[2]_2 (bank02_n_456),
        .\grn_reg[2]_3 (bank02_n_472),
        .\grn_reg[2]_4 (bank02_n_488),
        .\grn_reg[3] (bank02_n_427),
        .\grn_reg[3]_0 (bank02_n_433),
        .\grn_reg[3]_1 (bank02_n_449),
        .\grn_reg[3]_2 (bank02_n_455),
        .\grn_reg[3]_3 (bank02_n_471),
        .\grn_reg[3]_4 (bank02_n_487),
        .\grn_reg[4] (bank02_n_426),
        .\grn_reg[4]_0 (bank02_n_432),
        .\grn_reg[4]_1 (bank02_n_448),
        .\grn_reg[4]_2 (bank02_n_454),
        .\grn_reg[4]_3 (bank02_n_470),
        .\grn_reg[4]_4 (bank02_n_486),
        .\grn_reg[5] (bank02_n_425),
        .\grn_reg[5]_0 (bank02_n_431),
        .\grn_reg[5]_1 (bank02_n_447),
        .\grn_reg[5]_2 (bank02_n_453),
        .\grn_reg[5]_3 (bank02_n_469),
        .\grn_reg[5]_4 (bank02_n_485),
        .\grn_reg[6] (bank02_n_424),
        .\grn_reg[6]_0 (bank02_n_446),
        .\grn_reg[6]_1 (bank02_n_468),
        .\grn_reg[6]_2 (bank02_n_484),
        .\grn_reg[7] (bank02_n_423),
        .\grn_reg[7]_0 (bank02_n_445),
        .\grn_reg[7]_1 (bank02_n_467),
        .\grn_reg[7]_2 (bank02_n_483),
        .\grn_reg[8] (bank02_n_422),
        .\grn_reg[8]_0 (bank02_n_444),
        .\grn_reg[8]_1 (bank02_n_466),
        .\grn_reg[8]_2 (bank02_n_482),
        .\grn_reg[9] (bank02_n_421),
        .\grn_reg[9]_0 (bank02_n_443),
        .\grn_reg[9]_1 (bank02_n_465),
        .\grn_reg[9]_2 (bank02_n_481),
        .\i_/badr[15]_INST_0_i_15 (sreg_n_276),
        .\i_/bdatw[15]_INST_0_i_65 (\i_/bdatw[15]_INST_0_i_65 ),
        .\i_/bdatw[15]_INST_0_i_65_0 (\i_/bdatw[15]_INST_0_i_65_0 ),
        .\i_/bdatw[15]_INST_0_i_65_1 (\i_/bdatw[15]_INST_0_i_65_1 ),
        .\i_/bdatw[15]_INST_0_i_65_2 (\i_/bdatw[15]_INST_0_i_65_2 ),
        .\iv[0]_i_10_0 (\iv[0]_i_10 ),
        .\iv[0]_i_10_1 (\iv[0]_i_10_0 ),
        .\iv[0]_i_10_2 (\iv[0]_i_10_1 ),
        .\iv[0]_i_10_3 (sreg_n_142),
        .\iv[0]_i_19 (\iv[0]_i_19 ),
        .\iv[0]_i_22_0 (sreg_n_109),
        .\iv[0]_i_25 (\iv[0]_i_25 ),
        .\iv[0]_i_3 (\iv[0]_i_3 ),
        .\iv[0]_i_3_0 (sreg_n_75),
        .\iv[0]_i_3_1 (\iv[0]_i_3_1 ),
        .\iv[0]_i_6 (\iv[0]_i_6 ),
        .\iv[0]_i_6_0 (\iv[0]_i_6_0 ),
        .\iv[0]_i_7 (\iv[0]_i_7 ),
        .\iv[0]_i_8 (sreg_n_103),
        .\iv[0]_i_8_0 (sreg_n_102),
        .\iv[10]_i_10 (\iv[10]_i_10 ),
        .\iv[10]_i_10_0 (sreg_n_118),
        .\iv[10]_i_13 (sreg_n_145),
        .\iv[10]_i_2 (\iv[10]_i_2 ),
        .\iv[10]_i_22_0 (sreg_n_119),
        .\iv[10]_i_25 (sreg_n_157),
        .\iv[10]_i_2_0 (sreg_n_43),
        .\iv[10]_i_5 (\iv[10]_i_5 ),
        .\iv[11]_i_13 (sreg_n_128),
        .\iv[11]_i_25 (sreg_n_150),
        .\iv[12]_i_13 (sreg_n_143),
        .\iv[12]_i_2 (\iv[12]_i_2 ),
        .\iv[12]_i_27_0 (bank02_n_181),
        .\iv[13]_i_13 (sreg_n_123),
        .\iv[13]_i_17 (\iv[13]_i_17 ),
        .\iv[13]_i_17_0 (\iv[13]_i_17_0 ),
        .\iv[13]_i_17_1 (abus_0[21]),
        .\iv[13]_i_2 (\iv[13]_i_2 ),
        .\iv[13]_i_26 (sreg_n_151),
        .\iv[13]_i_26_0 (sreg_n_125),
        .\iv[13]_i_27 (\iv[13]_i_27 ),
        .\iv[13]_i_29_0 (bank02_n_182),
        .\iv[14]_i_32_0 (abus_0[30]),
        .\iv[14]_i_35_0 (\iv[14]_i_35 ),
        .\iv[14]_i_49 (\iv[14]_i_49 ),
        .\iv[14]_i_5 (\iv[14]_i_5 ),
        .\iv[15]_i_108 (\iv[15]_i_108 ),
        .\iv[15]_i_108_0 (\iv[15]_i_108_0 ),
        .\iv[15]_i_108_1 (\iv[15]_i_108_1 ),
        .\iv[15]_i_108_2 (\iv[15]_i_108_2 ),
        .\iv[15]_i_108_3 (\iv[15]_i_108_3 ),
        .\iv[15]_i_108_4 (\iv[15]_i_108_4 ),
        .\iv[15]_i_108_5 (\iv[15]_i_108_5 ),
        .\iv[15]_i_108_6 (\iv[15]_i_108_6 ),
        .\iv[15]_i_108_7 (\iv[15]_i_108_7 ),
        .\iv[15]_i_108_8 (\iv[15]_i_108_8 ),
        .\iv[15]_i_22_0 (sreg_n_148),
        .\iv[15]_i_60_0 (sreg_n_127),
        .\iv[15]_i_8 (\sr_reg[8]_36 ),
        .\iv[15]_i_8_0 (\iv[15]_i_8 ),
        .\iv[15]_i_8_1 (\iv[15]_i_8_0 ),
        .\iv[15]_i_8_2 (\iv[15]_i_8_1 ),
        .\iv[15]_i_94 (bank02_n_196),
        .\iv[1]_i_10 (\iv[1]_i_10 ),
        .\iv[1]_i_10_0 (\iv[1]_i_10_0 ),
        .\iv[1]_i_10_1 (\iv[1]_i_10_1 ),
        .\iv[1]_i_9 (\iv[1]_i_9 ),
        .\iv[2]_i_24 (sreg_n_156),
        .\iv[2]_i_9 (\iv[2]_i_9 ),
        .\iv[3]_i_10 (\iv[3]_i_10 ),
        .\iv[3]_i_10_0 (\iv[3]_i_10_0 ),
        .\iv[3]_i_10_1 (\iv[3]_i_10_1 ),
        .\iv[3]_i_15 (sreg_n_153),
        .\iv[3]_i_31 (sreg_n_149),
        .\iv[3]_i_9 (\iv[3]_i_9 ),
        .\iv[4]_i_14 (sreg_n_146),
        .\iv[4]_i_31 (\sr_reg[8]_125 ),
        .\iv[4]_i_6 (\iv[4]_i_6 ),
        .\iv[4]_i_9 (\iv[4]_i_9 ),
        .\iv[5]_i_14 (sreg_n_129),
        .\iv[5]_i_23 (bank02_n_203),
        .\iv[5]_i_30 (sreg_n_126),
        .\iv[5]_i_9 (\iv[5]_i_9 ),
        .\iv[6]_i_10 (\iv[6]_i_10 ),
        .\iv[6]_i_10_0 (\iv[6]_i_10_0 ),
        .\iv[6]_i_10_1 (\iv[6]_i_10_1 ),
        .\iv[6]_i_15 (sreg_n_95),
        .\iv[7]_i_17 (\iv[7]_i_17 ),
        .\iv[7]_i_17_0 (sreg_n_80),
        .\iv[7]_i_25 (\iv[7]_i_25 ),
        .\iv[7]_i_3 (sreg_n_69),
        .\iv[7]_i_33 (\iv[7]_i_33 ),
        .\iv[7]_i_37_0 (bank02_n_144),
        .\iv[7]_i_3_0 (sreg_n_107),
        .\iv[7]_i_3_1 (\iv[7]_i_3 ),
        .\iv[7]_i_7 (\iv[7]_i_7 ),
        .\iv[7]_i_7_0 (\iv[7]_i_7_0 ),
        .\iv[7]_i_7_1 (\iv[7]_i_7_1 ),
        .\iv[7]_i_9 (\iv[7]_i_9 ),
        .\iv[8]_i_2 (\iv[8]_i_2 ),
        .\iv[8]_i_20 (\iv[8]_i_20 ),
        .\iv[8]_i_30 (bank02_n_190),
        .\iv[8]_i_5 (\iv[8]_i_5 ),
        .\iv[8]_i_8 (\iv[8]_i_8 ),
        .\iv[9]_i_11 (\iv[9]_i_11 ),
        .\iv[9]_i_11_0 (sreg_n_101),
        .\iv[9]_i_2 (sreg_n_54),
        .\iv[9]_i_5 (\iv[9]_i_5 ),
        .\iv_reg[7]_i_12_0 (\sr_reg[6]_11 ),
        .mul_a(mul_a[32:16]),
        .\mul_b_reg[0] (\mul_b_reg[0] ),
        .\mul_b_reg[0]_0 (\mul_b_reg[0]_0 ),
        .\mul_b_reg[0]_1 (bbus_out_n_17),
        .\mul_b_reg[0]_2 (bbus_out_n_35),
        .\mul_b_reg[5] (\mul_b_reg[5]_0 ),
        .\mul_b_reg[5]_0 (\mul_b_reg[5] ),
        .\mul_b_reg[5]_1 (bbus_out_n_11),
        .\mul_b_reg[5]_2 (bbus_out_n_28),
        .mul_rslt(mul_rslt),
        .niho_dsp_a(niho_dsp_a[32:16]),
        .\niho_dsp_a[15]_INST_0_i_3 (\niho_dsp_a[15]_INST_0_i_3 ),
        .\niho_dsp_a[16] ({out[8],out[6],out[1:0]}),
        .\niho_dsp_a[16]_0 (\mul_a_reg[32] ),
        .\niho_dsp_a[32] (abus_out_n_5),
        .\niho_dsp_a[32]_0 (abus_out_n_4),
        .\niho_dsp_a[32]_1 (\mul_a_reg[15] ),
        .niho_dsp_c(niho_dsp_c),
        .out({bank02_n_0,bank02_n_1,bank02_n_2,bank02_n_3,bank02_n_4,bank02_n_5,bank02_n_6,bank02_n_7,bank02_n_8,bank02_n_9,bank02_n_10,bank02_n_11,bank02_n_12,bank02_n_13,bank02_n_14,bank02_n_15}),
        .p_0_in(p_0_in_0),
        .p_1_in(p_1_in),
        .p_2_in(p_2_in[5:0]),
        .\sr[4]_i_104_0 (sreg_n_132),
        .\sr[4]_i_108_0 (sreg_n_113),
        .\sr[4]_i_116_0 (\sr[4]_i_116 ),
        .\sr[4]_i_147_0 (\sr[4]_i_147 ),
        .\sr[4]_i_152 (sreg_n_131),
        .\sr[4]_i_152_0 (sreg_n_130),
        .\sr[4]_i_16_0 (\sr[4]_i_16_0 ),
        .\sr[4]_i_16_1 (sreg_n_269),
        .\sr[4]_i_16_2 (sreg_n_270),
        .\sr[4]_i_16_3 (\sr[4]_i_16 ),
        .\sr[4]_i_16_4 (sreg_n_45),
        .\sr[4]_i_16_5 (sreg_n_47),
        .\sr[4]_i_17 (sreg_n_268),
        .\sr[4]_i_17_0 (\sr_reg[8]_19 ),
        .\sr[4]_i_18 (sreg_n_26),
        .\sr[4]_i_18_0 (\sr[4]_i_18 ),
        .\sr[4]_i_19_0 (sreg_n_67),
        .\sr[4]_i_19_1 (sreg_n_263),
        .\sr[4]_i_19_2 (\sr[4]_i_19 ),
        .\sr[4]_i_20_0 (\sr[4]_i_20 ),
        .\sr[4]_i_20_1 (\sr[4]_i_20_0 ),
        .\sr[4]_i_20_2 (\sr[4]_i_20_1 ),
        .\sr[4]_i_20_3 (\sr[4]_i_20_2 ),
        .\sr[4]_i_21_0 (\sr[4]_i_21 ),
        .\sr[4]_i_21_1 (sreg_n_265),
        .\sr[4]_i_21_2 (\sr[4]_i_21_0 ),
        .\sr[4]_i_21_3 (\sr[4]_i_21_1 ),
        .\sr[4]_i_21_4 (sreg_n_266),
        .\sr[4]_i_21_5 (sreg_n_65),
        .\sr[4]_i_33_0 (\sr[4]_i_33 ),
        .\sr[4]_i_35_0 (\sr[4]_i_35 ),
        .\sr[4]_i_36 (abus_0[31]),
        .\sr[4]_i_36_0 (\sr[4]_i_36 ),
        .\sr[4]_i_37 (\sr_reg[8]_30 ),
        .\sr[4]_i_38_0 (\sr[4]_i_38 ),
        .\sr[4]_i_38_1 (\sr_reg[8]_33 ),
        .\sr[4]_i_39 (\sr_reg[8]_25 ),
        .\sr[4]_i_39_0 (\sr[4]_i_39 ),
        .\sr[4]_i_40 (\sr[4]_i_40 ),
        .\sr[4]_i_41_0 (\sr[4]_i_41 ),
        .\sr[4]_i_42 (sreg_n_79),
        .\sr[4]_i_43 (\sr_reg[8]_8 ),
        .\sr[4]_i_43_0 (\sr_reg[8]_9 ),
        .\sr[4]_i_43_1 (\sr[4]_i_43_0 ),
        .\sr[4]_i_44_0 (\sr[4]_i_44 ),
        .\sr[4]_i_44_1 (\sr[4]_i_44_0 ),
        .\sr[4]_i_44_2 (\sr[4]_i_44_1 ),
        .\sr[4]_i_45_0 (\sr[4]_i_45 ),
        .\sr[4]_i_45_1 (\sr[4]_i_45_0 ),
        .\sr[4]_i_45_2 (\sr_reg[8]_114 ),
        .\sr[4]_i_4_0 (\sr_reg[8]_0 ),
        .\sr[4]_i_51_0 (bank02_n_347),
        .\sr[4]_i_53_0 (sreg_n_138),
        .\sr[4]_i_58_0 (sreg_n_120),
        .\sr[4]_i_5_0 (\sr[4]_i_5 ),
        .\sr[4]_i_5_1 (sreg_n_24),
        .\sr[4]_i_5_2 (\sr[4]_i_5_0 ),
        .\sr[4]_i_5_3 (\sr[4]_i_5_1 ),
        .\sr[4]_i_5_4 (\sr[4]_i_5_2 ),
        .\sr[4]_i_5_5 (\iv[13]_i_10 ),
        .\sr[4]_i_61_0 (\sr[4]_i_61 ),
        .\sr[4]_i_64 (\sr_reg[8]_84 ),
        .\sr[4]_i_65_0 (\sr[4]_i_65 ),
        .\sr[4]_i_67 (\sr_reg[8]_88 ),
        .\sr[4]_i_75 (sreg_n_85),
        .\sr[4]_i_76_0 (sreg_n_76),
        .\sr[4]_i_80_0 (sreg_n_36),
        .\sr[4]_i_85_0 (sreg_n_122),
        .\sr[4]_i_88 (sreg_n_133),
        .\sr[4]_i_89_0 (\sr[4]_i_89 ),
        .\sr[4]_i_89_1 (sreg_n_74),
        .\sr[4]_i_98_0 (sreg_n_137),
        .\sr[6]_i_11 (sreg_n_147),
        .\sr[6]_i_11_0 (\sr[6]_i_11 ),
        .\sr[6]_i_12_0 (\sr_reg[8]_57 ),
        .\sr[6]_i_12_1 (\sr[6]_i_12 ),
        .\sr[6]_i_12_2 (\sr[6]_i_12_0 ),
        .\sr[6]_i_4 (sreg_n_152),
        .\sr[7]_i_7 (sreg_n_154),
        .\sr_reg[4] (\sr_reg[4]_2 ),
        .\sr_reg[4]_0 (\sr_reg[4]_3 ),
        .\sr_reg[6] (\sr_reg[6] ),
        .\sr_reg[6]_0 (bank02_n_261),
        .\sr_reg[6]_1 (bank02_n_267),
        .\sr_reg[6]_10 (\sr_reg[6]_7 ),
        .\sr_reg[6]_11 (\sr_reg[6]_8 ),
        .\sr_reg[6]_2 (\sr_reg[6]_0 ),
        .\sr_reg[6]_3 (bank02_n_272),
        .\sr_reg[6]_4 (\sr_reg[6]_1 ),
        .\sr_reg[6]_5 (\sr_reg[6]_2 ),
        .\sr_reg[6]_6 (\sr_reg[6]_3 ),
        .\sr_reg[6]_7 (bank02_n_300),
        .\sr_reg[6]_8 (\sr_reg[6]_4 ),
        .\sr_reg[6]_9 (\sr_reg[6]_6 ),
        .\sr_reg[8] (\sr_reg[8]_2 ),
        .\sr_reg[8]_0 (bank02_n_140),
        .\sr_reg[8]_1 (\sr_reg[8]_3 ),
        .\sr_reg[8]_10 (\sr_reg[8]_13 ),
        .\sr_reg[8]_100 (\sr_reg[8]_115 ),
        .\sr_reg[8]_101 (\sr_reg[8]_117 ),
        .\sr_reg[8]_102 (\sr_reg[8]_118 ),
        .\sr_reg[8]_103 (bank02_n_280),
        .\sr_reg[8]_104 (\sr_reg[8]_120 ),
        .\sr_reg[8]_105 (bank02_n_282),
        .\sr_reg[8]_106 (\sr_reg[8]_121 ),
        .\sr_reg[8]_107 (bank02_n_286),
        .\sr_reg[8]_108 (\sr_reg[8]_122 ),
        .\sr_reg[8]_109 (\sr_reg[8]_123 ),
        .\sr_reg[8]_11 (\sr_reg[8]_14 ),
        .\sr_reg[8]_110 (bank02_n_289),
        .\sr_reg[8]_111 (bank02_n_291),
        .\sr_reg[8]_112 (\sr_reg[8]_126 ),
        .\sr_reg[8]_113 (\sr_reg[8]_127 ),
        .\sr_reg[8]_114 (bank02_n_295),
        .\sr_reg[8]_115 (\sr_reg[8]_128 ),
        .\sr_reg[8]_116 (\sr_reg[8]_129 ),
        .\sr_reg[8]_117 (bank02_n_298),
        .\sr_reg[8]_118 (\sr_reg[8]_124 ),
        .\sr_reg[8]_119 (bank02_n_301),
        .\sr_reg[8]_12 (\sr_reg[8]_15 ),
        .\sr_reg[8]_120 (bank02_n_304),
        .\sr_reg[8]_121 (\sr_reg[8]_152 ),
        .\sr_reg[8]_122 (\sr_reg[8]_153 ),
        .\sr_reg[8]_123 (bank02_n_385),
        .\sr_reg[8]_124 (\sr_reg[8]_154 ),
        .\sr_reg[8]_125 (bank02_n_387),
        .\sr_reg[8]_126 (bank02_n_388),
        .\sr_reg[8]_127 (bank02_n_390),
        .\sr_reg[8]_128 (\sr_reg[8]_164 ),
        .\sr_reg[8]_129 (\sr_reg[8]_56 ),
        .\sr_reg[8]_13 (\sr_reg[8]_16 ),
        .\sr_reg[8]_130 (\sr_reg[8]_165 ),
        .\sr_reg[8]_131 (\sr_reg[8]_166 ),
        .\sr_reg[8]_132 (\sr_reg[8]_167 ),
        .\sr_reg[8]_14 (\sr_reg[8]_17 ),
        .\sr_reg[8]_15 (\sr_reg[8]_18 ),
        .\sr_reg[8]_16 (\sr_reg[8]_20 ),
        .\sr_reg[8]_17 (\sr_reg[8]_21 ),
        .\sr_reg[8]_18 (\sr_reg[8]_22 ),
        .\sr_reg[8]_19 (\sr_reg[8]_23 ),
        .\sr_reg[8]_2 (\sr_reg[8]_4 ),
        .\sr_reg[8]_20 (\sr_reg[8]_24 ),
        .\sr_reg[8]_21 (\sr_reg[8]_26 ),
        .\sr_reg[8]_22 (\sr_reg[8]_27 ),
        .\sr_reg[8]_23 (\sr_reg[8]_28 ),
        .\sr_reg[8]_24 (\sr_reg[8]_29 ),
        .\sr_reg[8]_25 (\sr_reg[8]_31 ),
        .\sr_reg[8]_26 (bank02_n_177),
        .\sr_reg[8]_27 (bank02_n_178),
        .\sr_reg[8]_28 (bank02_n_183),
        .\sr_reg[8]_29 (bank02_n_186),
        .\sr_reg[8]_3 (\sr_reg[8]_5 ),
        .\sr_reg[8]_30 (bank02_n_187),
        .\sr_reg[8]_31 (\sr_reg[8]_34 ),
        .\sr_reg[8]_32 (bank02_n_189),
        .\sr_reg[8]_33 (bank02_n_191),
        .\sr_reg[8]_34 (\sr_reg[8]_35 ),
        .\sr_reg[8]_35 (\sr_reg[8]_37 ),
        .\sr_reg[8]_36 (\sr_reg[8]_39 ),
        .\sr_reg[8]_37 (bank02_n_197),
        .\sr_reg[8]_38 (bank02_n_198),
        .\sr_reg[8]_39 (bank02_n_200),
        .\sr_reg[8]_4 (\sr_reg[8]_6 ),
        .\sr_reg[8]_40 (\sr_reg[8]_42 ),
        .\sr_reg[8]_41 (bank02_n_202),
        .\sr_reg[8]_42 (bank02_n_204),
        .\sr_reg[8]_43 (bank02_n_206),
        .\sr_reg[8]_44 (bank02_n_207),
        .\sr_reg[8]_45 (\sr_reg[8]_59 ),
        .\sr_reg[8]_46 (\sr_reg[8]_60 ),
        .\sr_reg[8]_47 (\sr_reg[8]_61 ),
        .\sr_reg[8]_48 (\sr_reg[8]_62 ),
        .\sr_reg[8]_49 (\sr_reg[8]_63 ),
        .\sr_reg[8]_5 (\sr_reg[8]_7 ),
        .\sr_reg[8]_50 (\sr_reg[8]_64 ),
        .\sr_reg[8]_51 (bank02_n_214),
        .\sr_reg[8]_52 (\sr_reg[8]_66 ),
        .\sr_reg[8]_53 (bank02_n_217),
        .\sr_reg[8]_54 (bank02_n_218),
        .\sr_reg[8]_55 (\sr_reg[8]_67 ),
        .\sr_reg[8]_56 (\sr_reg[8]_68 ),
        .\sr_reg[8]_57 (\sr_reg[8]_69 ),
        .\sr_reg[8]_58 (\sr_reg[8]_70 ),
        .\sr_reg[8]_59 (\sr_reg[8]_71 ),
        .\sr_reg[8]_6 (\sr_reg[8]_10 ),
        .\sr_reg[8]_60 (\sr_reg[8]_72 ),
        .\sr_reg[8]_61 (\sr_reg[8]_73 ),
        .\sr_reg[8]_62 (\sr_reg[8]_74 ),
        .\sr_reg[8]_63 (\sr_reg[8]_75 ),
        .\sr_reg[8]_64 (\sr_reg[8]_76 ),
        .\sr_reg[8]_65 (\sr_reg[8]_77 ),
        .\sr_reg[8]_66 (\sr_reg[8]_80 ),
        .\sr_reg[8]_67 (bank02_n_231),
        .\sr_reg[8]_68 (\sr_reg[8]_85 ),
        .\sr_reg[8]_69 (\sr_reg[8]_86 ),
        .\sr_reg[8]_7 (bank02_n_150),
        .\sr_reg[8]_70 (bank02_n_234),
        .\sr_reg[8]_71 (bank02_n_235),
        .\sr_reg[8]_72 (\sr_reg[8]_93 ),
        .\sr_reg[8]_73 (\sr_reg[8]_94 ),
        .\sr_reg[8]_74 (\sr_reg[8]_95 ),
        .\sr_reg[8]_75 (\sr_reg[8]_96 ),
        .\sr_reg[8]_76 (\sr_reg[8]_97 ),
        .\sr_reg[8]_77 (\sr_reg[8]_98 ),
        .\sr_reg[8]_78 (\sr_reg[8]_99 ),
        .\sr_reg[8]_79 (bank02_n_243),
        .\sr_reg[8]_8 (\sr_reg[8]_11 ),
        .\sr_reg[8]_80 (\sr_reg[8]_100 ),
        .\sr_reg[8]_81 (bank02_n_245),
        .\sr_reg[8]_82 (\sr_reg[8]_101 ),
        .\sr_reg[8]_83 (bank02_n_247),
        .\sr_reg[8]_84 (\sr_reg[8]_102 ),
        .\sr_reg[8]_85 (\sr_reg[8]_103 ),
        .\sr_reg[8]_86 (bank02_n_251),
        .\sr_reg[8]_87 (bank02_n_252),
        .\sr_reg[8]_88 (bank02_n_253),
        .\sr_reg[8]_89 (\sr_reg[8]_104 ),
        .\sr_reg[8]_9 (\sr_reg[8]_12 ),
        .\sr_reg[8]_90 (\sr_reg[8]_105 ),
        .\sr_reg[8]_91 (\sr_reg[8]_106 ),
        .\sr_reg[8]_92 (\sr_reg[8]_107 ),
        .\sr_reg[8]_93 (bank02_n_260),
        .\sr_reg[8]_94 (bank02_n_265),
        .\sr_reg[8]_95 (bank02_n_266),
        .\sr_reg[8]_96 (\sr_reg[8]_110 ),
        .\sr_reg[8]_97 (\sr_reg[8]_111 ),
        .\sr_reg[8]_98 (\sr_reg[8]_112 ),
        .\sr_reg[8]_99 (bank02_n_274),
        .\tr[16]_i_2_0 (sreg_n_84),
        .\tr[16]_i_6_0 (sreg_n_262),
        .\tr[16]_i_6_1 (sreg_n_136),
        .\tr[16]_i_6_2 (\tr[16]_i_6 ),
        .\tr[16]_i_6_3 (\tr[16]_i_6_0 ),
        .\tr[16]_i_9_0 (bank02_n_216),
        .\tr[17]_i_2 (\tr[17]_i_2 ),
        .\tr[17]_i_3_0 (abus_0[16]),
        .\tr[17]_i_3_1 (sreg_n_447),
        .\tr[17]_i_3_2 (sreg_n_264),
        .\tr[17]_i_3_3 (sreg_n_68),
        .\tr[17]_i_9_0 (\tr[17]_i_9 ),
        .\tr[18]_i_2 (\tr[18]_i_2 ),
        .\tr[18]_i_3_0 (sreg_n_452),
        .\tr[18]_i_3_1 (sreg_n_117),
        .\tr[18]_i_3_2 (abus_0[17]),
        .\tr[18]_i_3_3 (sreg_n_66),
        .\tr[18]_i_9_0 (\tr[18]_i_9 ),
        .\tr[19]_i_2_0 (\tr[19]_i_2 ),
        .\tr[19]_i_3_0 (\tr[19]_i_3 ),
        .\tr[19]_i_3_1 (sreg_n_449),
        .\tr[19]_i_3_2 (sreg_n_267),
        .\tr[19]_i_3_3 (abus_0[18]),
        .\tr[19]_i_3_4 (\tr[19]_i_3_0 ),
        .\tr[19]_i_3_5 (sreg_n_64),
        .\tr[20]_i_2 (\tr[20]_i_2 ),
        .\tr[20]_i_3_0 (sreg_n_468),
        .\tr[20]_i_3_1 (sreg_n_140),
        .\tr[20]_i_3_2 (abus_0[19]),
        .\tr[20]_i_3_3 (\tr[20]_i_3 ),
        .\tr[20]_i_9_0 (\tr[20]_i_9 ),
        .\tr[21]_i_2_0 (\tr[21]_i_2 ),
        .\tr[21]_i_3_0 (sreg_n_446),
        .\tr[21]_i_3_1 (sreg_n_108),
        .\tr[21]_i_3_2 (sreg_n_110),
        .\tr[21]_i_3_3 (abus_0[20]),
        .\tr[21]_i_3_4 (\tr[21]_i_3 ),
        .\tr[22]_i_11 (\tr[22]_i_11 ),
        .\tr[22]_i_2 (\tr[22]_i_2 ),
        .\tr[22]_i_3_0 (\tr[22]_i_3 ),
        .\tr[22]_i_3_1 (sreg_n_29),
        .\tr[22]_i_8_0 (\sr_reg[8]_116 ),
        .\tr[22]_i_9_0 (\tr[22]_i_9 ),
        .\tr[23]_i_2_0 (\tr[23]_i_2 ),
        .\tr[23]_i_2_1 (sreg_n_33),
        .\tr[23]_i_3_0 (sreg_n_135),
        .\tr[23]_i_3_1 (abus_0[22]),
        .\tr[23]_i_3_2 (sreg_n_28),
        .\tr[23]_i_6_0 (\sr_reg[8]_92 ),
        .\tr[23]_i_7_0 (sreg_n_73),
        .\tr[24]_i_10_0 (\tr[24]_i_10 ),
        .\tr[24]_i_10_1 (sreg_n_77),
        .\tr[24]_i_2 (\tr[24]_i_2 ),
        .\tr[24]_i_3_0 (sreg_n_144),
        .\tr[24]_i_3_1 (abus_0[23]),
        .\tr[24]_i_3_2 (\tr[24]_i_3 ),
        .\tr[24]_i_3_3 (sreg_n_57),
        .\tr[24]_i_3_4 (sreg_n_86),
        .\tr[24]_i_3_5 (\tr[24]_i_3_0 ),
        .\tr[25]_i_10_0 (sreg_n_124),
        .\tr[25]_i_2 (\tr[25]_i_2 ),
        .\tr[25]_i_3_0 (sreg_n_274),
        .\tr[25]_i_3_1 (abus_0[24]),
        .\tr[25]_i_3_2 (sreg_n_55),
        .\tr[25]_i_3_3 (sreg_n_467),
        .\tr[26]_i_2 (sreg_n_32),
        .\tr[26]_i_3_0 (sreg_n_448),
        .\tr[26]_i_3_1 (sreg_n_116),
        .\tr[26]_i_3_2 (abus_0[25]),
        .\tr[26]_i_3_3 (\tr[26]_i_3 ),
        .\tr[26]_i_3_4 (sreg_n_466),
        .\tr[26]_i_9_0 (\tr[26]_i_9 ),
        .\tr[27]_i_2_0 (sreg_n_31),
        .\tr[27]_i_3_0 (sreg_n_451),
        .\tr[27]_i_3_1 (abus_0[26]),
        .\tr[27]_i_3_2 (sreg_n_99),
        .\tr[27]_i_6_0 (sreg_n_134),
        .\tr[28]_i_2_0 (sreg_n_30),
        .\tr[28]_i_2_1 (\tr[28]_i_2 ),
        .\tr[28]_i_3_0 (abus_0[27]),
        .\tr[28]_i_6_0 (\sr_reg[8]_82 ),
        .\tr[29]_i_3_0 (sreg_n_469),
        .\tr[29]_i_3_1 (abus_0[28]),
        .\tr[29]_i_3_2 (sreg_n_62),
        .\tr[29]_i_3_3 (\tr[29]_i_3 ),
        .\tr[29]_i_8_0 (\sr_reg[8]_108 ),
        .\tr[30]_i_10_0 (\tr[30]_i_10 ),
        .\tr[30]_i_3_0 (sreg_n_445),
        .\tr[30]_i_3_1 (abus_0[29]),
        .\tr[30]_i_3_2 (sreg_n_94),
        .\tr[30]_i_3_3 (\tr[30]_i_3_0 ),
        .\tr[30]_i_3_4 (\tr[30]_i_3 ),
        .\tr[30]_i_9_0 (\sr_reg[8]_109 ),
        .\tr_reg[0] (\tr_reg[5] [0]),
        .\tr_reg[16] (sreg_n_70),
        .\tr_reg[19] (sreg_n_218),
        .\tr_reg[19]_0 (\tr_reg[19]_0 ),
        .\tr_reg[1] (\tr_reg[1] ),
        .\tr_reg[1]_0 (\tr_reg[1]_0 ),
        .\tr_reg[21] (sreg_n_219),
        .\tr_reg[21]_0 (\tr_reg[21]_0 ),
        .\tr_reg[23] (sreg_n_220),
        .\tr_reg[23]_0 (\tr_reg[23]_0 ),
        .\tr_reg[27] (\tr_reg[27]_0 ),
        .\tr_reg[27]_0 (sreg_n_221),
        .\tr_reg[27]_1 (\tr_reg[27]_1 ),
        .\tr_reg[28] (sreg_n_222),
        .\tr_reg[28]_0 (\tr_reg[28]_0 ),
        .\tr_reg[29] (sreg_n_223),
        .\tr_reg[29]_0 (\tr_reg[29]_0 ),
        .\tr_reg[5] (\tr_reg[5] [1]));
  niho_rgf_bank_0 bank13
       (.E(sreg_n_281),
        .SR(p_0_in),
        .abus_sel_0(abus_sel_0),
        .\badr[16]_INST_0_i_1 (sreg_n_429),
        .\badr[16]_INST_0_i_1_0 (sreg_n_413),
        .\badr[17]_INST_0_i_1 (sreg_n_430),
        .\badr[17]_INST_0_i_1_0 (sreg_n_414),
        .\badr[18]_INST_0_i_1 (sreg_n_431),
        .\badr[18]_INST_0_i_1_0 (sreg_n_415),
        .\badr[19]_INST_0_i_1 (sreg_n_432),
        .\badr[19]_INST_0_i_1_0 (sreg_n_416),
        .\badr[20]_INST_0_i_1 (sreg_n_433),
        .\badr[20]_INST_0_i_1_0 (sreg_n_417),
        .\badr[21]_INST_0_i_1 (sreg_n_434),
        .\badr[21]_INST_0_i_1_0 (sreg_n_418),
        .\badr[22]_INST_0_i_1 (sreg_n_435),
        .\badr[22]_INST_0_i_1_0 (sreg_n_419),
        .\badr[23]_INST_0_i_1 (sreg_n_436),
        .\badr[23]_INST_0_i_1_0 (sreg_n_420),
        .\badr[24]_INST_0_i_1 (sreg_n_437),
        .\badr[24]_INST_0_i_1_0 (sreg_n_421),
        .\badr[25]_INST_0_i_1 (sreg_n_438),
        .\badr[25]_INST_0_i_1_0 (sreg_n_422),
        .\badr[26]_INST_0_i_1 (sreg_n_439),
        .\badr[26]_INST_0_i_1_0 (sreg_n_423),
        .\badr[27]_INST_0_i_1 (sreg_n_440),
        .\badr[27]_INST_0_i_1_0 (sreg_n_424),
        .\badr[28]_INST_0_i_1 (sreg_n_441),
        .\badr[28]_INST_0_i_1_0 (sreg_n_425),
        .\badr[29]_INST_0_i_1 (sreg_n_442),
        .\badr[29]_INST_0_i_1_0 (sreg_n_426),
        .\badr[30]_INST_0_i_1 (sreg_n_443),
        .\badr[30]_INST_0_i_1_0 (sreg_n_427),
        .\badr[31]_INST_0_i_1 (sreg_n_444),
        .\badr[31]_INST_0_i_1_0 (sreg_n_428),
        .bbus_sel_0({bbus_sel_0[7],bbus_sel_0[4:0]}),
        .\bdatw[16]_INST_0_i_3 (sreg_n_380),
        .\bdatw[16]_INST_0_i_3_0 (sreg_n_364),
        .\bdatw[17]_INST_0_i_3 (sreg_n_379),
        .\bdatw[17]_INST_0_i_3_0 (sreg_n_363),
        .\bdatw[18]_INST_0_i_3 (sreg_n_378),
        .\bdatw[18]_INST_0_i_3_0 (sreg_n_362),
        .\bdatw[19]_INST_0_i_3 (sreg_n_377),
        .\bdatw[19]_INST_0_i_3_0 (sreg_n_361),
        .\bdatw[20]_INST_0_i_3 (sreg_n_376),
        .\bdatw[20]_INST_0_i_3_0 (sreg_n_360),
        .\bdatw[21]_INST_0_i_3 (sreg_n_375),
        .\bdatw[21]_INST_0_i_3_0 (sreg_n_359),
        .\bdatw[22]_INST_0_i_3 (sreg_n_374),
        .\bdatw[22]_INST_0_i_3_0 (sreg_n_358),
        .\bdatw[23]_INST_0_i_3 (sreg_n_373),
        .\bdatw[23]_INST_0_i_3_0 (sreg_n_357),
        .\bdatw[24]_INST_0_i_3 (sreg_n_372),
        .\bdatw[24]_INST_0_i_3_0 (sreg_n_356),
        .\bdatw[25]_INST_0_i_3 (sreg_n_371),
        .\bdatw[25]_INST_0_i_3_0 (sreg_n_355),
        .\bdatw[26]_INST_0_i_3 (sreg_n_370),
        .\bdatw[26]_INST_0_i_3_0 (sreg_n_354),
        .\bdatw[27]_INST_0_i_3 (sreg_n_369),
        .\bdatw[27]_INST_0_i_3_0 (sreg_n_353),
        .\bdatw[28]_INST_0_i_3 (sreg_n_368),
        .\bdatw[28]_INST_0_i_3_0 (sreg_n_352),
        .\bdatw[29]_INST_0_i_3 (sreg_n_367),
        .\bdatw[29]_INST_0_i_3_0 (sreg_n_351),
        .\bdatw[30]_INST_0_i_3 (sreg_n_366),
        .\bdatw[30]_INST_0_i_3_0 (sreg_n_350),
        .\bdatw[31]_INST_0_i_5 (sreg_n_365),
        .\bdatw[31]_INST_0_i_5_0 (sreg_n_349),
        .cbus(cbus[15:0]),
        .clk(clk),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .\grn_reg[0] (bank13_n_80),
        .\grn_reg[0]_0 (bank13_n_96),
        .\grn_reg[0]_1 (bank13_n_112),
        .\grn_reg[0]_10 (bank13_n_236),
        .\grn_reg[0]_11 (sreg_n_19),
        .\grn_reg[0]_12 (sreg_n_283),
        .\grn_reg[0]_13 (sreg_n_17),
        .\grn_reg[0]_2 (bank13_n_118),
        .\grn_reg[0]_3 (bank13_n_134),
        .\grn_reg[0]_4 (bank13_n_150),
        .\grn_reg[0]_5 (bank13_n_166),
        .\grn_reg[0]_6 (bank13_n_172),
        .\grn_reg[0]_7 (bank13_n_188),
        .\grn_reg[0]_8 (bank13_n_204),
        .\grn_reg[0]_9 (bank13_n_220),
        .\grn_reg[10] (bank13_n_70),
        .\grn_reg[10]_0 (bank13_n_86),
        .\grn_reg[10]_1 (bank13_n_102),
        .\grn_reg[10]_2 (bank13_n_124),
        .\grn_reg[10]_3 (bank13_n_140),
        .\grn_reg[10]_4 (bank13_n_156),
        .\grn_reg[10]_5 (bank13_n_178),
        .\grn_reg[10]_6 (bank13_n_194),
        .\grn_reg[10]_7 (bank13_n_210),
        .\grn_reg[10]_8 (bank13_n_226),
        .\grn_reg[11] (bank13_n_69),
        .\grn_reg[11]_0 (bank13_n_85),
        .\grn_reg[11]_1 (bank13_n_101),
        .\grn_reg[11]_2 (bank13_n_123),
        .\grn_reg[11]_3 (bank13_n_139),
        .\grn_reg[11]_4 (bank13_n_155),
        .\grn_reg[11]_5 (bank13_n_177),
        .\grn_reg[11]_6 (bank13_n_193),
        .\grn_reg[11]_7 (bank13_n_209),
        .\grn_reg[11]_8 (bank13_n_225),
        .\grn_reg[12] (bank13_n_68),
        .\grn_reg[12]_0 (bank13_n_84),
        .\grn_reg[12]_1 (bank13_n_100),
        .\grn_reg[12]_2 (bank13_n_122),
        .\grn_reg[12]_3 (bank13_n_138),
        .\grn_reg[12]_4 (bank13_n_154),
        .\grn_reg[12]_5 (bank13_n_176),
        .\grn_reg[12]_6 (bank13_n_192),
        .\grn_reg[12]_7 (bank13_n_208),
        .\grn_reg[12]_8 (bank13_n_224),
        .\grn_reg[13] (bank13_n_67),
        .\grn_reg[13]_0 (bank13_n_83),
        .\grn_reg[13]_1 (bank13_n_99),
        .\grn_reg[13]_2 (bank13_n_121),
        .\grn_reg[13]_3 (bank13_n_137),
        .\grn_reg[13]_4 (bank13_n_153),
        .\grn_reg[13]_5 (bank13_n_175),
        .\grn_reg[13]_6 (bank13_n_191),
        .\grn_reg[13]_7 (bank13_n_207),
        .\grn_reg[13]_8 (bank13_n_223),
        .\grn_reg[14] (bank13_n_66),
        .\grn_reg[14]_0 (bank13_n_82),
        .\grn_reg[14]_1 (bank13_n_98),
        .\grn_reg[14]_2 (bank13_n_120),
        .\grn_reg[14]_3 (bank13_n_136),
        .\grn_reg[14]_4 (bank13_n_152),
        .\grn_reg[14]_5 (bank13_n_174),
        .\grn_reg[14]_6 (bank13_n_190),
        .\grn_reg[14]_7 (bank13_n_206),
        .\grn_reg[14]_8 (bank13_n_222),
        .\grn_reg[15] ({bank13_n_16,bank13_n_17,bank13_n_18,bank13_n_19,bank13_n_20,bank13_n_21,bank13_n_22,bank13_n_23,bank13_n_24,bank13_n_25,bank13_n_26,bank13_n_27,bank13_n_28,bank13_n_29,bank13_n_30,bank13_n_31}),
        .\grn_reg[15]_0 ({bank13_n_32,bank13_n_33,bank13_n_34,bank13_n_35,bank13_n_36,bank13_n_37,bank13_n_38,bank13_n_39,bank13_n_40,bank13_n_41,bank13_n_42,bank13_n_43,bank13_n_44,bank13_n_45,bank13_n_46,bank13_n_47}),
        .\grn_reg[15]_1 ({bank13_n_48,bank13_n_49,bank13_n_50,bank13_n_51,bank13_n_52,bank13_n_53,bank13_n_54,bank13_n_55,bank13_n_56,bank13_n_57,bank13_n_58,bank13_n_59,bank13_n_60,bank13_n_61,bank13_n_62,bank13_n_63}),
        .\grn_reg[15]_10 (bank13_n_205),
        .\grn_reg[15]_11 (bank13_n_221),
        .\grn_reg[15]_12 (\grn_reg[15]_11 ),
        .\grn_reg[15]_13 (\grn_reg[15]_12 ),
        .\grn_reg[15]_14 (\grn_reg[15]_13 ),
        .\grn_reg[15]_15 (\grn_reg[15]_14 ),
        .\grn_reg[15]_16 (\grn_reg[15]_15 ),
        .\grn_reg[15]_17 (\grn_reg[15]_16 ),
        .\grn_reg[15]_18 (\grn_reg[15]_17 ),
        .\grn_reg[15]_19 (\grn_reg[15]_5 ),
        .\grn_reg[15]_2 (bank13_n_65),
        .\grn_reg[15]_20 (\grn_reg[15]_18 ),
        .\grn_reg[15]_21 (\grn_reg[15]_19 ),
        .\grn_reg[15]_22 (\grn_reg[15]_20 ),
        .\grn_reg[15]_23 (\grn_reg[15]_21 ),
        .\grn_reg[15]_24 (\grn_reg[15]_22 ),
        .\grn_reg[15]_3 (bank13_n_81),
        .\grn_reg[15]_4 (bank13_n_97),
        .\grn_reg[15]_5 (bank13_n_119),
        .\grn_reg[15]_6 (bank13_n_135),
        .\grn_reg[15]_7 (bank13_n_151),
        .\grn_reg[15]_8 (bank13_n_173),
        .\grn_reg[15]_9 (bank13_n_189),
        .\grn_reg[1] (bank13_n_79),
        .\grn_reg[1]_0 (bank13_n_95),
        .\grn_reg[1]_1 (bank13_n_111),
        .\grn_reg[1]_10 (bank13_n_235),
        .\grn_reg[1]_2 (bank13_n_117),
        .\grn_reg[1]_3 (bank13_n_133),
        .\grn_reg[1]_4 (bank13_n_149),
        .\grn_reg[1]_5 (bank13_n_165),
        .\grn_reg[1]_6 (bank13_n_171),
        .\grn_reg[1]_7 (bank13_n_187),
        .\grn_reg[1]_8 (bank13_n_203),
        .\grn_reg[1]_9 (bank13_n_219),
        .\grn_reg[2] (bank13_n_78),
        .\grn_reg[2]_0 (bank13_n_94),
        .\grn_reg[2]_1 (bank13_n_110),
        .\grn_reg[2]_10 (bank13_n_234),
        .\grn_reg[2]_2 (bank13_n_116),
        .\grn_reg[2]_3 (bank13_n_132),
        .\grn_reg[2]_4 (bank13_n_148),
        .\grn_reg[2]_5 (bank13_n_164),
        .\grn_reg[2]_6 (bank13_n_170),
        .\grn_reg[2]_7 (bank13_n_186),
        .\grn_reg[2]_8 (bank13_n_202),
        .\grn_reg[2]_9 (bank13_n_218),
        .\grn_reg[3] (bank13_n_77),
        .\grn_reg[3]_0 (bank13_n_93),
        .\grn_reg[3]_1 (bank13_n_109),
        .\grn_reg[3]_10 (bank13_n_233),
        .\grn_reg[3]_2 (bank13_n_115),
        .\grn_reg[3]_3 (bank13_n_131),
        .\grn_reg[3]_4 (bank13_n_147),
        .\grn_reg[3]_5 (bank13_n_163),
        .\grn_reg[3]_6 (bank13_n_169),
        .\grn_reg[3]_7 (bank13_n_185),
        .\grn_reg[3]_8 (bank13_n_201),
        .\grn_reg[3]_9 (bank13_n_217),
        .\grn_reg[4] (bank13_n_76),
        .\grn_reg[4]_0 (bank13_n_92),
        .\grn_reg[4]_1 (bank13_n_108),
        .\grn_reg[4]_10 (bank13_n_232),
        .\grn_reg[4]_2 (bank13_n_114),
        .\grn_reg[4]_3 (bank13_n_130),
        .\grn_reg[4]_4 (bank13_n_146),
        .\grn_reg[4]_5 (bank13_n_162),
        .\grn_reg[4]_6 (bank13_n_168),
        .\grn_reg[4]_7 (bank13_n_184),
        .\grn_reg[4]_8 (bank13_n_200),
        .\grn_reg[4]_9 (bank13_n_216),
        .\grn_reg[5] (bank13_n_75),
        .\grn_reg[5]_0 (bank13_n_91),
        .\grn_reg[5]_1 (bank13_n_107),
        .\grn_reg[5]_10 (bank13_n_231),
        .\grn_reg[5]_2 (bank13_n_113),
        .\grn_reg[5]_3 (bank13_n_129),
        .\grn_reg[5]_4 (bank13_n_145),
        .\grn_reg[5]_5 (bank13_n_161),
        .\grn_reg[5]_6 (bank13_n_167),
        .\grn_reg[5]_7 (bank13_n_183),
        .\grn_reg[5]_8 (bank13_n_199),
        .\grn_reg[5]_9 (bank13_n_215),
        .\grn_reg[6] (bank13_n_74),
        .\grn_reg[6]_0 (bank13_n_90),
        .\grn_reg[6]_1 (bank13_n_106),
        .\grn_reg[6]_2 (bank13_n_128),
        .\grn_reg[6]_3 (bank13_n_144),
        .\grn_reg[6]_4 (bank13_n_160),
        .\grn_reg[6]_5 (bank13_n_182),
        .\grn_reg[6]_6 (bank13_n_198),
        .\grn_reg[6]_7 (bank13_n_214),
        .\grn_reg[6]_8 (bank13_n_230),
        .\grn_reg[7] (bank13_n_73),
        .\grn_reg[7]_0 (bank13_n_89),
        .\grn_reg[7]_1 (bank13_n_105),
        .\grn_reg[7]_2 (bank13_n_127),
        .\grn_reg[7]_3 (bank13_n_143),
        .\grn_reg[7]_4 (bank13_n_159),
        .\grn_reg[7]_5 (bank13_n_181),
        .\grn_reg[7]_6 (bank13_n_197),
        .\grn_reg[7]_7 (bank13_n_213),
        .\grn_reg[7]_8 (bank13_n_229),
        .\grn_reg[8] (bank13_n_72),
        .\grn_reg[8]_0 (bank13_n_88),
        .\grn_reg[8]_1 (bank13_n_104),
        .\grn_reg[8]_2 (bank13_n_126),
        .\grn_reg[8]_3 (bank13_n_142),
        .\grn_reg[8]_4 (bank13_n_158),
        .\grn_reg[8]_5 (bank13_n_180),
        .\grn_reg[8]_6 (bank13_n_196),
        .\grn_reg[8]_7 (bank13_n_212),
        .\grn_reg[8]_8 (bank13_n_228),
        .\grn_reg[9] (bank13_n_71),
        .\grn_reg[9]_0 (bank13_n_87),
        .\grn_reg[9]_1 (bank13_n_103),
        .\grn_reg[9]_2 (bank13_n_125),
        .\grn_reg[9]_3 (bank13_n_141),
        .\grn_reg[9]_4 (bank13_n_157),
        .\grn_reg[9]_5 (bank13_n_179),
        .\grn_reg[9]_6 (bank13_n_195),
        .\grn_reg[9]_7 (bank13_n_211),
        .\grn_reg[9]_8 (bank13_n_227),
        .\i_/badr[15]_INST_0_i_17 (sreg_n_275),
        .\i_/badr[15]_INST_0_i_19 (sreg_n_280),
        .\i_/badr[15]_INST_0_i_20 ({out[8],out[1:0]}),
        .\i_/bdatw[15]_INST_0_i_27 (\i_/bdatw[15]_INST_0_i_27 ),
        .\i_/bdatw[15]_INST_0_i_27_0 (\i_/bdatw[15]_INST_0_i_27_0 ),
        .\i_/bdatw[15]_INST_0_i_66 (\i_/bdatw[15]_INST_0_i_65_2 ),
        .\i_/bdatw[15]_INST_0_i_66_0 (\i_/bdatw[15]_INST_0_i_65_0 ),
        .\i_/bdatw[15]_INST_0_i_66_1 (\i_/bdatw[15]_INST_0_i_65_1 ),
        .\i_/bdatw[15]_INST_0_i_66_2 (\i_/bdatw[15]_INST_0_i_65 ),
        .\i_/bdatw[15]_INST_0_i_67 (\i_/bdatw[15]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_67_0 (\i_/bdatw[15]_INST_0_i_67_0 ),
        .out({bank13_n_0,bank13_n_1,bank13_n_2,bank13_n_3,bank13_n_4,bank13_n_5,bank13_n_6,bank13_n_7,bank13_n_8,bank13_n_9,bank13_n_10,bank13_n_11,bank13_n_12,bank13_n_13,bank13_n_14,bank13_n_15}),
        .rst_n(rst_n));
  niho_rgf_bus_1 bbus_out
       (.bbus_sel_cr(bbus_sel_cr),
        .bbus_sr(bbus_sr),
        .\bdatw[15]_INST_0_i_9_0 (rgf_pc),
        .\bdatw[16]_INST_0_i_1 (bank13_n_236),
        .\bdatw[16]_INST_0_i_1_0 (bank13_n_220),
        .\bdatw[16]_INST_0_i_1_1 (sreg_n_300),
        .\bdatw[16]_INST_0_i_1_2 (sreg_n_316),
        .\bdatw[16]_INST_0_i_1_3 (sreg_n_332),
        .\bdatw[16]_INST_0_i_1_4 (sreg_n_348),
        .\bdatw[17]_INST_0_i_1 (bank13_n_235),
        .\bdatw[17]_INST_0_i_1_0 (bank13_n_219),
        .\bdatw[17]_INST_0_i_1_1 (sreg_n_299),
        .\bdatw[17]_INST_0_i_1_2 (sreg_n_315),
        .\bdatw[17]_INST_0_i_1_3 (sreg_n_331),
        .\bdatw[17]_INST_0_i_1_4 (sreg_n_347),
        .\bdatw[18]_INST_0_i_1 (bank13_n_234),
        .\bdatw[18]_INST_0_i_1_0 (bank13_n_218),
        .\bdatw[18]_INST_0_i_1_1 (sreg_n_298),
        .\bdatw[18]_INST_0_i_1_2 (sreg_n_314),
        .\bdatw[18]_INST_0_i_1_3 (sreg_n_330),
        .\bdatw[18]_INST_0_i_1_4 (sreg_n_346),
        .\bdatw[19]_INST_0_i_1 (bank13_n_233),
        .\bdatw[19]_INST_0_i_1_0 (bank13_n_217),
        .\bdatw[19]_INST_0_i_1_1 (sreg_n_297),
        .\bdatw[19]_INST_0_i_1_2 (sreg_n_313),
        .\bdatw[19]_INST_0_i_1_3 (sreg_n_329),
        .\bdatw[19]_INST_0_i_1_4 (sreg_n_345),
        .\bdatw[20]_INST_0_i_1 (bank13_n_232),
        .\bdatw[20]_INST_0_i_1_0 (bank13_n_216),
        .\bdatw[20]_INST_0_i_1_1 (sreg_n_296),
        .\bdatw[20]_INST_0_i_1_2 (sreg_n_312),
        .\bdatw[20]_INST_0_i_1_3 (sreg_n_328),
        .\bdatw[20]_INST_0_i_1_4 (sreg_n_344),
        .\bdatw[21]_INST_0_i_1 (bank13_n_231),
        .\bdatw[21]_INST_0_i_1_0 (bank13_n_215),
        .\bdatw[21]_INST_0_i_1_1 (sreg_n_295),
        .\bdatw[21]_INST_0_i_1_2 (sreg_n_311),
        .\bdatw[21]_INST_0_i_1_3 (sreg_n_327),
        .\bdatw[21]_INST_0_i_1_4 (sreg_n_343),
        .\bdatw[22]_INST_0_i_1 (bank13_n_230),
        .\bdatw[22]_INST_0_i_1_0 (bank13_n_214),
        .\bdatw[22]_INST_0_i_1_1 (sreg_n_294),
        .\bdatw[22]_INST_0_i_1_2 (sreg_n_310),
        .\bdatw[22]_INST_0_i_1_3 (sreg_n_326),
        .\bdatw[22]_INST_0_i_1_4 (sreg_n_342),
        .\bdatw[23]_INST_0_i_1 (bank13_n_229),
        .\bdatw[23]_INST_0_i_1_0 (bank13_n_213),
        .\bdatw[23]_INST_0_i_1_1 (sreg_n_293),
        .\bdatw[23]_INST_0_i_1_2 (sreg_n_309),
        .\bdatw[23]_INST_0_i_1_3 (sreg_n_325),
        .\bdatw[23]_INST_0_i_1_4 (sreg_n_341),
        .\bdatw[24]_INST_0_i_1 (bank13_n_228),
        .\bdatw[24]_INST_0_i_1_0 (bank13_n_212),
        .\bdatw[24]_INST_0_i_1_1 (sreg_n_292),
        .\bdatw[24]_INST_0_i_1_2 (sreg_n_308),
        .\bdatw[24]_INST_0_i_1_3 (sreg_n_324),
        .\bdatw[24]_INST_0_i_1_4 (sreg_n_340),
        .\bdatw[25]_INST_0_i_1 (bank13_n_227),
        .\bdatw[25]_INST_0_i_1_0 (bank13_n_211),
        .\bdatw[25]_INST_0_i_1_1 (sreg_n_291),
        .\bdatw[25]_INST_0_i_1_2 (sreg_n_307),
        .\bdatw[25]_INST_0_i_1_3 (sreg_n_323),
        .\bdatw[25]_INST_0_i_1_4 (sreg_n_339),
        .\bdatw[26]_INST_0_i_1 (bank13_n_226),
        .\bdatw[26]_INST_0_i_1_0 (bank13_n_210),
        .\bdatw[26]_INST_0_i_1_1 (sreg_n_290),
        .\bdatw[26]_INST_0_i_1_2 (sreg_n_306),
        .\bdatw[26]_INST_0_i_1_3 (sreg_n_322),
        .\bdatw[26]_INST_0_i_1_4 (sreg_n_338),
        .\bdatw[27]_INST_0_i_1 (bank13_n_225),
        .\bdatw[27]_INST_0_i_1_0 (bank13_n_209),
        .\bdatw[27]_INST_0_i_1_1 (sreg_n_289),
        .\bdatw[27]_INST_0_i_1_2 (sreg_n_305),
        .\bdatw[27]_INST_0_i_1_3 (sreg_n_321),
        .\bdatw[27]_INST_0_i_1_4 (sreg_n_337),
        .\bdatw[28]_INST_0_i_1 (bank13_n_224),
        .\bdatw[28]_INST_0_i_1_0 (bank13_n_208),
        .\bdatw[28]_INST_0_i_1_1 (sreg_n_288),
        .\bdatw[28]_INST_0_i_1_2 (sreg_n_304),
        .\bdatw[28]_INST_0_i_1_3 (sreg_n_320),
        .\bdatw[28]_INST_0_i_1_4 (sreg_n_336),
        .\bdatw[29]_INST_0_i_1 (bank13_n_223),
        .\bdatw[29]_INST_0_i_1_0 (bank13_n_207),
        .\bdatw[29]_INST_0_i_1_1 (sreg_n_287),
        .\bdatw[29]_INST_0_i_1_2 (sreg_n_303),
        .\bdatw[29]_INST_0_i_1_3 (sreg_n_319),
        .\bdatw[29]_INST_0_i_1_4 (sreg_n_335),
        .\bdatw[30]_INST_0_i_1 (bank13_n_222),
        .\bdatw[30]_INST_0_i_1_0 (bank13_n_206),
        .\bdatw[30]_INST_0_i_1_1 (sreg_n_286),
        .\bdatw[30]_INST_0_i_1_2 (sreg_n_302),
        .\bdatw[30]_INST_0_i_1_3 (sreg_n_318),
        .\bdatw[30]_INST_0_i_1_4 (sreg_n_334),
        .\bdatw[31]_INST_0_i_1 (\tr_reg[31] ),
        .\bdatw[31]_INST_0_i_1_0 ({p_0_in_1,\sp_reg[0] }),
        .\bdatw[31]_INST_0_i_1_1 (bank13_n_221),
        .\bdatw[31]_INST_0_i_1_2 (bank13_n_205),
        .\bdatw[31]_INST_0_i_1_3 (sreg_n_285),
        .\bdatw[31]_INST_0_i_1_4 (sreg_n_301),
        .\bdatw[31]_INST_0_i_1_5 (sreg_n_317),
        .\bdatw[31]_INST_0_i_1_6 (sreg_n_333),
        .\grn_reg[0] (bbus_out_n_16),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[5] (bbus_out_n_10),
        .\iv[12]_i_51 (bank02_n_452),
        .\iv[12]_i_51_0 (bank02_n_458),
        .\iv[12]_i_51_1 (bank02_n_430),
        .\iv[12]_i_51_2 (bank02_n_436),
        .\iv[15]_i_56 (bank02_n_447),
        .\iv[15]_i_56_0 (bank02_n_453),
        .\iv[15]_i_56_1 (bank02_n_425),
        .\iv[15]_i_56_2 (bank02_n_431),
        .\iv_reg[10] (\iv_reg[10] ),
        .\iv_reg[11] (\iv_reg[11] ),
        .\iv_reg[12] (\iv_reg[12] ),
        .\iv_reg[13] (\iv_reg[13] ),
        .\iv_reg[14] (\iv_reg[14] ),
        .\iv_reg[15] (\iv_reg[15] ),
        .\iv_reg[6] (\iv_reg[6] ),
        .\iv_reg[7] (\iv_reg[7] ),
        .\iv_reg[8] (\iv_reg[8] ),
        .\iv_reg[9] (\iv_reg[9] ),
        .\mul_b_reg[0] (bank13_n_112),
        .\mul_b_reg[0]_0 (bank13_n_118),
        .\mul_b_reg[0]_1 (bank13_n_172),
        .\mul_b_reg[0]_2 (bank13_n_166),
        .\mul_b_reg[10] (bank02_n_442),
        .\mul_b_reg[10]_0 (bank02_n_420),
        .\mul_b_reg[10]_1 (bank13_n_102),
        .\mul_b_reg[10]_2 (bank13_n_156),
        .\mul_b_reg[11] (bank02_n_441),
        .\mul_b_reg[11]_0 (bank02_n_419),
        .\mul_b_reg[11]_1 (bank13_n_101),
        .\mul_b_reg[11]_2 (bank13_n_155),
        .\mul_b_reg[12] (bank02_n_440),
        .\mul_b_reg[12]_0 (bank02_n_418),
        .\mul_b_reg[12]_1 (bank13_n_100),
        .\mul_b_reg[12]_2 (bank13_n_154),
        .\mul_b_reg[13] (bank02_n_439),
        .\mul_b_reg[13]_0 (bank02_n_417),
        .\mul_b_reg[13]_1 (bank13_n_99),
        .\mul_b_reg[13]_2 (bank13_n_153),
        .\mul_b_reg[14] (bank02_n_438),
        .\mul_b_reg[14]_0 (bank02_n_416),
        .\mul_b_reg[14]_1 (bank13_n_98),
        .\mul_b_reg[14]_2 (bank13_n_152),
        .\mul_b_reg[15] (bank02_n_437),
        .\mul_b_reg[15]_0 (bank02_n_415),
        .\mul_b_reg[15]_1 (\iv_reg[15]_0 ),
        .\mul_b_reg[15]_2 (bank13_n_97),
        .\mul_b_reg[15]_3 (bank13_n_151),
        .\mul_b_reg[1] (bank02_n_451),
        .\mul_b_reg[1]_0 (bank02_n_457),
        .\mul_b_reg[1]_1 (bank02_n_429),
        .\mul_b_reg[1]_2 (bank02_n_435),
        .\mul_b_reg[1]_3 (bank13_n_165),
        .\mul_b_reg[1]_4 (bank13_n_171),
        .\mul_b_reg[1]_5 (bank13_n_117),
        .\mul_b_reg[1]_6 (bank13_n_111),
        .\mul_b_reg[2] (bank02_n_450),
        .\mul_b_reg[2]_0 (bank02_n_456),
        .\mul_b_reg[2]_1 (bank02_n_428),
        .\mul_b_reg[2]_2 (bank02_n_434),
        .\mul_b_reg[2]_3 (bank13_n_164),
        .\mul_b_reg[2]_4 (bank13_n_170),
        .\mul_b_reg[2]_5 (bank13_n_116),
        .\mul_b_reg[2]_6 (bank13_n_110),
        .\mul_b_reg[3] (bank02_n_449),
        .\mul_b_reg[3]_0 (bank02_n_455),
        .\mul_b_reg[3]_1 (bank02_n_427),
        .\mul_b_reg[3]_2 (bank02_n_433),
        .\mul_b_reg[3]_3 (bank13_n_163),
        .\mul_b_reg[3]_4 (bank13_n_169),
        .\mul_b_reg[3]_5 (bank13_n_115),
        .\mul_b_reg[3]_6 (bank13_n_109),
        .\mul_b_reg[4] (bank02_n_448),
        .\mul_b_reg[4]_0 (bank02_n_454),
        .\mul_b_reg[4]_1 (bank02_n_426),
        .\mul_b_reg[4]_2 (bank02_n_432),
        .\mul_b_reg[4]_3 (bank13_n_162),
        .\mul_b_reg[4]_4 (bank13_n_168),
        .\mul_b_reg[4]_5 (bank13_n_114),
        .\mul_b_reg[4]_6 (bank13_n_108),
        .\mul_b_reg[5] (bank13_n_107),
        .\mul_b_reg[5]_0 (bank13_n_113),
        .\mul_b_reg[5]_1 (bank13_n_167),
        .\mul_b_reg[5]_2 (bank13_n_161),
        .\mul_b_reg[6] (bank02_n_446),
        .\mul_b_reg[6]_0 (bank02_n_424),
        .\mul_b_reg[6]_1 (bank13_n_106),
        .\mul_b_reg[6]_2 (bank13_n_160),
        .\mul_b_reg[7] (bank02_n_445),
        .\mul_b_reg[7]_0 (bank02_n_423),
        .\mul_b_reg[7]_1 (bank13_n_105),
        .\mul_b_reg[7]_2 (bank13_n_159),
        .\mul_b_reg[8] (bank02_n_444),
        .\mul_b_reg[8]_0 (bank02_n_422),
        .\mul_b_reg[8]_1 (bank13_n_104),
        .\mul_b_reg[8]_2 (bank13_n_158),
        .\mul_b_reg[9] (bank02_n_443),
        .\mul_b_reg[9]_0 (bank02_n_421),
        .\mul_b_reg[9]_1 (bank13_n_103),
        .\mul_b_reg[9]_2 (bank13_n_157),
        .out({p_0_in_2[15:14],out[12:9],p_0_in_2[9],out[8:1]}),
        .sp_dec_0(sp_dec_0),
        .\sp_reg[0] (bbus_out_n_35),
        .\sp_reg[16] (\sp_reg[16]_0 ),
        .\sp_reg[17] (\sp_reg[17]_0 ),
        .\sp_reg[18] (\sp_reg[18]_0 ),
        .\sp_reg[19] (\sp_reg[19]_0 ),
        .\sp_reg[1] (\sp_reg[1]_0 ),
        .\sp_reg[20] (\sp_reg[20]_0 ),
        .\sp_reg[21] (\sp_reg[21]_0 ),
        .\sp_reg[22] (\sp_reg[22]_0 ),
        .\sp_reg[23] (\sp_reg[23]_0 ),
        .\sp_reg[24] (\sp_reg[24]_0 ),
        .\sp_reg[25] (\sp_reg[25]_0 ),
        .\sp_reg[26] (\sp_reg[26]_0 ),
        .\sp_reg[27] (\sp_reg[27]_0 ),
        .\sp_reg[28] (\sp_reg[28]_0 ),
        .\sp_reg[29] (\sp_reg[29]_0 ),
        .\sp_reg[2] (\sp_reg[2]_0 ),
        .\sp_reg[30] (\sp_reg[30]_0 ),
        .\sp_reg[31] (\sp_reg[31]_0 ),
        .\sp_reg[3] (\sp_reg[3]_0 ),
        .\sp_reg[4] (\sp_reg[4]_0 ),
        .\sp_reg[5] (bbus_out_n_28),
        .\sp_reg[5]_0 (bbus_out_n_29),
        .\sr_reg[10] (\sr_reg[10] ),
        .\sr_reg[11] (\sr_reg[11] ),
        .\sr_reg[12] (\sr_reg[12] ),
        .\sr_reg[13] (\sr_reg[13] ),
        .\sr_reg[14] (\sr_reg[14] ),
        .\sr_reg[15] (\sr_reg[15] ),
        .\sr_reg[1] (\sr_reg[1] ),
        .\sr_reg[2] (\sr_reg[2] ),
        .\sr_reg[3] (\sr_reg[3] ),
        .\sr_reg[4] (\sr_reg[4] ),
        .\sr_reg[5] (bbus_out_n_30),
        .\sr_reg[6] (\sr_reg[6]_9 ),
        .\sr_reg[7] (\sr_reg[7]_3 ),
        .\sr_reg[8] (\sr_reg[8]_168 ),
        .\sr_reg[9] (\sr_reg[9] ),
        .\tr_reg[0] (bbus_out_n_17),
        .\tr_reg[16] (\tr_reg[16] ),
        .\tr_reg[17] (\tr_reg[17] ),
        .\tr_reg[18] (\tr_reg[18] ),
        .\tr_reg[19] (\tr_reg[19] ),
        .\tr_reg[20] (\tr_reg[20] ),
        .\tr_reg[21] (\tr_reg[21] ),
        .\tr_reg[22] (\tr_reg[22] ),
        .\tr_reg[23] (\tr_reg[23] ),
        .\tr_reg[24] (\tr_reg[24] ),
        .\tr_reg[25] (\tr_reg[25] ),
        .\tr_reg[26] (\tr_reg[26] ),
        .\tr_reg[27] (\tr_reg[27] ),
        .\tr_reg[28] (\tr_reg[28] ),
        .\tr_reg[29] (\tr_reg[29] ),
        .\tr_reg[30] (\tr_reg[30] ),
        .\tr_reg[31] (\tr_reg[31]_0 ),
        .\tr_reg[5] (bbus_out_n_11));
  niho_rgf_ivec ivec
       (.SR(p_0_in),
        .cbus(cbus[15:0]),
        .clk(clk),
        .\iv_reg[0]_0 (\tr_reg[0] [0]),
        .\iv_reg[15]_0 (\iv_reg[15]_0 ));
  niho_rgf_pcnt pcnt
       (.S(sreg_n_261),
        .SR(p_0_in),
        .clk(clk),
        .fch_pc(fch_pc),
        .out(rgf_pc),
        .\pc_reg[15]_0 (\pc_reg[15] ));
  niho_rgf_ctl rctl
       (.bank_sel(bank_sel),
        .out({out[8],out[1:0]}));
  niho_rgf_sptr sptr
       (.O(O),
        .SR(p_0_in),
        .abus_sel_cr(abus_sel_cr[3:2]),
        .abus_sp(abus_sp),
        .clk(clk),
        .ctl_sp_dec(ctl_sp_dec),
        .ctl_sp_id4(ctl_sp_id4),
        .ctl_sp_inc(ctl_sp_inc),
        .out({p_0_in_1,\sp_reg[0] }),
        .sp_dec_0(sp_dec_0),
        .\sp_reg[10]_0 (\sp_reg[10] ),
        .\sp_reg[11]_0 (\sp_reg[11] ),
        .\sp_reg[12]_0 (\sp_reg[12] ),
        .\sp_reg[13]_0 (\sp_reg[13] ),
        .\sp_reg[14]_0 (\sp_reg[14] ),
        .\sp_reg[15]_0 (\sp_reg[15] ),
        .\sp_reg[16]_0 (\sp_reg[16] ),
        .\sp_reg[17]_0 (\sp_reg[17] ),
        .\sp_reg[18]_0 (\sp_reg[18] ),
        .\sp_reg[19]_0 (\sp_reg[19] ),
        .\sp_reg[1]_0 (\sp_reg[1] ),
        .\sp_reg[20]_0 (\sp_reg[20] ),
        .\sp_reg[21]_0 (\sp_reg[21] ),
        .\sp_reg[22]_0 (\sp_reg[22] ),
        .\sp_reg[23]_0 (\sp_reg[23] ),
        .\sp_reg[24]_0 (\sp_reg[24] ),
        .\sp_reg[25]_0 (\sp_reg[25] ),
        .\sp_reg[26]_0 (\sp_reg[26] ),
        .\sp_reg[27]_0 (\sp_reg[27] ),
        .\sp_reg[28]_0 (\sp_reg[28] ),
        .\sp_reg[29]_0 (\sp_reg[29] ),
        .\sp_reg[2]_0 (\sp_reg[2] ),
        .\sp_reg[30]_0 (\sp_reg[30] ),
        .\sp_reg[31]_0 (\sp_reg[31] ),
        .\sp_reg[31]_1 (\sp_reg[31]_1 ),
        .\sp_reg[3]_0 (\sp_reg[3] ),
        .\sp_reg[4]_0 (\sp_reg[4] ),
        .\sp_reg[5]_0 (\sp_reg[5] ),
        .\sp_reg[6]_0 (\sp_reg[6] ),
        .\sp_reg[7]_0 (\sp_reg[7] ),
        .\sp_reg[8]_0 (\sp_reg[8] ),
        .\sp_reg[9]_0 (\sp_reg[9] ));
  niho_rgf_sreg sreg
       (.CO(bank02_n_364),
        .D(D),
        .DI(abus_0[15:12]),
        .E(sreg_n_281),
        .O(\sr_reg[8]_1 ),
        .Q(Q),
        .S(sreg_n_261),
        .SR(p_0_in),
        .abus_o(abus_o[31:16]),
        .\abus_o[16] (abus_o_16_sn_1),
        .abus_sel_0({abus_sel_0[6:5],abus_sel_0[2:1]}),
        .alu_sr_flag(alu_sr_flag),
        .\badr[0]_INST_0_i_1 (\badr[0]_INST_0_i_1_0 ),
        .\badr[16]_INST_0_i_1 (sreg_n_109),
        .\badr[16]_INST_0_i_1_0 (sreg_n_145),
        .\badr[17]_INST_0_i_1 (sreg_n_151),
        .\badr[18]_INST_0_i_1 (sreg_n_128),
        .\badr[1]_INST_0_i_1 (\badr[1]_INST_0_i_1 ),
        .\badr[2]_INST_0_i_1 (\badr[2]_INST_0_i_1 ),
        .\badr[31]_INST_0_i_69 (\badr[31]_INST_0_i_69 ),
        .\badr[4]_INST_0_i_1 (\badr[4]_INST_0_i_1 ),
        .\badr[5]_INST_0_i_1 (\badr[5]_INST_0_i_1_0 ),
        .\badr[6]_INST_0_i_1 (\badr[6]_INST_0_i_1 ),
        .bbus_0(bbus_0[2:0]),
        .bbus_sel_0(bbus_sel_0),
        .\bdatw[31]_INST_0_i_4 ({bank02_n_64,bank02_n_65,bank02_n_66,bank02_n_67,bank02_n_68,bank02_n_69,bank02_n_70,bank02_n_71,bank02_n_72,bank02_n_73,bank02_n_74,bank02_n_75,bank02_n_76,bank02_n_77,bank02_n_78,bank02_n_79}),
        .\bdatw[31]_INST_0_i_4_0 ({bank02_n_48,bank02_n_49,bank02_n_50,bank02_n_51,bank02_n_52,bank02_n_53,bank02_n_54,bank02_n_55,bank02_n_56,bank02_n_57,bank02_n_58,bank02_n_59,bank02_n_60,bank02_n_61,bank02_n_62,bank02_n_63}),
        .\bdatw[31]_INST_0_i_4_1 ({bank02_n_0,bank02_n_1,bank02_n_2,bank02_n_3,bank02_n_4,bank02_n_5,bank02_n_6,bank02_n_7,bank02_n_8,bank02_n_9,bank02_n_10,bank02_n_11,bank02_n_12,bank02_n_13,bank02_n_14,bank02_n_15}),
        .\bdatw[31]_INST_0_i_4_2 ({bank02_n_112,bank02_n_113,bank02_n_114,bank02_n_115,bank02_n_116,bank02_n_117,bank02_n_118,bank02_n_119,bank02_n_120,bank02_n_121,bank02_n_122,bank02_n_123,bank02_n_124,bank02_n_125,bank02_n_126,bank02_n_127}),
        .cbus_sel_0(cbus_sel_0),
        .clk(clk),
        .fch_irq_req(fch_irq_req),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\i_/badr[31]_INST_0_i_4 ({bank02_n_96,bank02_n_97,bank02_n_98,bank02_n_99,bank02_n_100,bank02_n_101,bank02_n_102,bank02_n_103,bank02_n_104,bank02_n_105,bank02_n_106,bank02_n_107,bank02_n_108,bank02_n_109,bank02_n_110,bank02_n_111}),
        .\i_/badr[31]_INST_0_i_4_0 ({bank02_n_80,bank02_n_81,bank02_n_82,bank02_n_83,bank02_n_84,bank02_n_85,bank02_n_86,bank02_n_87,bank02_n_88,bank02_n_89,bank02_n_90,bank02_n_91,bank02_n_92,bank02_n_93,bank02_n_94,bank02_n_95}),
        .\i_/badr[31]_INST_0_i_5 ({bank02_n_32,bank02_n_33,bank02_n_34,bank02_n_35,bank02_n_36,bank02_n_37,bank02_n_38,bank02_n_39,bank02_n_40,bank02_n_41,bank02_n_42,bank02_n_43,bank02_n_44,bank02_n_45,bank02_n_46,bank02_n_47}),
        .\i_/badr[31]_INST_0_i_5_0 ({bank02_n_16,bank02_n_17,bank02_n_18,bank02_n_19,bank02_n_20,bank02_n_21,bank02_n_22,bank02_n_23,bank02_n_24,bank02_n_25,bank02_n_26,bank02_n_27,bank02_n_28,bank02_n_29,bank02_n_30,bank02_n_31}),
        .\i_/badr[31]_INST_0_i_6 ({bank13_n_48,bank13_n_49,bank13_n_50,bank13_n_51,bank13_n_52,bank13_n_53,bank13_n_54,bank13_n_55,bank13_n_56,bank13_n_57,bank13_n_58,bank13_n_59,bank13_n_60,bank13_n_61,bank13_n_62,bank13_n_63}),
        .\i_/badr[31]_INST_0_i_6_0 ({bank13_n_32,bank13_n_33,bank13_n_34,bank13_n_35,bank13_n_36,bank13_n_37,bank13_n_38,bank13_n_39,bank13_n_40,bank13_n_41,bank13_n_42,bank13_n_43,bank13_n_44,bank13_n_45,bank13_n_46,bank13_n_47}),
        .\i_/badr[31]_INST_0_i_7 ({bank13_n_16,bank13_n_17,bank13_n_18,bank13_n_19,bank13_n_20,bank13_n_21,bank13_n_22,bank13_n_23,bank13_n_24,bank13_n_25,bank13_n_26,bank13_n_27,bank13_n_28,bank13_n_29,bank13_n_30,bank13_n_31}),
        .\i_/badr[31]_INST_0_i_7_0 ({bank13_n_0,bank13_n_1,bank13_n_2,bank13_n_3,bank13_n_4,bank13_n_5,bank13_n_6,bank13_n_7,bank13_n_8,bank13_n_9,bank13_n_10,bank13_n_11,bank13_n_12,bank13_n_13,bank13_n_14,bank13_n_15}),
        .irq(irq),
        .irq_lev(irq_lev),
        .irq_lev_0_sp_1(irq_lev_0_sn_1),
        .irq_lev_1_sp_1(irq_lev_1_sn_1),
        .\iv[0]_i_21 (\iv[0]_i_10 ),
        .\iv[0]_i_3 (bank02_n_231),
        .\iv[0]_i_31_0 (sreg_n_136),
        .\iv[0]_i_3_0 (\iv[0]_i_3_0 ),
        .\iv[0]_i_3_1 (bank02_n_387),
        .\iv[10]_i_29_0 (bank02_n_272),
        .\iv[10]_i_34 (sreg_n_116),
        .\iv[10]_i_4 (bank02_n_202),
        .\iv[10]_i_41_0 (sreg_n_66),
        .\iv[10]_i_44_0 (sreg_n_117),
        .\iv[10]_i_44_1 (bbus_out_n_16),
        .\iv[10]_i_44_2 (bbus_out_n_35),
        .\iv[10]_i_6 (bank02_n_245),
        .\iv[10]_i_9 (\iv[10]_i_9 ),
        .\iv[11]_i_10_0 (\sr_reg[8]_123 ),
        .\iv[11]_i_11_0 (\iv[11]_i_11 ),
        .\iv[11]_i_4_0 (bank02_n_150),
        .\iv[12]_i_25 (\badr[0]_INST_0_i_1 ),
        .\iv[12]_i_49 (sreg_n_140),
        .\iv[12]_i_9 (bank02_n_265),
        .\iv[13]_i_10_0 (\iv[13]_i_10 ),
        .\iv[13]_i_35 (sreg_n_108),
        .\iv[13]_i_45_0 (\mul_b_reg[0] ),
        .\iv[13]_i_45_1 (\mul_b_reg[0]_0 ),
        .\iv[13]_i_4_0 (\sr_reg[8]_42 ),
        .\iv[13]_i_4_1 (\sr_reg[8]_16 ),
        .\iv[13]_i_50 (sreg_n_110),
        .\iv[14]_i_11_0 (\iv[14]_i_11 ),
        .\iv[14]_i_13 (bank02_n_264),
        .\iv[14]_i_2 (\sr_reg[8]_28 ),
        .\iv[14]_i_30_0 (sreg_n_154),
        .\iv[15]_i_108 (\iv[15]_i_108_9 ),
        .\iv[15]_i_108_0 (\iv[15]_i_108_10 ),
        .\iv[15]_i_108_1 (\iv[15]_i_108_11 ),
        .\iv[15]_i_108_10 (\iv[15]_i_108_20 ),
        .\iv[15]_i_108_11 (\iv[15]_i_108_21 ),
        .\iv[15]_i_108_12 (\iv[15]_i_108_22 ),
        .\iv[15]_i_108_13 (\iv[15]_i_108_23 ),
        .\iv[15]_i_108_2 (\iv[15]_i_108_12 ),
        .\iv[15]_i_108_3 (\iv[15]_i_108_13 ),
        .\iv[15]_i_108_4 (\iv[15]_i_108_14 ),
        .\iv[15]_i_108_5 (\iv[15]_i_108_15 ),
        .\iv[15]_i_108_6 (\iv[15]_i_108_16 ),
        .\iv[15]_i_108_7 (\iv[15]_i_108_17 ),
        .\iv[15]_i_108_8 (\iv[15]_i_108_18 ),
        .\iv[15]_i_108_9 (\iv[15]_i_108_19 ),
        .\iv[15]_i_58 (bank02_n_284),
        .\iv[15]_i_8 (bank02_n_253),
        .\iv[15]_i_8_0 (bank02_n_252),
        .\iv[15]_i_8_1 (\iv[15]_i_8_2 ),
        .\iv[15]_i_8_2 (bank02_n_214),
        .\iv[15]_i_96 (bbus_out_n_29),
        .\iv[15]_i_96_0 (bbus_out_n_30),
        .\iv[15]_i_96_1 (bbus_out_n_10),
        .\iv[15]_i_96_2 (\mul_b_reg[5] ),
        .\iv[15]_i_96_3 (\mul_b_reg[5]_0 ),
        .\iv[15]_i_96_4 (\iv[15]_i_96 ),
        .\iv[15]_i_96_5 (\sp_reg[4]_0 ),
        .\iv[15]_i_96_6 (\sr_reg[4] ),
        .\iv[15]_i_96_7 (\grn_reg[4] ),
        .\iv[15]_i_96_8 (\iv[15]_i_96_0 ),
        .\iv[1]_i_8 (bank02_n_197),
        .\iv[2]_i_8 (bank02_n_198),
        .\iv[3]_i_41_0 (sreg_n_64),
        .\iv[3]_i_8 (\sr_reg[8]_56 ),
        .\iv[4]_i_27_0 (bank02_n_259),
        .\iv[4]_i_3 (\iv[4]_i_3 ),
        .\iv[4]_i_35_0 (\iv[4]_i_35 ),
        .\iv[5]_i_15 (bank02_n_279),
        .\iv[5]_i_3 (\iv[5]_i_3 ),
        .\iv[5]_i_7 (\iv[7]_i_7_0 ),
        .\iv[6]_i_10 (\sr_reg[8]_66 ),
        .\iv[6]_i_3 (bank02_n_234),
        .\iv[6]_i_8 (\iv[14]_i_49 ),
        .\iv[7]_i_8 (bank02_n_196),
        .\iv[8]_i_27 (bank02_n_261),
        .\iv[8]_i_34 (\iv[8]_i_34 ),
        .\iv[8]_i_38 (sreg_n_144),
        .\iv[8]_i_4 (\iv[0]_i_25 ),
        .\iv[9]_i_28 (\iv[0]_i_19 ),
        .\iv[9]_i_28_0 (bank02_n_283),
        .\iv[9]_i_4 (bank02_n_206),
        .\iv[9]_i_46_0 (sreg_n_68),
        .mul_a(mul_a[15:0]),
        .mul_a_i(mul_a_i),
        .\mul_a_reg[16] (abus_0[16]),
        .\mul_a_reg[17] (abus_0[17]),
        .\mul_a_reg[18] (abus_0[18]),
        .\mul_a_reg[19] (abus_0[19]),
        .\mul_a_reg[20] (abus_0[20]),
        .\mul_a_reg[21] (abus_0[21]),
        .\mul_a_reg[22] (abus_0[22]),
        .\mul_a_reg[23] (abus_0[23]),
        .\mul_a_reg[24] (abus_0[24]),
        .\mul_a_reg[25] (abus_0[25]),
        .\mul_a_reg[26] (abus_0[26]),
        .\mul_a_reg[27] (abus_0[27]),
        .\mul_a_reg[28] (abus_0[28]),
        .\mul_a_reg[29] (abus_0[29]),
        .\mul_a_reg[30] (abus_0[30]),
        .\mul_a_reg[32] (abus_0[31]),
        .\mul_a_reg[32]_0 (\mul_a_reg[32] ),
        .mul_rslt(mul_rslt),
        .mul_rslt0(mul_rslt0),
        .niho_dsp_a(niho_dsp_a[15:0]),
        .\niho_dsp_a[11] (abus_0[11:8]),
        .\niho_dsp_a[3] (abus_0[3:0]),
        .\niho_dsp_a[7] (abus_0[7:4]),
        .niho_dsp_a_15_sp_1(bank02_n_304),
        .niho_dsp_b(niho_dsp_b),
        .\niho_dsp_b[0]_0 (niho_dsp_b_0_sn_1),
        .\niho_dsp_b[5] (\tr_reg[5] [1]),
        .\niho_dsp_b[5]_0 (\niho_dsp_b[5] ),
        .\niho_dsp_b[5]_1 (\niho_dsp_b[5]_0 ),
        .niho_dsp_b_0_sp_1(\tr_reg[5] [0]),
        .out({p_0_in_2[15:14],out[12:9],p_0_in_2[9],out[8:0]}),
        .p_2_in(p_2_in[6]),
        .\pc_reg[3]_i_2 (rgf_pc[1]),
        .\quo_reg[19] (sreg_n_218),
        .\quo_reg[23] (sreg_n_220),
        .\quo_reg[27] (sreg_n_221),
        .\rem_reg[21] (sreg_n_219),
        .\rem_reg[28] (sreg_n_222),
        .\rem_reg[29] (sreg_n_223),
        .\remden_reg[16] (\remden_reg[16] ),
        .\remden_reg[17] (\remden_reg[17] ),
        .\remden_reg[18] (\remden_reg[18] ),
        .\remden_reg[19] (\remden_reg[19] ),
        .\remden_reg[20] (\remden_reg[20] ),
        .\remden_reg[21] (\remden_reg[21] ),
        .\remden_reg[22] (\remden_reg[22] ),
        .\remden_reg[23] (\remden_reg[23] ),
        .\remden_reg[24] (\remden_reg[24] ),
        .\remden_reg[25] (\remden_reg[25] ),
        .\remden_reg[26] (\remden_reg[26] ),
        .\remden_reg[26]_0 (\remden_reg[26]_0 ),
        .\remden_reg[27] (\remden_reg[27] ),
        .\remden_reg[28] (\remden_reg[28] ),
        .\remden_reg[29] (\remden_reg[29] ),
        .\remden_reg[30] (\remden_reg[30] ),
        .rst_n(rst_n),
        .\sr[4]_i_103 (\iv[3]_i_10_1 ),
        .\sr[4]_i_139_0 (\sr[4]_i_139 ),
        .\sr[4]_i_17 (bank02_n_200),
        .\sr[4]_i_19 (\tr_reg[1]_0 ),
        .\sr[4]_i_19_0 (bank02_n_144),
        .\sr[4]_i_19_1 (\sr[4]_i_16 ),
        .\sr[4]_i_3 (bank02_n_347),
        .\sr[4]_i_31 (\iv[4]_i_9 ),
        .\sr[4]_i_31_0 (bank02_n_181),
        .\sr[4]_i_32 (bank02_n_204),
        .\sr[4]_i_33 (\iv[5]_i_9 ),
        .\sr[4]_i_33_0 (bank02_n_182),
        .\sr[4]_i_34 (bank02_n_203),
        .\sr[4]_i_35 (\iv[10]_i_5 ),
        .\sr[4]_i_35_0 (bank02_n_189),
        .\sr[4]_i_37 (\sr[4]_i_37 ),
        .\sr[4]_i_37_0 (\iv[9]_i_5 ),
        .\sr[4]_i_37_1 (bank02_n_186),
        .\sr[4]_i_38 (\tr[22]_i_3 ),
        .\sr[4]_i_38_0 (\iv[13]_i_17_0 ),
        .\sr[4]_i_39 (\sr[4]_i_39_0 ),
        .\sr[4]_i_39_0 (\iv[8]_i_5 ),
        .\sr[4]_i_39_1 (bank02_n_190),
        .\sr[4]_i_3_0 (\sr[4]_i_3 ),
        .\sr[4]_i_40 (\sr[4]_i_40_0 ),
        .\sr[4]_i_40_0 (\iv[14]_i_5 ),
        .\sr[4]_i_40_1 (bank02_n_178),
        .\sr[4]_i_41 (\iv[1]_i_9 ),
        .\sr[4]_i_41_0 (bank02_n_187),
        .\sr[4]_i_42_0 (\tr[24]_i_3 ),
        .\sr[4]_i_42_1 (\sr[4]_i_42 ),
        .\sr[4]_i_42_2 (bank02_n_251),
        .\sr[4]_i_42_3 (bank02_n_218),
        .\sr[4]_i_42_4 (\iv[7]_i_9 ),
        .\sr[4]_i_42_5 (bank02_n_177),
        .\sr[4]_i_42_6 (\tr[16]_i_6 ),
        .\sr[4]_i_43 (\sr[4]_i_43 ),
        .\sr[4]_i_46 (\iv[3]_i_9 ),
        .\sr[4]_i_46_0 (bank02_n_183),
        .\sr[4]_i_47 (\iv[2]_i_9 ),
        .\sr[4]_i_47_0 (bank02_n_191),
        .\sr[4]_i_66 (bank02_n_247),
        .\sr[4]_i_69_0 (bank02_n_286),
        .\sr[4]_i_73 (\iv[6]_i_10_1 ),
        .\sr[4]_i_74 (\sr_reg[8]_62 ),
        .\sr[4]_i_86 (\iv[1]_i_10_1 ),
        .\sr[4]_i_87_0 (\sr[4]_i_87 ),
        .\sr[4]_i_90_0 (\sr_reg[8]_67 ),
        .\sr[4]_i_91 (\sr_reg[8]_5 ),
        .\sr[4]_i_91_0 (bank02_n_243),
        .\sr[4]_i_94_0 (bank02_n_291),
        .\sr[5]_i_2_0 (\sr[5]_i_2 ),
        .\sr[5]_i_3 (bank02_n_388),
        .\sr[5]_i_3_0 (\sr[4]_i_36 ),
        .\sr[5]_i_3_1 (bank02_n_217),
        .\sr[5]_i_3_2 (bank02_n_385),
        .\sr[5]_i_3_3 (bank02_n_390),
        .\sr[5]_i_3_4 (\sr[5]_i_3 ),
        .\sr[5]_i_3_5 (\tr[30]_i_3 ),
        .\sr[6]_i_10 (bank02_n_298),
        .\sr[6]_i_11_0 (\sr[4]_i_89 ),
        .\sr[6]_i_11_1 (\sr_reg[8]_12 ),
        .\sr[6]_i_13 (\sr[6]_i_13 ),
        .\sr[6]_i_38_0 (\sr[6]_i_12 ),
        .\sr[6]_i_4_0 (bank02_n_216),
        .\sr[6]_i_4_1 (bank02_n_235),
        .\sr[6]_i_4_2 (\sr[6]_i_4 ),
        .\sr[6]_i_4_3 (\iv[0]_i_10_1 ),
        .\sr_reg[0]_0 (sreg_n_280),
        .\sr_reg[0]_1 (sreg_n_285),
        .\sr_reg[0]_10 (sreg_n_294),
        .\sr_reg[0]_11 (sreg_n_295),
        .\sr_reg[0]_12 (sreg_n_296),
        .\sr_reg[0]_13 (sreg_n_297),
        .\sr_reg[0]_14 (sreg_n_298),
        .\sr_reg[0]_15 (sreg_n_299),
        .\sr_reg[0]_16 (sreg_n_300),
        .\sr_reg[0]_17 (sreg_n_301),
        .\sr_reg[0]_18 (sreg_n_302),
        .\sr_reg[0]_19 (sreg_n_303),
        .\sr_reg[0]_2 (sreg_n_286),
        .\sr_reg[0]_20 (sreg_n_304),
        .\sr_reg[0]_21 (sreg_n_305),
        .\sr_reg[0]_22 (sreg_n_306),
        .\sr_reg[0]_23 (sreg_n_307),
        .\sr_reg[0]_24 (sreg_n_308),
        .\sr_reg[0]_25 (sreg_n_309),
        .\sr_reg[0]_26 (sreg_n_310),
        .\sr_reg[0]_27 (sreg_n_311),
        .\sr_reg[0]_28 (sreg_n_312),
        .\sr_reg[0]_29 (sreg_n_313),
        .\sr_reg[0]_3 (sreg_n_287),
        .\sr_reg[0]_30 (sreg_n_314),
        .\sr_reg[0]_31 (sreg_n_315),
        .\sr_reg[0]_32 (sreg_n_316),
        .\sr_reg[0]_33 (sreg_n_317),
        .\sr_reg[0]_34 (sreg_n_318),
        .\sr_reg[0]_35 (sreg_n_319),
        .\sr_reg[0]_36 (sreg_n_320),
        .\sr_reg[0]_37 (sreg_n_321),
        .\sr_reg[0]_38 (sreg_n_322),
        .\sr_reg[0]_39 (sreg_n_323),
        .\sr_reg[0]_4 (sreg_n_288),
        .\sr_reg[0]_40 (sreg_n_324),
        .\sr_reg[0]_41 (sreg_n_325),
        .\sr_reg[0]_42 (sreg_n_326),
        .\sr_reg[0]_43 (sreg_n_327),
        .\sr_reg[0]_44 (sreg_n_328),
        .\sr_reg[0]_45 (sreg_n_329),
        .\sr_reg[0]_46 (sreg_n_330),
        .\sr_reg[0]_47 (sreg_n_331),
        .\sr_reg[0]_48 (sreg_n_332),
        .\sr_reg[0]_49 (sreg_n_333),
        .\sr_reg[0]_5 (sreg_n_289),
        .\sr_reg[0]_50 (sreg_n_334),
        .\sr_reg[0]_51 (sreg_n_335),
        .\sr_reg[0]_52 (sreg_n_336),
        .\sr_reg[0]_53 (sreg_n_337),
        .\sr_reg[0]_54 (sreg_n_338),
        .\sr_reg[0]_55 (sreg_n_339),
        .\sr_reg[0]_56 (sreg_n_340),
        .\sr_reg[0]_57 (sreg_n_341),
        .\sr_reg[0]_58 (sreg_n_342),
        .\sr_reg[0]_59 (sreg_n_343),
        .\sr_reg[0]_6 (sreg_n_290),
        .\sr_reg[0]_60 (sreg_n_344),
        .\sr_reg[0]_61 (sreg_n_345),
        .\sr_reg[0]_62 (sreg_n_346),
        .\sr_reg[0]_63 (sreg_n_347),
        .\sr_reg[0]_64 (sreg_n_348),
        .\sr_reg[0]_65 (sreg_n_349),
        .\sr_reg[0]_66 (sreg_n_350),
        .\sr_reg[0]_67 (sreg_n_351),
        .\sr_reg[0]_68 (sreg_n_352),
        .\sr_reg[0]_69 (sreg_n_353),
        .\sr_reg[0]_7 (sreg_n_291),
        .\sr_reg[0]_70 (sreg_n_354),
        .\sr_reg[0]_71 (sreg_n_355),
        .\sr_reg[0]_72 (sreg_n_356),
        .\sr_reg[0]_73 (sreg_n_357),
        .\sr_reg[0]_74 (sreg_n_358),
        .\sr_reg[0]_75 (sreg_n_359),
        .\sr_reg[0]_76 (sreg_n_360),
        .\sr_reg[0]_77 (sreg_n_361),
        .\sr_reg[0]_78 (sreg_n_362),
        .\sr_reg[0]_79 (sreg_n_363),
        .\sr_reg[0]_8 (sreg_n_292),
        .\sr_reg[0]_80 (sreg_n_364),
        .\sr_reg[0]_81 (sreg_n_365),
        .\sr_reg[0]_82 (sreg_n_366),
        .\sr_reg[0]_83 (sreg_n_367),
        .\sr_reg[0]_84 (sreg_n_368),
        .\sr_reg[0]_85 (sreg_n_369),
        .\sr_reg[0]_86 (sreg_n_370),
        .\sr_reg[0]_87 (sreg_n_371),
        .\sr_reg[0]_88 (sreg_n_372),
        .\sr_reg[0]_89 (sreg_n_373),
        .\sr_reg[0]_9 (sreg_n_293),
        .\sr_reg[0]_90 (sreg_n_374),
        .\sr_reg[0]_91 (sreg_n_375),
        .\sr_reg[0]_92 (sreg_n_376),
        .\sr_reg[0]_93 (sreg_n_377),
        .\sr_reg[0]_94 (sreg_n_378),
        .\sr_reg[0]_95 (sreg_n_379),
        .\sr_reg[0]_96 (sreg_n_380),
        .\sr_reg[0]_97 (\sr_reg[0] ),
        .\sr_reg[10]_0 (\sr_reg[10]_0 ),
        .\sr_reg[11]_0 (\sr_reg[11]_0 ),
        .\sr_reg[15]_0 (\sr_reg[15]_0 ),
        .\sr_reg[1]_0 (sreg_n_16),
        .\sr_reg[1]_1 (sreg_n_17),
        .\sr_reg[1]_2 (sreg_n_18),
        .\sr_reg[1]_3 (sreg_n_19),
        .\sr_reg[1]_4 (sreg_n_275),
        .\sr_reg[1]_5 (sreg_n_276),
        .\sr_reg[1]_6 (sreg_n_282),
        .\sr_reg[1]_7 (sreg_n_283),
        .\sr_reg[1]_8 (sreg_n_284),
        .\sr_reg[1]_9 (\sr_reg[1]_0 ),
        .\sr_reg[2]_0 (\sr_reg[2]_0 ),
        .\sr_reg[3]_0 (\sr_reg[3]_0 ),
        .\sr_reg[4]_0 (\sr_reg[4]_0 ),
        .\sr_reg[4]_1 (\sr_reg[4]_1 ),
        .\sr_reg[4]_2 (\sr_reg[4]_4 ),
        .\sr_reg[5]_0 (\sr_reg[5] ),
        .\sr_reg[5]_1 (\sr_reg[5]_0 ),
        .\sr_reg[5]_2 (\sr_reg[5]_1 ),
        .\sr_reg[5]_3 (\art/add/sr[5]_i_14 [3]),
        .\sr_reg[5]_4 (\sr_reg[5]_2 ),
        .\sr_reg[6]_0 (sreg_n_126),
        .\sr_reg[6]_1 (sreg_n_127),
        .\sr_reg[6]_2 (sreg_n_137),
        .\sr_reg[6]_3 (\sr_reg[6]_5 ),
        .\sr_reg[6]_4 (\sr_reg[6]_10 ),
        .\sr_reg[6]_5 (\sr_reg[6]_11 ),
        .\sr_reg[6]_6 (\sr_reg[6]_12 ),
        .\sr_reg[6]_i_6_0 (\sr_reg[6]_i_6 ),
        .\sr_reg[6]_i_6_1 (\sr_reg[6]_i_6_0 ),
        .\sr_reg[6]_i_6_2 (\sr_reg[6]_i_6_1 ),
        .\sr_reg[7]_0 (\sr_reg[7] ),
        .\sr_reg[7]_1 (\sr_reg[7]_0 ),
        .\sr_reg[7]_2 (\sr_reg[7]_1 ),
        .\sr_reg[7]_3 (\sr_reg[7]_2 ),
        .\sr_reg[7]_4 (\sr_reg[7]_4 ),
        .\sr_reg[8]_0 (\sr_reg[8] ),
        .\sr_reg[8]_1 (\sr_reg[8]_0 ),
        .\sr_reg[8]_10 (sreg_n_32),
        .\sr_reg[8]_100 (sreg_n_143),
        .\sr_reg[8]_101 (sreg_n_146),
        .\sr_reg[8]_102 (sreg_n_147),
        .\sr_reg[8]_103 (sreg_n_148),
        .\sr_reg[8]_104 (sreg_n_149),
        .\sr_reg[8]_105 (sreg_n_150),
        .\sr_reg[8]_106 (sreg_n_152),
        .\sr_reg[8]_107 (sreg_n_153),
        .\sr_reg[8]_108 (\sr_reg[8]_116 ),
        .\sr_reg[8]_109 (sreg_n_156),
        .\sr_reg[8]_11 (sreg_n_33),
        .\sr_reg[8]_110 (sreg_n_157),
        .\sr_reg[8]_111 (\sr_reg[8]_130 ),
        .\sr_reg[8]_112 (\sr_reg[8]_131 ),
        .\sr_reg[8]_113 (\sr_reg[8]_132 ),
        .\sr_reg[8]_114 (\sr_reg[8]_133 ),
        .\sr_reg[8]_115 (\sr_reg[8]_134 ),
        .\sr_reg[8]_116 (\sr_reg[8]_135 ),
        .\sr_reg[8]_117 (\sr_reg[8]_136 ),
        .\sr_reg[8]_118 (\sr_reg[8]_137 ),
        .\sr_reg[8]_119 (\sr_reg[8]_138 ),
        .\sr_reg[8]_12 (\sr_reg[8]_38 ),
        .\sr_reg[8]_120 (\sr_reg[8]_139 ),
        .\sr_reg[8]_121 (\sr_reg[8]_140 ),
        .\sr_reg[8]_122 (\sr_reg[8]_141 ),
        .\sr_reg[8]_123 (\sr_reg[8]_142 ),
        .\sr_reg[8]_124 (\sr_reg[8]_143 ),
        .\sr_reg[8]_125 (\sr_reg[8]_144 ),
        .\sr_reg[8]_126 (\sr_reg[8]_145 ),
        .\sr_reg[8]_127 (\sr_reg[8]_146 ),
        .\sr_reg[8]_128 (\sr_reg[8]_147 ),
        .\sr_reg[8]_129 (\sr_reg[8]_148 ),
        .\sr_reg[8]_13 (sreg_n_36),
        .\sr_reg[8]_130 (\sr_reg[8]_149 ),
        .\sr_reg[8]_131 (\sr_reg[8]_150 ),
        .\sr_reg[8]_132 (\sr_reg[8]_151 ),
        .\sr_reg[8]_133 (sreg_n_262),
        .\sr_reg[8]_134 (sreg_n_263),
        .\sr_reg[8]_135 (sreg_n_264),
        .\sr_reg[8]_136 (sreg_n_265),
        .\sr_reg[8]_137 (sreg_n_266),
        .\sr_reg[8]_138 (sreg_n_267),
        .\sr_reg[8]_139 (sreg_n_268),
        .\sr_reg[8]_14 (\sr_reg[8]_40 ),
        .\sr_reg[8]_140 (sreg_n_269),
        .\sr_reg[8]_141 (sreg_n_270),
        .\sr_reg[8]_142 (\sr_reg[8]_155 ),
        .\sr_reg[8]_143 (\sr_reg[8]_156 ),
        .\sr_reg[8]_144 (\sr_reg[8]_157 ),
        .\sr_reg[8]_145 (sreg_n_274),
        .\sr_reg[8]_146 (sreg_n_381),
        .\sr_reg[8]_147 (sreg_n_382),
        .\sr_reg[8]_148 (sreg_n_383),
        .\sr_reg[8]_149 (sreg_n_384),
        .\sr_reg[8]_15 (\sr_reg[8]_41 ),
        .\sr_reg[8]_150 (sreg_n_385),
        .\sr_reg[8]_151 (sreg_n_386),
        .\sr_reg[8]_152 (sreg_n_387),
        .\sr_reg[8]_153 (sreg_n_388),
        .\sr_reg[8]_154 (sreg_n_389),
        .\sr_reg[8]_155 (sreg_n_390),
        .\sr_reg[8]_156 (sreg_n_391),
        .\sr_reg[8]_157 (sreg_n_392),
        .\sr_reg[8]_158 (sreg_n_393),
        .\sr_reg[8]_159 (sreg_n_394),
        .\sr_reg[8]_16 (\sr_reg[8]_43 ),
        .\sr_reg[8]_160 (sreg_n_395),
        .\sr_reg[8]_161 (sreg_n_396),
        .\sr_reg[8]_162 (sreg_n_397),
        .\sr_reg[8]_163 (sreg_n_398),
        .\sr_reg[8]_164 (sreg_n_399),
        .\sr_reg[8]_165 (sreg_n_400),
        .\sr_reg[8]_166 (sreg_n_401),
        .\sr_reg[8]_167 (sreg_n_402),
        .\sr_reg[8]_168 (sreg_n_403),
        .\sr_reg[8]_169 (sreg_n_404),
        .\sr_reg[8]_17 (sreg_n_43),
        .\sr_reg[8]_170 (sreg_n_405),
        .\sr_reg[8]_171 (sreg_n_406),
        .\sr_reg[8]_172 (sreg_n_407),
        .\sr_reg[8]_173 (sreg_n_408),
        .\sr_reg[8]_174 (sreg_n_409),
        .\sr_reg[8]_175 (sreg_n_410),
        .\sr_reg[8]_176 (sreg_n_411),
        .\sr_reg[8]_177 (sreg_n_412),
        .\sr_reg[8]_178 (sreg_n_413),
        .\sr_reg[8]_179 (sreg_n_414),
        .\sr_reg[8]_18 (\sr_reg[8]_44 ),
        .\sr_reg[8]_180 (sreg_n_415),
        .\sr_reg[8]_181 (sreg_n_416),
        .\sr_reg[8]_182 (sreg_n_417),
        .\sr_reg[8]_183 (sreg_n_418),
        .\sr_reg[8]_184 (sreg_n_419),
        .\sr_reg[8]_185 (sreg_n_420),
        .\sr_reg[8]_186 (sreg_n_421),
        .\sr_reg[8]_187 (sreg_n_422),
        .\sr_reg[8]_188 (sreg_n_423),
        .\sr_reg[8]_189 (sreg_n_424),
        .\sr_reg[8]_19 (sreg_n_45),
        .\sr_reg[8]_190 (sreg_n_425),
        .\sr_reg[8]_191 (sreg_n_426),
        .\sr_reg[8]_192 (sreg_n_427),
        .\sr_reg[8]_193 (sreg_n_428),
        .\sr_reg[8]_194 (sreg_n_429),
        .\sr_reg[8]_195 (sreg_n_430),
        .\sr_reg[8]_196 (sreg_n_431),
        .\sr_reg[8]_197 (sreg_n_432),
        .\sr_reg[8]_198 (sreg_n_433),
        .\sr_reg[8]_199 (sreg_n_434),
        .\sr_reg[8]_2 (sreg_n_24),
        .\sr_reg[8]_20 (\sr_reg[8]_45 ),
        .\sr_reg[8]_200 (sreg_n_435),
        .\sr_reg[8]_201 (sreg_n_436),
        .\sr_reg[8]_202 (sreg_n_437),
        .\sr_reg[8]_203 (sreg_n_438),
        .\sr_reg[8]_204 (sreg_n_439),
        .\sr_reg[8]_205 (sreg_n_440),
        .\sr_reg[8]_206 (sreg_n_441),
        .\sr_reg[8]_207 (sreg_n_442),
        .\sr_reg[8]_208 (sreg_n_443),
        .\sr_reg[8]_209 (sreg_n_444),
        .\sr_reg[8]_21 (sreg_n_47),
        .\sr_reg[8]_210 (sreg_n_445),
        .\sr_reg[8]_211 (sreg_n_446),
        .\sr_reg[8]_212 (sreg_n_447),
        .\sr_reg[8]_213 (sreg_n_448),
        .\sr_reg[8]_214 (sreg_n_449),
        .\sr_reg[8]_215 (\sr_reg[8]_9 ),
        .\sr_reg[8]_216 (sreg_n_451),
        .\sr_reg[8]_217 (sreg_n_452),
        .\sr_reg[8]_218 (\sr_reg[8]_158 ),
        .\sr_reg[8]_219 (\sr_reg[8]_159 ),
        .\sr_reg[8]_22 (\sr_reg[8]_46 ),
        .\sr_reg[8]_220 (\sr_reg[8]_160 ),
        .\sr_reg[8]_221 (\sr_reg[8]_161 ),
        .\sr_reg[8]_222 (\sr_reg[8]_162 ),
        .\sr_reg[8]_223 (\sr_reg[8]_163 ),
        .\sr_reg[8]_224 (sreg_n_466),
        .\sr_reg[8]_225 (sreg_n_467),
        .\sr_reg[8]_226 (sreg_n_468),
        .\sr_reg[8]_227 (sreg_n_469),
        .\sr_reg[8]_228 (\sr_reg[8]_169 ),
        .\sr_reg[8]_23 (\sr_reg[8]_47 ),
        .\sr_reg[8]_24 (\sr_reg[8]_48 ),
        .\sr_reg[8]_25 (\sr_reg[8]_49 ),
        .\sr_reg[8]_26 (\sr_reg[8]_50 ),
        .\sr_reg[8]_27 (sreg_n_54),
        .\sr_reg[8]_28 (sreg_n_55),
        .\sr_reg[8]_29 (\sr_reg[8]_51 ),
        .\sr_reg[8]_3 (\sr_reg[8]_32 ),
        .\sr_reg[8]_30 (sreg_n_57),
        .\sr_reg[8]_31 (\sr_reg[8]_52 ),
        .\sr_reg[8]_32 (\sr_reg[8]_53 ),
        .\sr_reg[8]_33 (\sr_reg[8]_54 ),
        .\sr_reg[8]_34 (sreg_n_62),
        .\sr_reg[8]_35 (\sr_reg[8]_55 ),
        .\sr_reg[8]_36 (sreg_n_65),
        .\sr_reg[8]_37 (sreg_n_67),
        .\sr_reg[8]_38 (sreg_n_69),
        .\sr_reg[8]_39 (sreg_n_70),
        .\sr_reg[8]_4 (sreg_n_26),
        .\sr_reg[8]_40 (\sr_reg[8]_57 ),
        .\sr_reg[8]_41 (\sr_reg[8]_58 ),
        .\sr_reg[8]_42 (sreg_n_73),
        .\sr_reg[8]_43 (sreg_n_74),
        .\sr_reg[8]_44 (sreg_n_75),
        .\sr_reg[8]_45 (sreg_n_76),
        .\sr_reg[8]_46 (sreg_n_77),
        .\sr_reg[8]_47 (\sr_reg[8]_65 ),
        .\sr_reg[8]_48 (sreg_n_79),
        .\sr_reg[8]_49 (sreg_n_80),
        .\sr_reg[8]_5 (\sr_reg[8]_33 ),
        .\sr_reg[8]_50 (\sr_reg[8]_78 ),
        .\sr_reg[8]_51 (\sr_reg[8]_79 ),
        .\sr_reg[8]_52 (sreg_n_84),
        .\sr_reg[8]_53 (sreg_n_85),
        .\sr_reg[8]_54 (sreg_n_86),
        .\sr_reg[8]_55 (\sr_reg[8]_8 ),
        .\sr_reg[8]_56 (\sr_reg[8]_81 ),
        .\sr_reg[8]_57 (\sr_reg[8]_82 ),
        .\sr_reg[8]_58 (\sr_reg[8]_19 ),
        .\sr_reg[8]_59 (\sr_reg[8]_83 ),
        .\sr_reg[8]_6 (sreg_n_28),
        .\sr_reg[8]_60 (\sr_reg[8]_84 ),
        .\sr_reg[8]_61 (\sr_reg[8]_25 ),
        .\sr_reg[8]_62 (sreg_n_94),
        .\sr_reg[8]_63 (sreg_n_95),
        .\sr_reg[8]_64 (\sr_reg[8]_30 ),
        .\sr_reg[8]_65 (\sr_reg[8]_87 ),
        .\sr_reg[8]_66 (\sr_reg[8]_88 ),
        .\sr_reg[8]_67 (sreg_n_99),
        .\sr_reg[8]_68 (\sr_reg[8]_89 ),
        .\sr_reg[8]_69 (sreg_n_101),
        .\sr_reg[8]_7 (sreg_n_29),
        .\sr_reg[8]_70 (sreg_n_102),
        .\sr_reg[8]_71 (sreg_n_103),
        .\sr_reg[8]_72 (\sr_reg[8]_90 ),
        .\sr_reg[8]_73 (\sr_reg[8]_91 ),
        .\sr_reg[8]_74 (\sr_reg[8]_92 ),
        .\sr_reg[8]_75 (sreg_n_107),
        .\sr_reg[8]_76 (\sr_reg[8]_109 ),
        .\sr_reg[8]_77 (\sr_reg[8]_113 ),
        .\sr_reg[8]_78 (sreg_n_113),
        .\sr_reg[8]_79 (\sr_reg[8]_36 ),
        .\sr_reg[8]_8 (sreg_n_30),
        .\sr_reg[8]_80 (\sr_reg[8]_114 ),
        .\sr_reg[8]_81 (sreg_n_118),
        .\sr_reg[8]_82 (sreg_n_119),
        .\sr_reg[8]_83 (sreg_n_120),
        .\sr_reg[8]_84 (\sr_reg[8]_119 ),
        .\sr_reg[8]_85 (sreg_n_122),
        .\sr_reg[8]_86 (sreg_n_123),
        .\sr_reg[8]_87 (sreg_n_124),
        .\sr_reg[8]_88 (sreg_n_125),
        .\sr_reg[8]_89 (sreg_n_129),
        .\sr_reg[8]_9 (sreg_n_31),
        .\sr_reg[8]_90 (sreg_n_130),
        .\sr_reg[8]_91 (sreg_n_131),
        .\sr_reg[8]_92 (sreg_n_132),
        .\sr_reg[8]_93 (sreg_n_133),
        .\sr_reg[8]_94 (sreg_n_134),
        .\sr_reg[8]_95 (sreg_n_135),
        .\sr_reg[8]_96 (sreg_n_138),
        .\sr_reg[8]_97 (\sr_reg[8]_125 ),
        .\sr_reg[8]_98 (\sr_reg[8]_108 ),
        .\sr_reg[8]_99 (sreg_n_142),
        .\stat[0]_i_6 (\stat[0]_i_6 ),
        .\stat_reg[0] (\stat_reg[0] ),
        .\stat_reg[1] (\stat_reg[1] ),
        .\tr[16]_i_2 (bank02_n_140),
        .\tr[16]_i_2_0 (\sr_reg[8]_37 ),
        .\tr[18]_i_9 (bank02_n_274),
        .\tr[19]_i_2 (\tr[19]_i_2_0 ),
        .\tr[19]_i_2_0 (\tr[19]_i_2_1 ),
        .\tr[19]_i_6 (bank02_n_300),
        .\tr[19]_i_7 (bank02_n_207),
        .\tr[20]_i_8 (bank02_n_289),
        .\tr[20]_i_9 (\sr_reg[8]_129 ),
        .\tr[21]_i_8 (bank02_n_266),
        .\tr[21]_i_9 (\sr_reg[8]_97 ),
        .\tr[21]_i_9_0 (bank02_n_267),
        .\tr[21]_i_9_1 (\sr_reg[8]_110 ),
        .\tr[22]_i_9 (\sr_reg[6]_1 ),
        .\tr[23]_i_3 (\sr_reg[8]_3 ),
        .\tr[23]_i_5 (\tr[22]_i_11 ),
        .\tr[23]_i_6 (\sr_reg[8]_124 ),
        .\tr[23]_i_6_0 (\sr[4]_i_61 ),
        .\tr[23]_i_7 (\sr_reg[8]_77 ),
        .\tr[24]_i_9 (\sr_reg[8]_126 ),
        .\tr[25]_i_9 (\sr_reg[8]_61 ),
        .\tr[26]_i_6 (\sr_reg[8]_73 ),
        .\tr[26]_i_7 (\sr_reg[8]_111 ),
        .\tr[26]_i_7_0 (bank02_n_280),
        .\tr[27]_i_7 (bank02_n_301),
        .\tr[27]_i_9 (\tr[24]_i_3_0 ),
        .\tr[28]_i_3 (\tr[19]_i_3_0 ),
        .\tr[28]_i_8_0 (bank02_n_260),
        .\tr[28]_i_9 (bank02_n_295),
        .\tr[29]_i_2 (\tr[29]_i_2 ),
        .\tr[30]_i_10 (bank02_n_282),
        .\tr_reg[23]_i_11_0 (\tr_reg[23]_i_11 ),
        .\tr_reg[23]_i_11_1 (\tr_reg[23]_i_11_0 ),
        .\tr_reg[23]_i_11_2 (\tr_reg[23]_i_11_1 ),
        .\tr_reg[23]_i_11_3 (\tr_reg[23]_i_11_2 ),
        .\tr_reg[31] (\tr_reg[31]_1 ),
        .\tr_reg[31]_0 (\tr_reg[31]_2 ),
        .\tr_reg[31]_i_13_0 (\tr_reg[31]_i_13 ),
        .\tr_reg[31]_i_13_1 (\tr_reg[31]_i_13_0 ),
        .\tr_reg[31]_i_13_2 (\tr_reg[31]_i_13_1 ),
        .\tr_reg[31]_i_32_0 (\tr_reg[31]_i_32 ),
        .\tr_reg[31]_i_32_1 (\tr_reg[31]_i_32_0 ),
        .\tr_reg[31]_i_32_2 (\tr_reg[31]_i_32_1 ),
        .\tr_reg[31]_i_32_3 (\tr_reg[31]_i_32_2 ));
  niho_rgf_treg treg
       (.SR(p_0_in),
        .cbus(cbus),
        .clk(clk),
        .\tr_reg[0]_0 (\tr_reg[0] [1]),
        .\tr_reg[31]_0 (\tr_reg[31] ));
endmodule

module niho_rgf_bank
   (.out({gr20[15],gr20[14],gr20[13],gr20[12],gr20[11],gr20[10],gr20[9],gr20[8],gr20[7],gr20[6],gr20[5],gr20[4],gr20[3],gr20[2],gr20[1],gr20[0]}),
    .\grn_reg[15] ({gr21[15],gr21[14],gr21[13],gr21[12],gr21[11],gr21[10],gr21[9],gr21[8],gr21[7],gr21[6],gr21[5],gr21[4],gr21[3],gr21[2],gr21[1],gr21[0]}),
    .\grn_reg[15]_0 ({gr22[15],gr22[14],gr22[13],gr22[12],gr22[11],gr22[10],gr22[9],gr22[8],gr22[7],gr22[6],gr22[5],gr22[4],gr22[3],gr22[2],gr22[1],gr22[0]}),
    .\grn_reg[15]_1 ({gr23[15],gr23[14],gr23[13],gr23[12],gr23[11],gr23[10],gr23[9],gr23[8],gr23[7],gr23[6],gr23[5],gr23[4],gr23[3],gr23[2],gr23[1],gr23[0]}),
    .\grn_reg[15]_2 ({gr24[15],gr24[14],gr24[13],gr24[12],gr24[11],gr24[10],gr24[9],gr24[8],gr24[7],gr24[6],gr24[5],gr24[4],gr24[3],gr24[2],gr24[1],gr24[0]}),
    .\grn_reg[15]_3 ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_4 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    .\grn_reg[15]_5 ({gr27[15],gr27[14],gr27[13],gr27[12],gr27[11],gr27[10],gr27[9],gr27[8],gr27[7],gr27[6],gr27[5],gr27[4],gr27[3],gr27[2],gr27[1],gr27[0]}),
    p_2_in,
    \badr[21]_INST_0_i_1 ,
    \tr_reg[5] ,
    \bdatw[8]_INST_0_i_2 ,
    \tr_reg[0] ,
    \iv[7]_i_33 ,
    \sr_reg[8] ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr[4]_i_21_0 ,
    \sr_reg[8]_2 ,
    \iv[7]_i_37_0 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr[4]_i_147_0 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr[4]_i_65_0 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \iv[13]_i_27 ,
    \sr_reg[8]_21 ,
    \iv[8]_i_20 ,
    \sr_reg[8]_22 ,
    \iv[14]_i_35_0 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr[4]_i_116_0 ,
    \sr_reg[8]_25 ,
    \tr[17]_i_9_0 ,
    \tr[24]_i_10_0 ,
    \tr[30]_i_10_0 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \tr[20]_i_9_0 ,
    \tr[22]_i_9_0 ,
    \iv[12]_i_27_0 ,
    \iv[13]_i_29_0 ,
    \sr_reg[8]_28 ,
    \tr[18]_i_9_0 ,
    \tr[26]_i_9_0 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \iv[8]_i_30 ,
    \sr_reg[8]_33 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \sr_reg[8]_36 ,
    \iv[7]_i_17 ,
    \iv[15]_i_94 ,
    \sr_reg[8]_37 ,
    \sr_reg[8]_38 ,
    \iv[10]_i_10 ,
    \sr_reg[8]_39 ,
    \sr_reg[8]_40 ,
    \sr_reg[8]_41 ,
    \iv[5]_i_23 ,
    \sr_reg[8]_42 ,
    \iv[9]_i_11 ,
    \sr_reg[8]_43 ,
    \sr_reg[8]_44 ,
    \sr_reg[8]_45 ,
    \sr_reg[8]_46 ,
    \sr_reg[8]_47 ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    \sr_reg[8]_50 ,
    \sr_reg[8]_51 ,
    \sr_reg[8]_52 ,
    \tr[16]_i_9_0 ,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    \sr_reg[8]_57 ,
    \sr_reg[8]_58 ,
    \sr_reg[8]_59 ,
    \sr_reg[8]_60 ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    \sr_reg[8]_63 ,
    \sr_reg[8]_64 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    \sr_reg[8]_67 ,
    \sr_reg[8]_68 ,
    \sr_reg[8]_69 ,
    \sr_reg[8]_70 ,
    \sr_reg[8]_71 ,
    \sr_reg[8]_72 ,
    \sr_reg[8]_73 ,
    \sr_reg[8]_74 ,
    \sr_reg[8]_75 ,
    \sr_reg[8]_76 ,
    \sr_reg[8]_77 ,
    \sr_reg[8]_78 ,
    \sr_reg[8]_79 ,
    \sr_reg[8]_80 ,
    \sr_reg[8]_81 ,
    \sr_reg[8]_82 ,
    \sr_reg[8]_83 ,
    \sr_reg[8]_84 ,
    \sr_reg[8]_85 ,
    \iv[7]_i_25 ,
    \sr_reg[8]_86 ,
    \sr_reg[8]_87 ,
    \sr_reg[8]_88 ,
    \sr_reg[8]_89 ,
    \sr_reg[8]_90 ,
    \sr_reg[8]_91 ,
    \sr_reg[6] ,
    \sr_reg[8]_92 ,
    \badr[14]_INST_0_i_1 ,
    \sr_reg[8]_93 ,
    \sr_reg[6]_0 ,
    \badr[0]_INST_0_i_1 ,
    \iv[0]_i_25 ,
    \badr[15]_INST_0_i_1 ,
    \sr_reg[8]_94 ,
    \sr_reg[8]_95 ,
    \sr_reg[6]_1 ,
    \sr_reg[8]_96 ,
    \sr_reg[8]_97 ,
    \sr_reg[6]_2 ,
    \sr_reg[8]_98 ,
    \sr_reg[6]_3 ,
    \sr_reg[6]_4 ,
    \sr_reg[8]_99 ,
    \sr_reg[8]_100 ,
    \iv[14]_i_49 ,
    \sr_reg[8]_101 ,
    \sr_reg[8]_102 ,
    \badr[14]_INST_0_i_1_0 ,
    \sr_reg[8]_103 ,
    \sr_reg[8]_104 ,
    \sr_reg[8]_105 ,
    \badr[0]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1 ,
    \sr_reg[8]_106 ,
    \sr_reg[8]_107 ,
    \sr_reg[8]_108 ,
    \sr_reg[8]_109 ,
    \sr_reg[8]_110 ,
    \sr_reg[6]_5 ,
    \sr_reg[8]_111 ,
    \sr_reg[8]_112 ,
    \sr_reg[8]_113 ,
    \sr_reg[6]_6 ,
    \sr_reg[8]_114 ,
    \sr_reg[8]_115 ,
    \sr_reg[8]_116 ,
    \sr_reg[8]_117 ,
    \sr_reg[8]_118 ,
    \sr_reg[6]_7 ,
    \sr_reg[8]_119 ,
    \badr[5]_INST_0_i_1 ,
    \niho_dsp_a[15]_INST_0_i_3 ,
    \sr_reg[8]_120 ,
    p_0_in,
    p_1_in,
    \iv[15]_i_108 ,
    \iv[15]_i_108_0 ,
    \iv[15]_i_108_1 ,
    \iv[15]_i_108_2 ,
    \iv[15]_i_108_3 ,
    \iv[15]_i_108_4 ,
    \iv[15]_i_108_5 ,
    \iv[15]_i_108_6 ,
    \iv[15]_i_108_7 ,
    \iv[15]_i_108_8 ,
    \sr[4]_i_51_0 ,
    \art/add/iv[7]_i_32 ,
    \art/add/sr[5]_i_14 ,
    \sr_reg[6]_8 ,
    \art/add/sr[5]_i_18 ,
    CO,
    abus_o,
    bbus_o,
    \sr_reg[8]_121 ,
    \sr_reg[8]_122 ,
    \sr_reg[8]_123 ,
    \sr_reg[8]_124 ,
    \sr_reg[8]_125 ,
    \sr_reg[8]_126 ,
    \sr_reg[6]_9 ,
    \sr_reg[8]_127 ,
    \sr_reg[6]_10 ,
    \sr_reg[6]_11 ,
    niho_dsp_a,
    \sr_reg[8]_128 ,
    \sr_reg[8]_129 ,
    \sr_reg[8]_130 ,
    \sr_reg[8]_131 ,
    \sr_reg[8]_132 ,
    \grn_reg[15]_6 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_7 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[15]_8 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_9 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    \tr_reg[27] ,
    niho_dsp_c,
    \tr_reg[23] ,
    \tr_reg[23]_0 ,
    \tr_reg[29] ,
    \tr_reg[29]_0 ,
    \tr_reg[28] ,
    \tr_reg[28]_0 ,
    \tr_reg[21] ,
    \tr_reg[21]_0 ,
    \tr_reg[19] ,
    \tr_reg[19]_0 ,
    \tr_reg[27]_0 ,
    \tr_reg[27]_1 ,
    DI,
    bbus_0,
    \iv[13]_i_17 ,
    \iv[13]_i_17_0 ,
    \iv[13]_i_17_1 ,
    \tr[17]_i_3_0 ,
    \abus_o[11] ,
    \sr[4]_i_36 ,
    \abus_o[7] ,
    \iv[7]_i_7 ,
    \iv[7]_i_7_0 ,
    \iv[7]_i_7_1 ,
    \tr_reg[1] ,
    \tr_reg[16] ,
    \tr_reg[1]_0 ,
    \niho_dsp_a[16] ,
    \tr[16]_i_6_0 ,
    \tr[16]_i_6_1 ,
    \sr_reg[4] ,
    \sr_reg[4]_0 ,
    \sr[4]_i_5_0 ,
    \sr[4]_i_5_1 ,
    \sr[4]_i_5_2 ,
    \sr[4]_i_42 ,
    \tr[23]_i_7_0 ,
    \sr[4]_i_89_0 ,
    \sr[4]_i_43 ,
    \sr[4]_i_43_0 ,
    \tr[17]_i_3_1 ,
    \sr[4]_i_5_3 ,
    \sr[4]_i_21_1 ,
    \tr[18]_i_3_0 ,
    \sr[4]_i_21_2 ,
    \sr[4]_i_21_3 ,
    \sr[4]_i_21_4 ,
    \tr[19]_i_3_0 ,
    \tr[19]_i_3_1 ,
    \sr[4]_i_5_4 ,
    \sr[4]_i_5_5 ,
    \sr[4]_i_20_0 ,
    \sr[4]_i_20_1 ,
    \iv[13]_i_2 ,
    \tr[30]_i_3_0 ,
    \sr[4]_i_20_2 ,
    \sr[4]_i_20_3 ,
    \iv[12]_i_2 ,
    \tr[29]_i_3_0 ,
    \sr[4]_i_44_0 ,
    \iv[0]_i_3 ,
    \iv[0]_i_3_0 ,
    \sr[4]_i_17 ,
    \sr[4]_i_17_0 ,
    \iv[10]_i_2 ,
    \tr[27]_i_3_0 ,
    \sr[4]_i_16_0 ,
    \sr[4]_i_16_1 ,
    \tr[21]_i_3_0 ,
    \sr[4]_i_33_0 ,
    \sr[4]_i_16_2 ,
    \tr[21]_i_3_1 ,
    \tr[20]_i_3_0 ,
    \sr[4]_i_39 ,
    \sr[4]_i_39_0 ,
    \iv[8]_i_2 ,
    \sr[4]_i_40 ,
    \sr[4]_i_80_0 ,
    \sr[4]_i_37 ,
    \tr[26]_i_3_0 ,
    \tr[24]_i_2 ,
    \tr[24]_i_3_0 ,
    \tr[24]_i_3_1 ,
    \tr[24]_i_3_2 ,
    \tr[30]_i_3_1 ,
    \tr[23]_i_2_0 ,
    \tr[23]_i_2_1 ,
    \tr[23]_i_3_0 ,
    \tr[23]_i_3_1 ,
    \tr[17]_i_2 ,
    \tr[17]_i_3_2 ,
    \tr[21]_i_2_0 ,
    \tr[21]_i_3_2 ,
    \tr[21]_i_3_3 ,
    \tr[22]_i_2 ,
    \tr[20]_i_2 ,
    \tr[20]_i_3_1 ,
    \tr[20]_i_3_2 ,
    \sr[4]_i_4_0 ,
    \tr[26]_i_2 ,
    \tr[26]_i_3_1 ,
    \tr[26]_i_3_2 ,
    \tr[29]_i_3_1 ,
    \tr[18]_i_2 ,
    \tr[18]_i_3_1 ,
    \tr[18]_i_3_2 ,
    \tr[27]_i_2_0 ,
    \tr[27]_i_3_1 ,
    \tr[28]_i_2_0 ,
    \tr[28]_i_2_1 ,
    \tr[28]_i_3_0 ,
    \tr[25]_i_2 ,
    \tr[25]_i_3_0 ,
    \tr[25]_i_3_1 ,
    \tr[19]_i_2_0 ,
    \tr[19]_i_3_2 ,
    \tr[19]_i_3_3 ,
    \iv[15]_i_8 ,
    \iv[15]_i_8_0 ,
    \iv[15]_i_8_1 ,
    \iv[15]_i_8_2 ,
    \tr[19]_i_3_4 ,
    \tr[19]_i_3_5 ,
    \tr[25]_i_3_2 ,
    \tr[18]_i_3_3 ,
    \tr[29]_i_3_2 ,
    \tr[17]_i_3_3 ,
    \tr[30]_i_3_2 ,
    \tr[24]_i_3_3 ,
    \tr[30]_i_3_3 ,
    \tr[30]_i_3_4 ,
    \tr[23]_i_3_2 ,
    \tr[26]_i_3_3 ,
    \tr[26]_i_3_4 ,
    \tr[29]_i_3_3 ,
    \tr[27]_i_3_2 ,
    \sr[4]_i_16_3 ,
    \iv[7]_i_3 ,
    \sr[4]_i_36_0 ,
    \sr[4]_i_19_0 ,
    \sr[4]_i_21_5 ,
    \iv[10]_i_2_0 ,
    \sr[4]_i_16_4 ,
    \sr[4]_i_16_5 ,
    \iv[9]_i_2 ,
    \tr[25]_i_3_3 ,
    \iv[0]_i_3_1 ,
    \tr[24]_i_10_1 ,
    \tr[25]_i_10_0 ,
    \iv[0]_i_10_0 ,
    \tr[16]_i_2_0 ,
    \iv[1]_i_10 ,
    \iv[1]_i_10_0 ,
    \iv[1]_i_10_1 ,
    \iv[3]_i_10 ,
    \iv[3]_i_10_0 ,
    \iv[3]_i_10_1 ,
    \sr[4]_i_45_0 ,
    \sr[4]_i_44_1 ,
    \sr[4]_i_35_0 ,
    \iv[6]_i_10 ,
    \iv[6]_i_10_0 ,
    \iv[6]_i_10_1 ,
    \iv[15]_i_22_0 ,
    \iv[0]_i_10_1 ,
    \sr[6]_i_12_0 ,
    \sr[6]_i_12_1 ,
    \sr[6]_i_12_2 ,
    \tr[16]_i_6_2 ,
    \tr[16]_i_6_3 ,
    \iv[7]_i_9 ,
    \sr[4]_i_43_1 ,
    \iv[1]_i_9 ,
    \iv[2]_i_9 ,
    \iv[3]_i_9 ,
    \sr[4]_i_45_1 ,
    \sr[4]_i_44_2 ,
    \iv[0]_i_8 ,
    \iv[0]_i_8_0 ,
    \iv[10]_i_5 ,
    \iv[5]_i_9 ,
    \iv[4]_i_9 ,
    \iv[8]_i_5 ,
    \sr[7]_i_7 ,
    \iv[14]_i_5 ,
    \iv[9]_i_5 ,
    \sr[4]_i_38_0 ,
    \tr[21]_i_3_4 ,
    \tr[22]_i_3_0 ,
    \tr[22]_i_3_1 ,
    \tr[20]_i_3_3 ,
    \iv[0]_i_10_2 ,
    \iv[0]_i_10_3 ,
    \sr[6]_i_11 ,
    \sr[6]_i_11_0 ,
    \sr[4]_i_38_1 ,
    \sr[4]_i_53_0 ,
    \sr[4]_i_58_0 ,
    \sr[4]_i_104_0 ,
    \sr[4]_i_108_0 ,
    \sr[4]_i_41_0 ,
    \sr[4]_i_85_0 ,
    \iv[0]_i_19 ,
    \iv[7]_i_3_0 ,
    \iv[7]_i_3_1 ,
    \sr[4]_i_76_0 ,
    \iv[0]_i_22_0 ,
    \sr[4]_i_75 ,
    \tr[29]_i_8_0 ,
    \iv[12]_i_13 ,
    \iv[5]_i_30 ,
    \iv[2]_i_24 ,
    \tr[22]_i_8_0 ,
    \iv[6]_i_15 ,
    \iv[10]_i_22_0 ,
    \iv[13]_i_26 ,
    \iv[13]_i_26_0 ,
    \tr[30]_i_9_0 ,
    \iv[13]_i_13 ,
    \iv[5]_i_14 ,
    \sr[4]_i_152 ,
    \tr[28]_i_6_0 ,
    \sr[4]_i_88 ,
    \iv[11]_i_13 ,
    \iv[4]_i_31 ,
    \sr[4]_i_152_0 ,
    \iv[7]_i_17_0 ,
    \iv[11]_i_25 ,
    \iv[3]_i_31 ,
    \iv[10]_i_13 ,
    \tr[23]_i_6_0 ,
    \iv[15]_i_60_0 ,
    \iv[10]_i_25 ,
    \iv[0]_i_7 ,
    \abus_o[3] ,
    \niho_dsp_a[32] ,
    \niho_dsp_a[32]_0 ,
    \niho_dsp_a[32]_1 ,
    \tr[22]_i_11 ,
    \iv[0]_i_6 ,
    \iv[0]_i_6_0 ,
    \iv[4]_i_6 ,
    \iv[8]_i_8 ,
    S,
    \mul_b_reg[5] ,
    \mul_b_reg[5]_0 ,
    \mul_b_reg[5]_1 ,
    \mul_b_reg[5]_2 ,
    \mul_b_reg[0] ,
    \mul_b_reg[0]_0 ,
    \mul_b_reg[0]_1 ,
    \mul_b_reg[0]_2 ,
    .abus_o_0_sp_1(abus_o_0_sn_1),
    \sr[4]_i_19_1 ,
    \sr[4]_i_19_2 ,
    \sr[4]_i_18 ,
    \sr[4]_i_18_0 ,
    \sr[4]_i_45_2 ,
    \sr[4]_i_61_0 ,
    \sr[6]_i_4 ,
    \iv[14]_i_32_0 ,
    \niho_dsp_a[16]_0 ,
    mul_rslt,
    mul_a,
    \tr[24]_i_3_4 ,
    \tr[24]_i_3_5 ,
    \sr[4]_i_64 ,
    \sr[4]_i_89_1 ,
    \iv[3]_i_15 ,
    \sr[4]_i_98_0 ,
    \tr[27]_i_6_0 ,
    \iv[9]_i_11_0 ,
    \sr[4]_i_67 ,
    \iv[10]_i_10_0 ,
    \iv[4]_i_14 ,
    \iv_reg[7]_i_12_0 ,
    abus_sel_0,
    bank_sel,
    bbus_sel_0,
    \i_/bdatw[15]_INST_0_i_65 ,
    ctl_selb_rn,
    \i_/bdatw[15]_INST_0_i_65_0 ,
    \i_/bdatw[15]_INST_0_i_65_1 ,
    ctl_selb_0,
    \i_/bdatw[15]_INST_0_i_65_2 ,
    \i_/badr[15]_INST_0_i_15 ,
    \badr[31]_INST_0_i_1 ,
    \badr[30]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1_0 ,
    \badr[31]_INST_0_i_1_0 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1_1 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1_1 ,
    SR,
    E,
    cbus,
    clk,
    \grn_reg[15]_10 ,
    \grn_reg[15]_11 ,
    \grn_reg[0]_5 ,
    \grn_reg[15]_12 ,
    \grn_reg[0]_6 ,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    \grn_reg[15]_15 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[0]_7 ,
    \grn_reg[15]_19 ,
    \grn_reg[0]_8 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 );
  output [5:0]p_2_in;
  output \badr[21]_INST_0_i_1 ;
  output \tr_reg[5] ;
  output \bdatw[8]_INST_0_i_2 ;
  output \tr_reg[0] ;
  output \iv[7]_i_33 ;
  output \sr_reg[8] ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr[4]_i_21_0 ;
  output \sr_reg[8]_2 ;
  output \iv[7]_i_37_0 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr[4]_i_147_0 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr[4]_i_65_0 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \iv[13]_i_27 ;
  output \sr_reg[8]_21 ;
  output \iv[8]_i_20 ;
  output \sr_reg[8]_22 ;
  output \iv[14]_i_35_0 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr[4]_i_116_0 ;
  output \sr_reg[8]_25 ;
  output \tr[17]_i_9_0 ;
  output \tr[24]_i_10_0 ;
  output \tr[30]_i_10_0 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \tr[20]_i_9_0 ;
  output \tr[22]_i_9_0 ;
  output \iv[12]_i_27_0 ;
  output \iv[13]_i_29_0 ;
  output \sr_reg[8]_28 ;
  output \tr[18]_i_9_0 ;
  output \tr[26]_i_9_0 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \iv[8]_i_30 ;
  output \sr_reg[8]_33 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \sr_reg[8]_36 ;
  output \iv[7]_i_17 ;
  output \iv[15]_i_94 ;
  output \sr_reg[8]_37 ;
  output \sr_reg[8]_38 ;
  output \iv[10]_i_10 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[8]_40 ;
  output \sr_reg[8]_41 ;
  output \iv[5]_i_23 ;
  output \sr_reg[8]_42 ;
  output \iv[9]_i_11 ;
  output \sr_reg[8]_43 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[8]_45 ;
  output \sr_reg[8]_46 ;
  output \sr_reg[8]_47 ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output \sr_reg[8]_50 ;
  output \sr_reg[8]_51 ;
  output \sr_reg[8]_52 ;
  output \tr[16]_i_9_0 ;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output \sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output \sr_reg[8]_57 ;
  output \sr_reg[8]_58 ;
  output \sr_reg[8]_59 ;
  output \sr_reg[8]_60 ;
  output \sr_reg[8]_61 ;
  output \sr_reg[8]_62 ;
  output \sr_reg[8]_63 ;
  output \sr_reg[8]_64 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output \sr_reg[8]_67 ;
  output \sr_reg[8]_68 ;
  output \sr_reg[8]_69 ;
  output \sr_reg[8]_70 ;
  output \sr_reg[8]_71 ;
  output \sr_reg[8]_72 ;
  output \sr_reg[8]_73 ;
  output \sr_reg[8]_74 ;
  output \sr_reg[8]_75 ;
  output \sr_reg[8]_76 ;
  output \sr_reg[8]_77 ;
  output \sr_reg[8]_78 ;
  output \sr_reg[8]_79 ;
  output \sr_reg[8]_80 ;
  output \sr_reg[8]_81 ;
  output \sr_reg[8]_82 ;
  output \sr_reg[8]_83 ;
  output \sr_reg[8]_84 ;
  output \sr_reg[8]_85 ;
  output \iv[7]_i_25 ;
  output \sr_reg[8]_86 ;
  output \sr_reg[8]_87 ;
  output \sr_reg[8]_88 ;
  output \sr_reg[8]_89 ;
  output \sr_reg[8]_90 ;
  output \sr_reg[8]_91 ;
  output \sr_reg[6] ;
  output \sr_reg[8]_92 ;
  output \badr[14]_INST_0_i_1 ;
  output \sr_reg[8]_93 ;
  output \sr_reg[6]_0 ;
  output \badr[0]_INST_0_i_1 ;
  output \iv[0]_i_25 ;
  output \badr[15]_INST_0_i_1 ;
  output \sr_reg[8]_94 ;
  output \sr_reg[8]_95 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[8]_96 ;
  output \sr_reg[8]_97 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[8]_98 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[6]_4 ;
  output \sr_reg[8]_99 ;
  output \sr_reg[8]_100 ;
  output \iv[14]_i_49 ;
  output \sr_reg[8]_101 ;
  output \sr_reg[8]_102 ;
  output \badr[14]_INST_0_i_1_0 ;
  output \sr_reg[8]_103 ;
  output \sr_reg[8]_104 ;
  output \sr_reg[8]_105 ;
  output \badr[0]_INST_0_i_1_0 ;
  output \badr[16]_INST_0_i_1 ;
  output \sr_reg[8]_106 ;
  output \sr_reg[8]_107 ;
  output \sr_reg[8]_108 ;
  output \sr_reg[8]_109 ;
  output \sr_reg[8]_110 ;
  output \sr_reg[6]_5 ;
  output \sr_reg[8]_111 ;
  output \sr_reg[8]_112 ;
  output \sr_reg[8]_113 ;
  output \sr_reg[6]_6 ;
  output \sr_reg[8]_114 ;
  output \sr_reg[8]_115 ;
  output \sr_reg[8]_116 ;
  output \sr_reg[8]_117 ;
  output \sr_reg[8]_118 ;
  output \sr_reg[6]_7 ;
  output \sr_reg[8]_119 ;
  output \badr[5]_INST_0_i_1 ;
  output \niho_dsp_a[15]_INST_0_i_3 ;
  output \sr_reg[8]_120 ;
  output [15:0]p_0_in;
  output [15:0]p_1_in;
  output \iv[15]_i_108 ;
  output \iv[15]_i_108_0 ;
  output \iv[15]_i_108_1 ;
  output \iv[15]_i_108_2 ;
  output \iv[15]_i_108_3 ;
  output \iv[15]_i_108_4 ;
  output \iv[15]_i_108_5 ;
  output \iv[15]_i_108_6 ;
  output \iv[15]_i_108_7 ;
  output \iv[15]_i_108_8 ;
  output \sr[4]_i_51_0 ;
  output [3:0]\art/add/iv[7]_i_32 ;
  output [3:0]\art/add/sr[5]_i_14 ;
  output [3:0]\sr_reg[6]_8 ;
  output [3:0]\art/add/sr[5]_i_18 ;
  output [0:0]CO;
  output [15:0]abus_o;
  output [1:0]bbus_o;
  output \sr_reg[8]_121 ;
  output \sr_reg[8]_122 ;
  output \sr_reg[8]_123 ;
  output \sr_reg[8]_124 ;
  output \sr_reg[8]_125 ;
  output \sr_reg[8]_126 ;
  output \sr_reg[6]_9 ;
  output \sr_reg[8]_127 ;
  output \sr_reg[6]_10 ;
  output \sr_reg[6]_11 ;
  output [16:0]niho_dsp_a;
  output \sr_reg[8]_128 ;
  output \sr_reg[8]_129 ;
  output \sr_reg[8]_130 ;
  output \sr_reg[8]_131 ;
  output \sr_reg[8]_132 ;
  output \grn_reg[15]_6 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_9 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  input \tr_reg[27] ;
  input [5:0]niho_dsp_c;
  input \tr_reg[23] ;
  input \tr_reg[23]_0 ;
  input \tr_reg[29] ;
  input \tr_reg[29]_0 ;
  input \tr_reg[28] ;
  input \tr_reg[28]_0 ;
  input \tr_reg[21] ;
  input \tr_reg[21]_0 ;
  input \tr_reg[19] ;
  input \tr_reg[19]_0 ;
  input \tr_reg[27]_0 ;
  input \tr_reg[27]_1 ;
  input [3:0]DI;
  input [3:0]bbus_0;
  input \iv[13]_i_17 ;
  input \iv[13]_i_17_0 ;
  input \iv[13]_i_17_1 ;
  input \tr[17]_i_3_0 ;
  input [3:0]\abus_o[11] ;
  input \sr[4]_i_36 ;
  input [3:0]\abus_o[7] ;
  input \iv[7]_i_7 ;
  input \iv[7]_i_7_0 ;
  input \iv[7]_i_7_1 ;
  input \tr_reg[1] ;
  input \tr_reg[16] ;
  input \tr_reg[1]_0 ;
  input [3:0]\niho_dsp_a[16] ;
  input \tr[16]_i_6_0 ;
  input \tr[16]_i_6_1 ;
  input \sr_reg[4] ;
  input \sr_reg[4]_0 ;
  input \sr[4]_i_5_0 ;
  input \sr[4]_i_5_1 ;
  input \sr[4]_i_5_2 ;
  input \sr[4]_i_42 ;
  input \tr[23]_i_7_0 ;
  input \sr[4]_i_89_0 ;
  input \sr[4]_i_43 ;
  input \sr[4]_i_43_0 ;
  input \tr[17]_i_3_1 ;
  input \sr[4]_i_5_3 ;
  input \sr[4]_i_21_1 ;
  input \tr[18]_i_3_0 ;
  input \sr[4]_i_21_2 ;
  input \sr[4]_i_21_3 ;
  input \sr[4]_i_21_4 ;
  input \tr[19]_i_3_0 ;
  input \tr[19]_i_3_1 ;
  input \sr[4]_i_5_4 ;
  input \sr[4]_i_5_5 ;
  input \sr[4]_i_20_0 ;
  input \sr[4]_i_20_1 ;
  input \iv[13]_i_2 ;
  input \tr[30]_i_3_0 ;
  input \sr[4]_i_20_2 ;
  input \sr[4]_i_20_3 ;
  input \iv[12]_i_2 ;
  input \tr[29]_i_3_0 ;
  input \sr[4]_i_44_0 ;
  input \iv[0]_i_3 ;
  input \iv[0]_i_3_0 ;
  input \sr[4]_i_17 ;
  input \sr[4]_i_17_0 ;
  input \iv[10]_i_2 ;
  input \tr[27]_i_3_0 ;
  input \sr[4]_i_16_0 ;
  input \sr[4]_i_16_1 ;
  input \tr[21]_i_3_0 ;
  input \sr[4]_i_33_0 ;
  input \sr[4]_i_16_2 ;
  input \tr[21]_i_3_1 ;
  input \tr[20]_i_3_0 ;
  input \sr[4]_i_39 ;
  input \sr[4]_i_39_0 ;
  input \iv[8]_i_2 ;
  input \sr[4]_i_40 ;
  input \sr[4]_i_80_0 ;
  input \sr[4]_i_37 ;
  input \tr[26]_i_3_0 ;
  input \tr[24]_i_2 ;
  input \tr[24]_i_3_0 ;
  input \tr[24]_i_3_1 ;
  input \tr[24]_i_3_2 ;
  input \tr[30]_i_3_1 ;
  input \tr[23]_i_2_0 ;
  input \tr[23]_i_2_1 ;
  input \tr[23]_i_3_0 ;
  input \tr[23]_i_3_1 ;
  input \tr[17]_i_2 ;
  input \tr[17]_i_3_2 ;
  input \tr[21]_i_2_0 ;
  input \tr[21]_i_3_2 ;
  input \tr[21]_i_3_3 ;
  input \tr[22]_i_2 ;
  input \tr[20]_i_2 ;
  input \tr[20]_i_3_1 ;
  input \tr[20]_i_3_2 ;
  input \sr[4]_i_4_0 ;
  input \tr[26]_i_2 ;
  input \tr[26]_i_3_1 ;
  input \tr[26]_i_3_2 ;
  input \tr[29]_i_3_1 ;
  input \tr[18]_i_2 ;
  input \tr[18]_i_3_1 ;
  input \tr[18]_i_3_2 ;
  input \tr[27]_i_2_0 ;
  input \tr[27]_i_3_1 ;
  input \tr[28]_i_2_0 ;
  input \tr[28]_i_2_1 ;
  input \tr[28]_i_3_0 ;
  input \tr[25]_i_2 ;
  input \tr[25]_i_3_0 ;
  input \tr[25]_i_3_1 ;
  input \tr[19]_i_2_0 ;
  input \tr[19]_i_3_2 ;
  input \tr[19]_i_3_3 ;
  input \iv[15]_i_8 ;
  input \iv[15]_i_8_0 ;
  input \iv[15]_i_8_1 ;
  input \iv[15]_i_8_2 ;
  input \tr[19]_i_3_4 ;
  input \tr[19]_i_3_5 ;
  input \tr[25]_i_3_2 ;
  input \tr[18]_i_3_3 ;
  input \tr[29]_i_3_2 ;
  input \tr[17]_i_3_3 ;
  input \tr[30]_i_3_2 ;
  input \tr[24]_i_3_3 ;
  input \tr[30]_i_3_3 ;
  input \tr[30]_i_3_4 ;
  input \tr[23]_i_3_2 ;
  input \tr[26]_i_3_3 ;
  input \tr[26]_i_3_4 ;
  input \tr[29]_i_3_3 ;
  input \tr[27]_i_3_2 ;
  input \sr[4]_i_16_3 ;
  input \iv[7]_i_3 ;
  input \sr[4]_i_36_0 ;
  input \sr[4]_i_19_0 ;
  input \sr[4]_i_21_5 ;
  input \iv[10]_i_2_0 ;
  input \sr[4]_i_16_4 ;
  input \sr[4]_i_16_5 ;
  input \iv[9]_i_2 ;
  input \tr[25]_i_3_3 ;
  input \iv[0]_i_3_1 ;
  input \tr[24]_i_10_1 ;
  input \tr[25]_i_10_0 ;
  input \iv[0]_i_10_0 ;
  input \tr[16]_i_2_0 ;
  input \iv[1]_i_10 ;
  input \iv[1]_i_10_0 ;
  input \iv[1]_i_10_1 ;
  input \iv[3]_i_10 ;
  input \iv[3]_i_10_0 ;
  input \iv[3]_i_10_1 ;
  input \sr[4]_i_45_0 ;
  input \sr[4]_i_44_1 ;
  input \sr[4]_i_35_0 ;
  input \iv[6]_i_10 ;
  input \iv[6]_i_10_0 ;
  input \iv[6]_i_10_1 ;
  input \iv[15]_i_22_0 ;
  input \iv[0]_i_10_1 ;
  input \sr[6]_i_12_0 ;
  input \sr[6]_i_12_1 ;
  input \sr[6]_i_12_2 ;
  input \tr[16]_i_6_2 ;
  input \tr[16]_i_6_3 ;
  input \iv[7]_i_9 ;
  input \sr[4]_i_43_1 ;
  input \iv[1]_i_9 ;
  input \iv[2]_i_9 ;
  input \iv[3]_i_9 ;
  input \sr[4]_i_45_1 ;
  input \sr[4]_i_44_2 ;
  input \iv[0]_i_8 ;
  input \iv[0]_i_8_0 ;
  input \iv[10]_i_5 ;
  input \iv[5]_i_9 ;
  input \iv[4]_i_9 ;
  input \iv[8]_i_5 ;
  input \sr[7]_i_7 ;
  input \iv[14]_i_5 ;
  input \iv[9]_i_5 ;
  input \sr[4]_i_38_0 ;
  input \tr[21]_i_3_4 ;
  input \tr[22]_i_3_0 ;
  input \tr[22]_i_3_1 ;
  input \tr[20]_i_3_3 ;
  input \iv[0]_i_10_2 ;
  input \iv[0]_i_10_3 ;
  input \sr[6]_i_11 ;
  input \sr[6]_i_11_0 ;
  input \sr[4]_i_38_1 ;
  input \sr[4]_i_53_0 ;
  input \sr[4]_i_58_0 ;
  input \sr[4]_i_104_0 ;
  input \sr[4]_i_108_0 ;
  input \sr[4]_i_41_0 ;
  input \sr[4]_i_85_0 ;
  input \iv[0]_i_19 ;
  input \iv[7]_i_3_0 ;
  input \iv[7]_i_3_1 ;
  input \sr[4]_i_76_0 ;
  input \iv[0]_i_22_0 ;
  input \sr[4]_i_75 ;
  input \tr[29]_i_8_0 ;
  input \iv[12]_i_13 ;
  input \iv[5]_i_30 ;
  input \iv[2]_i_24 ;
  input \tr[22]_i_8_0 ;
  input \iv[6]_i_15 ;
  input \iv[10]_i_22_0 ;
  input \iv[13]_i_26 ;
  input \iv[13]_i_26_0 ;
  input \tr[30]_i_9_0 ;
  input \iv[13]_i_13 ;
  input \iv[5]_i_14 ;
  input \sr[4]_i_152 ;
  input \tr[28]_i_6_0 ;
  input \sr[4]_i_88 ;
  input \iv[11]_i_13 ;
  input \iv[4]_i_31 ;
  input \sr[4]_i_152_0 ;
  input \iv[7]_i_17_0 ;
  input \iv[11]_i_25 ;
  input \iv[3]_i_31 ;
  input \iv[10]_i_13 ;
  input \tr[23]_i_6_0 ;
  input \iv[15]_i_60_0 ;
  input \iv[10]_i_25 ;
  input \iv[0]_i_7 ;
  input [3:0]\abus_o[3] ;
  input \niho_dsp_a[32] ;
  input \niho_dsp_a[32]_0 ;
  input \niho_dsp_a[32]_1 ;
  input \tr[22]_i_11 ;
  input \iv[0]_i_6 ;
  input [2:0]\iv[0]_i_6_0 ;
  input [2:0]\iv[4]_i_6 ;
  input [3:0]\iv[8]_i_8 ;
  input [3:0]S;
  input \mul_b_reg[5] ;
  input \mul_b_reg[5]_0 ;
  input \mul_b_reg[5]_1 ;
  input \mul_b_reg[5]_2 ;
  input \mul_b_reg[0] ;
  input \mul_b_reg[0]_0 ;
  input \mul_b_reg[0]_1 ;
  input \mul_b_reg[0]_2 ;
  input \sr[4]_i_19_1 ;
  input \sr[4]_i_19_2 ;
  input \sr[4]_i_18 ;
  input \sr[4]_i_18_0 ;
  input \sr[4]_i_45_2 ;
  input \sr[4]_i_61_0 ;
  input \sr[6]_i_4 ;
  input \iv[14]_i_32_0 ;
  input \niho_dsp_a[16]_0 ;
  input mul_rslt;
  input [16:0]mul_a;
  input \tr[24]_i_3_4 ;
  input \tr[24]_i_3_5 ;
  input \sr[4]_i_64 ;
  input \sr[4]_i_89_1 ;
  input \iv[3]_i_15 ;
  input \sr[4]_i_98_0 ;
  input \tr[27]_i_6_0 ;
  input \iv[9]_i_11_0 ;
  input \sr[4]_i_67 ;
  input \iv[10]_i_10_0 ;
  input \iv[4]_i_14 ;
  input \iv_reg[7]_i_12_0 ;
  input [7:0]abus_sel_0;
  input [0:0]bank_sel;
  input [5:0]bbus_sel_0;
  input \i_/bdatw[15]_INST_0_i_65 ;
  input [1:0]ctl_selb_rn;
  input \i_/bdatw[15]_INST_0_i_65_0 ;
  input \i_/bdatw[15]_INST_0_i_65_1 ;
  input [0:0]ctl_selb_0;
  input \i_/bdatw[15]_INST_0_i_65_2 ;
  input \i_/badr[15]_INST_0_i_15 ;
  input \badr[31]_INST_0_i_1 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1_0 ;
  input \badr[31]_INST_0_i_1_0 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1_1 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1_1 ;
  input [0:0]SR;
  input [0:0]E;
  input [15:0]cbus;
  input clk;
  input [0:0]\grn_reg[15]_10 ;
  input [0:0]\grn_reg[15]_11 ;
  input [0:0]\grn_reg[0]_5 ;
  input [0:0]\grn_reg[15]_12 ;
  input [0:0]\grn_reg[0]_6 ;
  input [0:0]\grn_reg[15]_13 ;
  input [0:0]\grn_reg[15]_14 ;
  input [0:0]\grn_reg[15]_15 ;
  input [15:0]\grn_reg[15]_16 ;
  input [0:0]\grn_reg[15]_17 ;
  input [0:0]\grn_reg[15]_18 ;
  input [0:0]\grn_reg[0]_7 ;
  input [0:0]\grn_reg[15]_19 ;
  input [0:0]\grn_reg[0]_8 ;
  input [0:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
     output [15:0]gr20;
     output [15:0]gr21;
     output [15:0]gr22;
     output [15:0]gr23;
     output [15:0]gr24;
     output [15:0]gr25;
     output [15:0]gr26;
     output [15:0]gr27;
  input abus_o_0_sn_1;

  wire \<const0> ;
  wire [0:0]CO;
  wire [3:0]DI;
  wire [0:0]E;
  wire [3:0]S;
  wire [0:0]SR;
  wire [15:0]abus_o;
  wire [3:0]\abus_o[11] ;
  wire [3:0]\abus_o[3] ;
  wire [3:0]\abus_o[7] ;
  wire abus_o_0_sn_1;
  wire [7:0]abus_sel_0;
  wire \art/add/iv[3]_i_26_n_0 ;
  wire \art/add/iv[7]_i_31_n_0 ;
  wire [3:0]\art/add/iv[7]_i_32 ;
  wire [3:0]\art/add/sr[5]_i_14 ;
  wire [3:0]\art/add/sr[5]_i_18 ;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[0]_INST_0_i_1_0 ;
  wire \badr[14]_INST_0_i_1 ;
  wire \badr[14]_INST_0_i_1_0 ;
  wire \badr[15]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[16]_INST_0_i_1_1 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1_1 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire \badr[31]_INST_0_i_1 ;
  wire \badr[31]_INST_0_i_1_0 ;
  wire \badr[5]_INST_0_i_1 ;
  wire [0:0]bank_sel;
  wire [3:0]bbus_0;
  wire [1:0]bbus_o;
  wire [5:0]bbus_sel_0;
  wire bbuso2l_n_10;
  wire bbuso2l_n_16;
  wire bbuso_n_10;
  wire bbuso_n_16;
  wire \bdatw[8]_INST_0_i_2 ;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire grn27_n_10;
  wire grn27_n_11;
  wire grn27_n_13;
  wire grn27_n_15;
  wire grn27_n_20;
  wire grn27_n_22;
  wire grn27_n_27;
  wire grn27_n_3;
  wire grn27_n_30;
  wire grn27_n_33;
  wire grn27_n_37;
  wire grn27_n_44;
  wire grn27_n_57;
  wire grn27_n_58;
  wire grn27_n_7;
  wire grn27_n_8;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire [0:0]\grn_reg[0]_5 ;
  wire [0:0]\grn_reg[0]_6 ;
  wire [0:0]\grn_reg[0]_7 ;
  wire [0:0]\grn_reg[0]_8 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire [0:0]\grn_reg[15]_10 ;
  wire [0:0]\grn_reg[15]_11 ;
  wire [0:0]\grn_reg[15]_12 ;
  wire [0:0]\grn_reg[15]_13 ;
  wire [0:0]\grn_reg[15]_14 ;
  wire [0:0]\grn_reg[15]_15 ;
  wire [15:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [0:0]\grn_reg[15]_18 ;
  wire [0:0]\grn_reg[15]_19 ;
  wire [0:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \i_/badr[15]_INST_0_i_15 ;
  wire \i_/bdatw[15]_INST_0_i_65 ;
  wire \i_/bdatw[15]_INST_0_i_65_0 ;
  wire \i_/bdatw[15]_INST_0_i_65_1 ;
  wire \i_/bdatw[15]_INST_0_i_65_2 ;
  wire \iv[0]_i_10_0 ;
  wire \iv[0]_i_10_1 ;
  wire \iv[0]_i_10_2 ;
  wire \iv[0]_i_10_3 ;
  wire \iv[0]_i_17_n_0 ;
  wire \iv[0]_i_18_n_0 ;
  wire \iv[0]_i_19 ;
  wire \iv[0]_i_21_n_0 ;
  wire \iv[0]_i_22_0 ;
  wire \iv[0]_i_22_n_0 ;
  wire \iv[0]_i_23_n_0 ;
  wire \iv[0]_i_25 ;
  wire \iv[0]_i_3 ;
  wire \iv[0]_i_30_n_0 ;
  wire \iv[0]_i_3_0 ;
  wire \iv[0]_i_3_1 ;
  wire \iv[0]_i_6 ;
  wire [2:0]\iv[0]_i_6_0 ;
  wire \iv[0]_i_7 ;
  wire \iv[0]_i_8 ;
  wire \iv[0]_i_8_0 ;
  wire \iv[10]_i_10 ;
  wire \iv[10]_i_10_0 ;
  wire \iv[10]_i_13 ;
  wire \iv[10]_i_2 ;
  wire \iv[10]_i_22_0 ;
  wire \iv[10]_i_24_n_0 ;
  wire \iv[10]_i_25 ;
  wire \iv[10]_i_2_0 ;
  wire \iv[10]_i_35_n_0 ;
  wire \iv[10]_i_38_n_0 ;
  wire \iv[10]_i_39_n_0 ;
  wire \iv[10]_i_45_n_0 ;
  wire \iv[10]_i_5 ;
  wire \iv[11]_i_13 ;
  wire \iv[11]_i_25 ;
  wire \iv[11]_i_26_n_0 ;
  wire \iv[11]_i_30_n_0 ;
  wire \iv[11]_i_31_n_0 ;
  wire \iv[12]_i_13 ;
  wire \iv[12]_i_2 ;
  wire \iv[12]_i_25_n_0 ;
  wire \iv[12]_i_27_0 ;
  wire \iv[12]_i_29_n_0 ;
  wire \iv[12]_i_30_n_0 ;
  wire \iv[12]_i_35_n_0 ;
  wire \iv[12]_i_50_n_0 ;
  wire \iv[13]_i_13 ;
  wire \iv[13]_i_17 ;
  wire \iv[13]_i_17_0 ;
  wire \iv[13]_i_17_1 ;
  wire \iv[13]_i_2 ;
  wire \iv[13]_i_25_n_0 ;
  wire \iv[13]_i_26 ;
  wire \iv[13]_i_26_0 ;
  wire \iv[13]_i_27 ;
  wire \iv[13]_i_29_0 ;
  wire \iv[13]_i_31_n_0 ;
  wire \iv[13]_i_32_n_0 ;
  wire \iv[13]_i_36_n_0 ;
  wire \iv[13]_i_37_n_0 ;
  wire \iv[14]_i_32_0 ;
  wire \iv[14]_i_35_0 ;
  wire \iv[14]_i_42_n_0 ;
  wire \iv[14]_i_43_n_0 ;
  wire \iv[14]_i_44_n_0 ;
  wire \iv[14]_i_45_n_0 ;
  wire \iv[14]_i_46_n_0 ;
  wire \iv[14]_i_47_n_0 ;
  wire \iv[14]_i_48_n_0 ;
  wire \iv[14]_i_49 ;
  wire \iv[14]_i_5 ;
  wire \iv[14]_i_57_n_0 ;
  wire \iv[14]_i_59_n_0 ;
  wire \iv[14]_i_60_n_0 ;
  wire \iv[14]_i_61_n_0 ;
  wire \iv[14]_i_62_n_0 ;
  wire \iv[14]_i_63_n_0 ;
  wire \iv[14]_i_64_n_0 ;
  wire \iv[15]_i_104_n_0 ;
  wire \iv[15]_i_106_n_0 ;
  wire \iv[15]_i_108 ;
  wire \iv[15]_i_108_0 ;
  wire \iv[15]_i_108_1 ;
  wire \iv[15]_i_108_2 ;
  wire \iv[15]_i_108_3 ;
  wire \iv[15]_i_108_4 ;
  wire \iv[15]_i_108_5 ;
  wire \iv[15]_i_108_6 ;
  wire \iv[15]_i_108_7 ;
  wire \iv[15]_i_108_8 ;
  wire \iv[15]_i_149_n_0 ;
  wire \iv[15]_i_150_n_0 ;
  wire \iv[15]_i_151_n_0 ;
  wire \iv[15]_i_152_n_0 ;
  wire \iv[15]_i_153_n_0 ;
  wire \iv[15]_i_154_n_0 ;
  wire \iv[15]_i_155_n_0 ;
  wire \iv[15]_i_157_n_0 ;
  wire \iv[15]_i_22_0 ;
  wire \iv[15]_i_55_n_0 ;
  wire \iv[15]_i_60_0 ;
  wire \iv[15]_i_60_n_0 ;
  wire \iv[15]_i_8 ;
  wire \iv[15]_i_8_0 ;
  wire \iv[15]_i_8_1 ;
  wire \iv[15]_i_8_2 ;
  wire \iv[15]_i_94 ;
  wire \iv[1]_i_10 ;
  wire \iv[1]_i_10_0 ;
  wire \iv[1]_i_10_1 ;
  wire \iv[1]_i_18_n_0 ;
  wire \iv[1]_i_25_n_0 ;
  wire \iv[1]_i_9 ;
  wire \iv[2]_i_17_n_0 ;
  wire \iv[2]_i_24 ;
  wire \iv[2]_i_26_n_0 ;
  wire \iv[2]_i_31_n_0 ;
  wire \iv[2]_i_9 ;
  wire \iv[3]_i_10 ;
  wire \iv[3]_i_10_0 ;
  wire \iv[3]_i_10_1 ;
  wire \iv[3]_i_15 ;
  wire \iv[3]_i_18_n_0 ;
  wire \iv[3]_i_30_n_0 ;
  wire \iv[3]_i_31 ;
  wire \iv[3]_i_9 ;
  wire \iv[4]_i_14 ;
  wire \iv[4]_i_18_n_0 ;
  wire \iv[4]_i_31 ;
  wire \iv[4]_i_34_n_0 ;
  wire [2:0]\iv[4]_i_6 ;
  wire \iv[4]_i_9 ;
  wire \iv[5]_i_14 ;
  wire \iv[5]_i_18_n_0 ;
  wire \iv[5]_i_23 ;
  wire \iv[5]_i_28_n_0 ;
  wire \iv[5]_i_30 ;
  wire \iv[5]_i_33_n_0 ;
  wire \iv[5]_i_9 ;
  wire \iv[6]_i_10 ;
  wire \iv[6]_i_10_0 ;
  wire \iv[6]_i_10_1 ;
  wire \iv[6]_i_15 ;
  wire \iv[6]_i_29_n_0 ;
  wire \iv[6]_i_30_n_0 ;
  wire \iv[7]_i_17 ;
  wire \iv[7]_i_17_0 ;
  wire \iv[7]_i_25 ;
  wire \iv[7]_i_3 ;
  wire \iv[7]_i_33 ;
  wire \iv[7]_i_37_0 ;
  wire \iv[7]_i_37_n_0 ;
  wire \iv[7]_i_38_n_0 ;
  wire \iv[7]_i_3_0 ;
  wire \iv[7]_i_3_1 ;
  wire \iv[7]_i_43_n_0 ;
  wire \iv[7]_i_46_n_0 ;
  wire \iv[7]_i_7 ;
  wire \iv[7]_i_7_0 ;
  wire \iv[7]_i_7_1 ;
  wire \iv[7]_i_9 ;
  wire \iv[8]_i_2 ;
  wire \iv[8]_i_20 ;
  wire \iv[8]_i_26_n_0 ;
  wire \iv[8]_i_27_n_0 ;
  wire \iv[8]_i_30 ;
  wire \iv[8]_i_41_n_0 ;
  wire \iv[8]_i_5 ;
  wire [3:0]\iv[8]_i_8 ;
  wire \iv[9]_i_11 ;
  wire \iv[9]_i_11_0 ;
  wire \iv[9]_i_2 ;
  wire \iv[9]_i_28_n_0 ;
  wire \iv[9]_i_5 ;
  wire \iv[9]_i_51_n_0 ;
  wire \iv_reg[3]_i_11_n_0 ;
  wire \iv_reg[3]_i_11_n_1 ;
  wire \iv_reg[3]_i_11_n_2 ;
  wire \iv_reg[3]_i_11_n_3 ;
  wire \iv_reg[7]_i_12_0 ;
  wire \iv_reg[7]_i_12_n_0 ;
  wire \iv_reg[7]_i_12_n_1 ;
  wire \iv_reg[7]_i_12_n_2 ;
  wire \iv_reg[7]_i_12_n_3 ;
  wire [16:0]mul_a;
  wire \mul_b_reg[0] ;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[0]_1 ;
  wire \mul_b_reg[0]_2 ;
  wire \mul_b_reg[5] ;
  wire \mul_b_reg[5]_0 ;
  wire \mul_b_reg[5]_1 ;
  wire \mul_b_reg[5]_2 ;
  wire mul_rslt;
  wire [16:0]niho_dsp_a;
  wire \niho_dsp_a[15]_INST_0_i_3 ;
  wire [3:0]\niho_dsp_a[16] ;
  wire \niho_dsp_a[16]_0 ;
  wire \niho_dsp_a[32] ;
  wire \niho_dsp_a[32]_0 ;
  wire \niho_dsp_a[32]_1 ;
  wire [5:0]niho_dsp_c;
  wire [15:0]p_0_in;
  wire [15:0]p_1_in;
  wire [5:0]p_2_in;
  wire \sr[4]_i_101_n_0 ;
  wire \sr[4]_i_102_n_0 ;
  wire \sr[4]_i_104_0 ;
  wire \sr[4]_i_104_n_0 ;
  wire \sr[4]_i_106_n_0 ;
  wire \sr[4]_i_107_n_0 ;
  wire \sr[4]_i_108_0 ;
  wire \sr[4]_i_108_n_0 ;
  wire \sr[4]_i_110_n_0 ;
  wire \sr[4]_i_113_n_0 ;
  wire \sr[4]_i_114_n_0 ;
  wire \sr[4]_i_116_0 ;
  wire \sr[4]_i_118_n_0 ;
  wire \sr[4]_i_122_n_0 ;
  wire \sr[4]_i_127_n_0 ;
  wire \sr[4]_i_12_n_0 ;
  wire \sr[4]_i_134_n_0 ;
  wire \sr[4]_i_13_n_0 ;
  wire \sr[4]_i_142_n_0 ;
  wire \sr[4]_i_147_0 ;
  wire \sr[4]_i_149_n_0 ;
  wire \sr[4]_i_14_n_0 ;
  wire \sr[4]_i_152 ;
  wire \sr[4]_i_152_0 ;
  wire \sr[4]_i_159_n_0 ;
  wire \sr[4]_i_15_n_0 ;
  wire \sr[4]_i_162_n_0 ;
  wire \sr[4]_i_168_n_0 ;
  wire \sr[4]_i_16_0 ;
  wire \sr[4]_i_16_1 ;
  wire \sr[4]_i_16_2 ;
  wire \sr[4]_i_16_3 ;
  wire \sr[4]_i_16_4 ;
  wire \sr[4]_i_16_5 ;
  wire \sr[4]_i_16_n_0 ;
  wire \sr[4]_i_17 ;
  wire \sr[4]_i_17_0 ;
  wire \sr[4]_i_18 ;
  wire \sr[4]_i_18_0 ;
  wire \sr[4]_i_19_0 ;
  wire \sr[4]_i_19_1 ;
  wire \sr[4]_i_19_2 ;
  wire \sr[4]_i_19_n_0 ;
  wire \sr[4]_i_20_0 ;
  wire \sr[4]_i_20_1 ;
  wire \sr[4]_i_20_2 ;
  wire \sr[4]_i_20_3 ;
  wire \sr[4]_i_20_n_0 ;
  wire \sr[4]_i_21_0 ;
  wire \sr[4]_i_21_1 ;
  wire \sr[4]_i_21_2 ;
  wire \sr[4]_i_21_3 ;
  wire \sr[4]_i_21_4 ;
  wire \sr[4]_i_21_5 ;
  wire \sr[4]_i_21_n_0 ;
  wire \sr[4]_i_31_n_0 ;
  wire \sr[4]_i_32_n_0 ;
  wire \sr[4]_i_33_0 ;
  wire \sr[4]_i_33_n_0 ;
  wire \sr[4]_i_34_n_0 ;
  wire \sr[4]_i_35_0 ;
  wire \sr[4]_i_36 ;
  wire \sr[4]_i_36_0 ;
  wire \sr[4]_i_37 ;
  wire \sr[4]_i_38_0 ;
  wire \sr[4]_i_38_1 ;
  wire \sr[4]_i_39 ;
  wire \sr[4]_i_39_0 ;
  wire \sr[4]_i_40 ;
  wire \sr[4]_i_41_0 ;
  wire \sr[4]_i_41_n_0 ;
  wire \sr[4]_i_42 ;
  wire \sr[4]_i_43 ;
  wire \sr[4]_i_43_0 ;
  wire \sr[4]_i_43_1 ;
  wire \sr[4]_i_44_0 ;
  wire \sr[4]_i_44_1 ;
  wire \sr[4]_i_44_2 ;
  wire \sr[4]_i_44_n_0 ;
  wire \sr[4]_i_45_0 ;
  wire \sr[4]_i_45_1 ;
  wire \sr[4]_i_45_2 ;
  wire \sr[4]_i_45_n_0 ;
  wire \sr[4]_i_46_n_0 ;
  wire \sr[4]_i_47_n_0 ;
  wire \sr[4]_i_4_0 ;
  wire \sr[4]_i_50_n_0 ;
  wire \sr[4]_i_51_0 ;
  wire \sr[4]_i_51_n_0 ;
  wire \sr[4]_i_52_n_0 ;
  wire \sr[4]_i_53_0 ;
  wire \sr[4]_i_53_n_0 ;
  wire \sr[4]_i_55_n_0 ;
  wire \sr[4]_i_56_n_0 ;
  wire \sr[4]_i_57_n_0 ;
  wire \sr[4]_i_58_0 ;
  wire \sr[4]_i_58_n_0 ;
  wire \sr[4]_i_5_0 ;
  wire \sr[4]_i_5_1 ;
  wire \sr[4]_i_5_2 ;
  wire \sr[4]_i_5_3 ;
  wire \sr[4]_i_5_4 ;
  wire \sr[4]_i_5_5 ;
  wire \sr[4]_i_60_n_0 ;
  wire \sr[4]_i_61_0 ;
  wire \sr[4]_i_61_n_0 ;
  wire \sr[4]_i_62_n_0 ;
  wire \sr[4]_i_63_n_0 ;
  wire \sr[4]_i_64 ;
  wire \sr[4]_i_65_0 ;
  wire \sr[4]_i_65_n_0 ;
  wire \sr[4]_i_67 ;
  wire \sr[4]_i_70_n_0 ;
  wire \sr[4]_i_71_n_0 ;
  wire \sr[4]_i_72_n_0 ;
  wire \sr[4]_i_75 ;
  wire \sr[4]_i_76_0 ;
  wire \sr[4]_i_80_0 ;
  wire \sr[4]_i_82_n_0 ;
  wire \sr[4]_i_83_n_0 ;
  wire \sr[4]_i_85_0 ;
  wire \sr[4]_i_85_n_0 ;
  wire \sr[4]_i_88 ;
  wire \sr[4]_i_89_0 ;
  wire \sr[4]_i_89_1 ;
  wire \sr[4]_i_95_n_0 ;
  wire \sr[4]_i_97_n_0 ;
  wire \sr[4]_i_98_0 ;
  wire \sr[4]_i_98_n_0 ;
  wire \sr[4]_i_99_n_0 ;
  wire \sr[6]_i_11 ;
  wire \sr[6]_i_11_0 ;
  wire \sr[6]_i_12_0 ;
  wire \sr[6]_i_12_1 ;
  wire \sr[6]_i_12_2 ;
  wire \sr[6]_i_27_n_0 ;
  wire \sr[6]_i_28_n_0 ;
  wire \sr[6]_i_35_n_0 ;
  wire \sr[6]_i_39_n_0 ;
  wire \sr[6]_i_4 ;
  wire \sr[6]_i_40_n_0 ;
  wire \sr[7]_i_17_n_0 ;
  wire \sr[7]_i_34_n_0 ;
  wire \sr[7]_i_35_n_0 ;
  wire \sr[7]_i_36_n_0 ;
  wire \sr[7]_i_41_n_0 ;
  wire \sr[7]_i_42_n_0 ;
  wire \sr[7]_i_43_n_0 ;
  wire \sr[7]_i_7 ;
  wire \sr_reg[4] ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[5]_i_10_n_0 ;
  wire \sr_reg[5]_i_10_n_1 ;
  wire \sr_reg[5]_i_10_n_2 ;
  wire \sr_reg[5]_i_10_n_3 ;
  wire \sr_reg[5]_i_5_n_1 ;
  wire \sr_reg[5]_i_5_n_2 ;
  wire \sr_reg[5]_i_5_n_3 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_10 ;
  wire \sr_reg[6]_11 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_7 ;
  wire [3:0]\sr_reg[6]_8 ;
  wire \sr_reg[6]_9 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_100 ;
  wire \sr_reg[8]_101 ;
  wire \sr_reg[8]_102 ;
  wire \sr_reg[8]_103 ;
  wire \sr_reg[8]_104 ;
  wire \sr_reg[8]_105 ;
  wire \sr_reg[8]_106 ;
  wire \sr_reg[8]_107 ;
  wire \sr_reg[8]_108 ;
  wire \sr_reg[8]_109 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_110 ;
  wire \sr_reg[8]_111 ;
  wire \sr_reg[8]_112 ;
  wire \sr_reg[8]_113 ;
  wire \sr_reg[8]_114 ;
  wire \sr_reg[8]_115 ;
  wire \sr_reg[8]_116 ;
  wire \sr_reg[8]_117 ;
  wire \sr_reg[8]_118 ;
  wire \sr_reg[8]_119 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_120 ;
  wire \sr_reg[8]_121 ;
  wire \sr_reg[8]_122 ;
  wire \sr_reg[8]_123 ;
  wire \sr_reg[8]_124 ;
  wire \sr_reg[8]_125 ;
  wire \sr_reg[8]_126 ;
  wire \sr_reg[8]_127 ;
  wire \sr_reg[8]_128 ;
  wire \sr_reg[8]_129 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_130 ;
  wire \sr_reg[8]_131 ;
  wire \sr_reg[8]_132 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_51 ;
  wire \sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire \sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire \sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_60 ;
  wire \sr_reg[8]_61 ;
  wire \sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire \sr_reg[8]_71 ;
  wire \sr_reg[8]_72 ;
  wire \sr_reg[8]_73 ;
  wire \sr_reg[8]_74 ;
  wire \sr_reg[8]_75 ;
  wire \sr_reg[8]_76 ;
  wire \sr_reg[8]_77 ;
  wire \sr_reg[8]_78 ;
  wire \sr_reg[8]_79 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_80 ;
  wire \sr_reg[8]_81 ;
  wire \sr_reg[8]_82 ;
  wire \sr_reg[8]_83 ;
  wire \sr_reg[8]_84 ;
  wire \sr_reg[8]_85 ;
  wire \sr_reg[8]_86 ;
  wire \sr_reg[8]_87 ;
  wire \sr_reg[8]_88 ;
  wire \sr_reg[8]_89 ;
  wire \sr_reg[8]_9 ;
  wire \sr_reg[8]_90 ;
  wire \sr_reg[8]_91 ;
  wire \sr_reg[8]_92 ;
  wire \sr_reg[8]_93 ;
  wire \sr_reg[8]_94 ;
  wire \sr_reg[8]_95 ;
  wire \sr_reg[8]_96 ;
  wire \sr_reg[8]_97 ;
  wire \sr_reg[8]_98 ;
  wire \sr_reg[8]_99 ;
  wire \tr[16]_i_12_n_0 ;
  wire \tr[16]_i_13_n_0 ;
  wire \tr[16]_i_16_n_0 ;
  wire \tr[16]_i_17_n_0 ;
  wire \tr[16]_i_24_n_0 ;
  wire \tr[16]_i_26_n_0 ;
  wire \tr[16]_i_28_n_0 ;
  wire \tr[16]_i_2_0 ;
  wire \tr[16]_i_32_n_0 ;
  wire \tr[16]_i_5_n_0 ;
  wire \tr[16]_i_6_0 ;
  wire \tr[16]_i_6_1 ;
  wire \tr[16]_i_6_2 ;
  wire \tr[16]_i_6_3 ;
  wire \tr[16]_i_6_n_0 ;
  wire \tr[16]_i_9_0 ;
  wire \tr[17]_i_16_n_0 ;
  wire \tr[17]_i_2 ;
  wire \tr[17]_i_3_0 ;
  wire \tr[17]_i_3_1 ;
  wire \tr[17]_i_3_2 ;
  wire \tr[17]_i_3_3 ;
  wire \tr[17]_i_6_n_0 ;
  wire \tr[17]_i_7_n_0 ;
  wire \tr[17]_i_9_0 ;
  wire \tr[17]_i_9_n_0 ;
  wire \tr[18]_i_2 ;
  wire \tr[18]_i_3_0 ;
  wire \tr[18]_i_3_1 ;
  wire \tr[18]_i_3_2 ;
  wire \tr[18]_i_3_3 ;
  wire \tr[18]_i_7_n_0 ;
  wire \tr[18]_i_8_n_0 ;
  wire \tr[18]_i_9_0 ;
  wire \tr[18]_i_9_n_0 ;
  wire \tr[19]_i_2_0 ;
  wire \tr[19]_i_3_0 ;
  wire \tr[19]_i_3_1 ;
  wire \tr[19]_i_3_2 ;
  wire \tr[19]_i_3_3 ;
  wire \tr[19]_i_3_4 ;
  wire \tr[19]_i_3_5 ;
  wire \tr[19]_i_3_n_0 ;
  wire \tr[19]_i_6_n_0 ;
  wire \tr[19]_i_7_n_0 ;
  wire \tr[19]_i_9_n_0 ;
  wire \tr[20]_i_16_n_0 ;
  wire \tr[20]_i_19_n_0 ;
  wire \tr[20]_i_2 ;
  wire \tr[20]_i_3_0 ;
  wire \tr[20]_i_3_1 ;
  wire \tr[20]_i_3_2 ;
  wire \tr[20]_i_3_3 ;
  wire \tr[20]_i_7_n_0 ;
  wire \tr[20]_i_8_n_0 ;
  wire \tr[20]_i_9_0 ;
  wire \tr[20]_i_9_n_0 ;
  wire \tr[21]_i_15_n_0 ;
  wire \tr[21]_i_2_0 ;
  wire \tr[21]_i_3_0 ;
  wire \tr[21]_i_3_1 ;
  wire \tr[21]_i_3_2 ;
  wire \tr[21]_i_3_3 ;
  wire \tr[21]_i_3_4 ;
  wire \tr[21]_i_3_n_0 ;
  wire \tr[21]_i_7_n_0 ;
  wire \tr[21]_i_8_n_0 ;
  wire \tr[21]_i_9_n_0 ;
  wire \tr[22]_i_11 ;
  wire \tr[22]_i_2 ;
  wire \tr[22]_i_3_0 ;
  wire \tr[22]_i_3_1 ;
  wire \tr[22]_i_6_n_0 ;
  wire \tr[22]_i_8_0 ;
  wire \tr[22]_i_8_n_0 ;
  wire \tr[22]_i_9_0 ;
  wire \tr[22]_i_9_n_0 ;
  wire \tr[23]_i_10_n_0 ;
  wire \tr[23]_i_2_0 ;
  wire \tr[23]_i_2_1 ;
  wire \tr[23]_i_3_0 ;
  wire \tr[23]_i_3_1 ;
  wire \tr[23]_i_3_2 ;
  wire \tr[23]_i_3_n_0 ;
  wire \tr[23]_i_6_0 ;
  wire \tr[23]_i_6_n_0 ;
  wire \tr[23]_i_7_0 ;
  wire \tr[23]_i_7_n_0 ;
  wire \tr[24]_i_10_0 ;
  wire \tr[24]_i_10_1 ;
  wire \tr[24]_i_10_n_0 ;
  wire \tr[24]_i_2 ;
  wire \tr[24]_i_3_0 ;
  wire \tr[24]_i_3_1 ;
  wire \tr[24]_i_3_2 ;
  wire \tr[24]_i_3_3 ;
  wire \tr[24]_i_3_4 ;
  wire \tr[24]_i_3_5 ;
  wire \tr[24]_i_6_n_0 ;
  wire \tr[24]_i_7_n_0 ;
  wire \tr[24]_i_9_n_0 ;
  wire \tr[25]_i_10_0 ;
  wire \tr[25]_i_10_n_0 ;
  wire \tr[25]_i_2 ;
  wire \tr[25]_i_3_0 ;
  wire \tr[25]_i_3_1 ;
  wire \tr[25]_i_3_2 ;
  wire \tr[25]_i_3_3 ;
  wire \tr[25]_i_6_n_0 ;
  wire \tr[25]_i_7_n_0 ;
  wire \tr[25]_i_9_n_0 ;
  wire \tr[26]_i_2 ;
  wire \tr[26]_i_3_0 ;
  wire \tr[26]_i_3_1 ;
  wire \tr[26]_i_3_2 ;
  wire \tr[26]_i_3_3 ;
  wire \tr[26]_i_3_4 ;
  wire \tr[26]_i_6_n_0 ;
  wire \tr[26]_i_7_n_0 ;
  wire \tr[26]_i_9_0 ;
  wire \tr[26]_i_9_n_0 ;
  wire \tr[27]_i_2_0 ;
  wire \tr[27]_i_3_0 ;
  wire \tr[27]_i_3_1 ;
  wire \tr[27]_i_3_2 ;
  wire \tr[27]_i_3_n_0 ;
  wire \tr[27]_i_6_0 ;
  wire \tr[27]_i_6_n_0 ;
  wire \tr[27]_i_7_n_0 ;
  wire \tr[27]_i_9_n_0 ;
  wire \tr[28]_i_2_0 ;
  wire \tr[28]_i_2_1 ;
  wire \tr[28]_i_3_0 ;
  wire \tr[28]_i_3_n_0 ;
  wire \tr[28]_i_6_0 ;
  wire \tr[28]_i_6_n_0 ;
  wire \tr[28]_i_7_n_0 ;
  wire \tr[29]_i_3_0 ;
  wire \tr[29]_i_3_1 ;
  wire \tr[29]_i_3_2 ;
  wire \tr[29]_i_3_3 ;
  wire \tr[29]_i_3_n_0 ;
  wire \tr[29]_i_6_n_0 ;
  wire \tr[29]_i_7_n_0 ;
  wire \tr[29]_i_8_0 ;
  wire \tr[29]_i_8_n_0 ;
  wire \tr[29]_i_9_n_0 ;
  wire \tr[30]_i_10_0 ;
  wire \tr[30]_i_10_n_0 ;
  wire \tr[30]_i_3_0 ;
  wire \tr[30]_i_3_1 ;
  wire \tr[30]_i_3_2 ;
  wire \tr[30]_i_3_3 ;
  wire \tr[30]_i_3_4 ;
  wire \tr[30]_i_7_n_0 ;
  wire \tr[30]_i_8_n_0 ;
  wire \tr[30]_i_9_0 ;
  wire \tr[30]_i_9_n_0 ;
  wire \tr_reg[0] ;
  wire \tr_reg[16] ;
  wire \tr_reg[19] ;
  wire \tr_reg[19]_0 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;
  wire \tr_reg[21] ;
  wire \tr_reg[21]_0 ;
  wire \tr_reg[23] ;
  wire \tr_reg[23]_0 ;
  wire \tr_reg[27] ;
  wire \tr_reg[27]_0 ;
  wire \tr_reg[27]_1 ;
  wire \tr_reg[28] ;
  wire \tr_reg[28]_0 ;
  wire \tr_reg[29] ;
  wire \tr_reg[29]_0 ;
  wire \tr_reg[5] ;

  GND GND
       (.G(\<const0> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[0]_INST_0 
       (.I0(\abus_o[3] [0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[10]_INST_0 
       (.I0(\abus_o[11] [2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[11]_INST_0 
       (.I0(\abus_o[11] [3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[12]_INST_0 
       (.I0(DI[0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[13]_INST_0 
       (.I0(DI[1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[14]_INST_0 
       (.I0(DI[2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[15]_INST_0 
       (.I0(DI[3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[15]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[1]_INST_0 
       (.I0(\abus_o[3] [1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[2]_INST_0 
       (.I0(\abus_o[3] [2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[3]_INST_0 
       (.I0(\abus_o[3] [3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[4]_INST_0 
       (.I0(\abus_o[7] [0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[5]_INST_0 
       (.I0(\abus_o[7] [1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[6]_INST_0 
       (.I0(\abus_o[7] [2]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[7]_INST_0 
       (.I0(\abus_o[7] [3]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[8]_INST_0 
       (.I0(\abus_o[11] [0]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[9]_INST_0 
       (.I0(\abus_o[11] [1]),
        .I1(abus_o_0_sn_1),
        .O(abus_o[9]));
  niho_rgf_bank_bus_22 abuso
       (.abus_sel_0(abus_sel_0),
        .bank_sel(bank_sel),
        .\i_/badr[15]_INST_0_i_10_0 ({\niho_dsp_a[16] [3],\niho_dsp_a[16] [1:0]}),
        .\i_/badr[15]_INST_0_i_11_0 (gr02),
        .\i_/badr[15]_INST_0_i_11_1 (gr01),
        .\i_/badr[15]_INST_0_i_3_0 (gr00),
        .\i_/badr[15]_INST_0_i_3_1 (gr07),
        .\i_/badr[15]_INST_0_i_3_2 (gr03),
        .\i_/badr[15]_INST_0_i_3_3 (gr04),
        .\mul_a_reg[15] (gr05),
        .out(gr06),
        .p_1_in(p_1_in));
  niho_rgf_bank_bus_23 abuso2h
       (.abus_sel_0({abus_sel_0[7],abus_sel_0[4:3],abus_sel_0[0]}),
        .\badr[16]_INST_0_i_1 (\badr[16]_INST_0_i_1_0 ),
        .\badr[16]_INST_0_i_1_0 (\badr[16]_INST_0_i_1_1 ),
        .\badr[17]_INST_0_i_1 (\badr[17]_INST_0_i_1 ),
        .\badr[17]_INST_0_i_1_0 (\badr[17]_INST_0_i_1_0 ),
        .\badr[18]_INST_0_i_1 (\badr[18]_INST_0_i_1 ),
        .\badr[18]_INST_0_i_1_0 (\badr[18]_INST_0_i_1_0 ),
        .\badr[19]_INST_0_i_1 (\badr[19]_INST_0_i_1 ),
        .\badr[19]_INST_0_i_1_0 (\badr[19]_INST_0_i_1_0 ),
        .\badr[20]_INST_0_i_1 (\badr[20]_INST_0_i_1 ),
        .\badr[20]_INST_0_i_1_0 (\badr[20]_INST_0_i_1_0 ),
        .\badr[21]_INST_0_i_1 (\badr[21]_INST_0_i_1_0 ),
        .\badr[21]_INST_0_i_1_0 (\badr[21]_INST_0_i_1_1 ),
        .\badr[22]_INST_0_i_1 (\badr[22]_INST_0_i_1 ),
        .\badr[22]_INST_0_i_1_0 (\badr[22]_INST_0_i_1_0 ),
        .\badr[23]_INST_0_i_1 (\badr[23]_INST_0_i_1 ),
        .\badr[23]_INST_0_i_1_0 (\badr[23]_INST_0_i_1_0 ),
        .\badr[24]_INST_0_i_1 (\badr[24]_INST_0_i_1 ),
        .\badr[24]_INST_0_i_1_0 (\badr[24]_INST_0_i_1_0 ),
        .\badr[25]_INST_0_i_1 (\badr[25]_INST_0_i_1 ),
        .\badr[25]_INST_0_i_1_0 (\badr[25]_INST_0_i_1_0 ),
        .\badr[26]_INST_0_i_1 (\badr[26]_INST_0_i_1 ),
        .\badr[26]_INST_0_i_1_0 (\badr[26]_INST_0_i_1_0 ),
        .\badr[27]_INST_0_i_1 (\badr[27]_INST_0_i_1 ),
        .\badr[27]_INST_0_i_1_0 (\badr[27]_INST_0_i_1_0 ),
        .\badr[28]_INST_0_i_1 (\badr[28]_INST_0_i_1 ),
        .\badr[28]_INST_0_i_1_0 (\badr[28]_INST_0_i_1_0 ),
        .\badr[29]_INST_0_i_1 (\badr[29]_INST_0_i_1 ),
        .\badr[29]_INST_0_i_1_0 (\badr[29]_INST_0_i_1_0 ),
        .\badr[30]_INST_0_i_1 (\badr[30]_INST_0_i_1 ),
        .\badr[30]_INST_0_i_1_0 (\badr[30]_INST_0_i_1_0 ),
        .\badr[31]_INST_0_i_1 (gr20),
        .\badr[31]_INST_0_i_1_0 (\badr[31]_INST_0_i_1 ),
        .\badr[31]_INST_0_i_1_1 (gr23),
        .\badr[31]_INST_0_i_1_2 (gr24),
        .\badr[31]_INST_0_i_1_3 (\badr[31]_INST_0_i_1_0 ),
        .\grn_reg[0] (\grn_reg[0]_3 ),
        .\grn_reg[0]_0 (\grn_reg[0]_4 ),
        .\grn_reg[10] (\grn_reg[10]_1 ),
        .\grn_reg[10]_0 (\grn_reg[10]_2 ),
        .\grn_reg[11] (\grn_reg[11]_1 ),
        .\grn_reg[11]_0 (\grn_reg[11]_2 ),
        .\grn_reg[12] (\grn_reg[12]_1 ),
        .\grn_reg[12]_0 (\grn_reg[12]_2 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[13]_0 (\grn_reg[13]_2 ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[14]_0 (\grn_reg[14]_2 ),
        .\grn_reg[15] (\grn_reg[15]_8 ),
        .\grn_reg[15]_0 (\grn_reg[15]_9 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[1]_0 (\grn_reg[1]_4 ),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[2]_0 (\grn_reg[2]_4 ),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[4] (\grn_reg[4]_3 ),
        .\grn_reg[4]_0 (\grn_reg[4]_4 ),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\grn_reg[6] (\grn_reg[6]_1 ),
        .\grn_reg[6]_0 (\grn_reg[6]_2 ),
        .\grn_reg[7] (\grn_reg[7]_1 ),
        .\grn_reg[7]_0 (\grn_reg[7]_2 ),
        .\grn_reg[8] (\grn_reg[8]_1 ),
        .\grn_reg[8]_0 (\grn_reg[8]_2 ),
        .\grn_reg[9] (\grn_reg[9]_1 ),
        .\grn_reg[9]_0 (\grn_reg[9]_2 ),
        .\i_/badr[31]_INST_0_i_5_0 ({\niho_dsp_a[16] [3],\niho_dsp_a[16] [0]}),
        .out(gr27));
  niho_rgf_bank_bus_24 abuso2l
       (.abus_sel_0(abus_sel_0),
        .\i_/badr[15]_INST_0_i_14_0 ({\niho_dsp_a[16] [3],\niho_dsp_a[16] [1:0]}),
        .\i_/badr[15]_INST_0_i_15_0 (gr22),
        .\i_/badr[15]_INST_0_i_15_1 (gr21),
        .\i_/badr[15]_INST_0_i_15_2 (\i_/badr[15]_INST_0_i_15 ),
        .\i_/badr[15]_INST_0_i_4_0 (gr27),
        .\i_/badr[15]_INST_0_i_4_1 (gr23),
        .\i_/badr[15]_INST_0_i_4_2 (gr24),
        .\mul_a_reg[15] (gr26),
        .\mul_a_reg[15]_0 (gr25),
        .out(gr20),
        .p_0_in(p_0_in));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[3]_i_26 
       (.I0(\abus_o[3] [0]),
        .I1(\iv_reg[7]_i_12_0 ),
        .I2(\tr_reg[0] ),
        .O(\art/add/iv[3]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'h69)) 
    \art/add/iv[7]_i_31 
       (.I0(\abus_o[7] [1]),
        .I1(\iv_reg[7]_i_12_0 ),
        .I2(\tr_reg[5] ),
        .O(\art/add/iv[7]_i_31_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[0]_INST_0 
       (.I0(\tr_reg[0] ),
        .I1(abus_o_0_sn_1),
        .O(bbus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \bbus_o[5]_INST_0 
       (.I0(\tr_reg[5] ),
        .I1(abus_o_0_sn_1),
        .O(bbus_o[1]));
  niho_rgf_bank_bus_25 bbuso
       (.bank_sel(bank_sel),
        .bbus_sel_0(bbus_sel_0),
        .\bdatw[15]_INST_0_i_8 (gr03),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .\grn_reg[0] (bbuso_n_16),
        .\grn_reg[0]_0 (\grn_reg[0] ),
        .\grn_reg[0]_1 (\grn_reg[0]_0 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[15] (\grn_reg[15]_6 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (\grn_reg[4]_0 ),
        .\grn_reg[5] (bbuso_n_10),
        .\grn_reg[5]_0 (\grn_reg[5] ),
        .\grn_reg[5]_1 (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\i_/bdatw[15]_INST_0_i_24_0 (gr07),
        .\i_/bdatw[15]_INST_0_i_24_1 (gr00),
        .\i_/bdatw[15]_INST_0_i_24_2 (gr02),
        .\i_/bdatw[15]_INST_0_i_24_3 (gr01),
        .\i_/bdatw[15]_INST_0_i_48_0 ({\niho_dsp_a[16] [3],\niho_dsp_a[16] [1:0]}),
        .\i_/bdatw[15]_INST_0_i_48_1 (gr06),
        .\i_/bdatw[15]_INST_0_i_48_2 (gr05),
        .\i_/bdatw[15]_INST_0_i_65_0 (\i_/bdatw[15]_INST_0_i_65 ),
        .\i_/bdatw[15]_INST_0_i_65_1 (\i_/bdatw[15]_INST_0_i_65_0 ),
        .\i_/bdatw[15]_INST_0_i_65_2 (\i_/bdatw[15]_INST_0_i_65_1 ),
        .\i_/bdatw[15]_INST_0_i_65_3 (\i_/bdatw[15]_INST_0_i_65_2 ),
        .out(gr04));
  niho_rgf_bank_bus_26 bbuso2l
       (.bbus_sel_0(bbus_sel_0),
        .\bdatw[15]_INST_0_i_8 (gr23),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .\grn_reg[0] (bbuso2l_n_16),
        .\grn_reg[0]_0 (\grn_reg[0]_1 ),
        .\grn_reg[0]_1 (\grn_reg[0]_2 ),
        .\grn_reg[10] (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14]_0 ),
        .\grn_reg[15] (\grn_reg[15]_7 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (\grn_reg[1]_2 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (\grn_reg[2]_2 ),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (\grn_reg[3]_2 ),
        .\grn_reg[4] (\grn_reg[4]_1 ),
        .\grn_reg[4]_0 (\grn_reg[4]_2 ),
        .\grn_reg[5] (bbuso2l_n_10),
        .\grn_reg[5]_0 (\grn_reg[5]_1 ),
        .\grn_reg[5]_1 (\grn_reg[5]_2 ),
        .\grn_reg[6] (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7]_0 ),
        .\grn_reg[8] (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9]_0 ),
        .\i_/bdatw[15]_INST_0_i_23_0 (gr27),
        .\i_/bdatw[15]_INST_0_i_23_1 (gr20),
        .\i_/bdatw[15]_INST_0_i_23_2 (gr22),
        .\i_/bdatw[15]_INST_0_i_23_3 (gr21),
        .\i_/bdatw[15]_INST_0_i_46_0 ({\niho_dsp_a[16] [3],\niho_dsp_a[16] [1:0]}),
        .\i_/bdatw[15]_INST_0_i_46_1 (gr26),
        .\i_/bdatw[15]_INST_0_i_46_2 (gr25),
        .\i_/bdatw[15]_INST_0_i_64_0 (\i_/badr[15]_INST_0_i_15 ),
        .\i_/bdatw[15]_INST_0_i_64_1 (\i_/bdatw[15]_INST_0_i_65_2 ),
        .\i_/bdatw[15]_INST_0_i_64_2 (\i_/bdatw[15]_INST_0_i_65_0 ),
        .\i_/bdatw[15]_INST_0_i_64_3 (\i_/bdatw[15]_INST_0_i_65_1 ),
        .\i_/bdatw[15]_INST_0_i_64_4 (\i_/bdatw[15]_INST_0_i_65 ),
        .out(gr24));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_1 
       (.I0(\mul_b_reg[5] ),
        .I1(\mul_b_reg[5]_0 ),
        .I2(\mul_b_reg[5]_1 ),
        .I3(bbuso_n_10),
        .I4(bbuso2l_n_10),
        .I5(\mul_b_reg[5]_2 ),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_1 
       (.I0(\mul_b_reg[0] ),
        .I1(\mul_b_reg[0]_0 ),
        .I2(\mul_b_reg[0]_1 ),
        .I3(bbuso_n_16),
        .I4(bbuso2l_n_16),
        .I5(\mul_b_reg[0]_2 ),
        .O(\tr_reg[0] ));
  niho_rgf_grn_27 grn00
       (.E(E),
        .Q(gr00),
        .SR(SR),
        .cbus(cbus),
        .clk(clk));
  niho_rgf_grn_28 grn01
       (.Q(gr01),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_10 ));
  niho_rgf_grn_29 grn02
       (.Q(gr02),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_11 ));
  niho_rgf_grn_30 grn03
       (.Q(gr03),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_5 ));
  niho_rgf_grn_31 grn04
       (.Q(gr04),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_12 ));
  niho_rgf_grn_32 grn05
       (.Q(gr05),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_6 ));
  niho_rgf_grn_33 grn06
       (.Q(gr06),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_13 ));
  niho_rgf_grn_34 grn07
       (.Q(gr07),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ));
  niho_rgf_grn_35 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_15 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ));
  niho_rgf_grn_36 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_17 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ));
  niho_rgf_grn_37 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_18 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ));
  niho_rgf_grn_38 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_7 ),
        .\grn_reg[15]_0 (\grn_reg[15]_16 ));
  niho_rgf_grn_39 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_19 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ));
  niho_rgf_grn_40 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_8 ),
        .\grn_reg[15]_0 (\grn_reg[15]_16 ));
  niho_rgf_grn_41 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_20 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ));
  niho_rgf_grn_42 grn27
       (.DI({DI[3],DI[1]}),
        .Q(gr27),
        .SR(SR),
        .\badr[5]_INST_0_i_1 (\badr[5]_INST_0_i_1 ),
        .bbus_0(bbus_0[2:1]),
        .\bdatw[12]_INST_0_i_1 (grn27_n_37),
        .\bdatw[12]_INST_0_i_1_0 (grn27_n_44),
        .\bdatw[8]_INST_0_i_2 (\bdatw[8]_INST_0_i_2 ),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_21 ),
        .\grn_reg[15]_1 (\grn_reg[15]_16 ),
        .\iv[0]_i_25 (\iv[0]_i_25 ),
        .\iv[0]_i_7 (\iv[13]_i_17 ),
        .\iv[0]_i_7_0 (\abus_o[11] [0]),
        .\iv[0]_i_7_1 (\iv[0]_i_7 ),
        .\iv[10]_i_10 (\iv[10]_i_10 ),
        .\iv[10]_i_2 (\iv[10]_i_2 ),
        .\iv[10]_i_2_0 (\sr[4]_i_17_0 ),
        .\iv[10]_i_2_1 (\sr_reg[8]_39 ),
        .\iv[10]_i_2_2 (\iv[10]_i_2_0 ),
        .\iv[10]_i_5_0 (\iv[10]_i_24_n_0 ),
        .\iv[10]_i_5_1 (\tr[27]_i_3_0 ),
        .\iv[10]_i_5_2 (\tr[26]_i_3_1 ),
        .\iv[10]_i_5_3 (\sr_reg[8]_32 ),
        .\iv[10]_i_5_4 (\iv[10]_i_5 ),
        .\iv[10]_i_6 (\sr[4]_i_35_0 ),
        .\iv[11]_i_18 (\iv[14]_i_63_n_0 ),
        .\iv[11]_i_18_0 (\iv[15]_i_155_n_0 ),
        .\iv[11]_i_2 (\sr[4]_i_43 ),
        .\iv[11]_i_5_0 (\sr[4]_i_43_0 ),
        .\iv[11]_i_5_1 (\iv[11]_i_26_n_0 ),
        .\iv[11]_i_5_2 (\iv[11]_i_30_n_0 ),
        .\iv[11]_i_5_3 (\iv[11]_i_31_n_0 ),
        .\iv[11]_i_5_4 (\sr[4]_i_43_1 ),
        .\iv[11]_i_6_0 (\sr_reg[8]_45 ),
        .\iv[12]_i_15 (\sr_reg[6] ),
        .\iv[12]_i_15_0 (\sr_reg[8]_116 ),
        .\iv[12]_i_2 (\iv[12]_i_2 ),
        .\iv[12]_i_21 (\badr[15]_INST_0_i_1 ),
        .\iv[12]_i_21_0 (\sr_reg[8]_93 ),
        .\iv[12]_i_21_1 (\iv[15]_i_149_n_0 ),
        .\iv[12]_i_2_0 (\sr[4]_i_20_3 ),
        .\iv[12]_i_5_0 (\tr[29]_i_3_0 ),
        .\iv[12]_i_5_1 (\iv[12]_i_25_n_0 ),
        .\iv[12]_i_5_2 (\iv[12]_i_29_n_0 ),
        .\iv[12]_i_5_3 (\iv[12]_i_30_n_0 ),
        .\iv[12]_i_5_4 (\sr[4]_i_44_2 ),
        .\iv[12]_i_6 (\sr[4]_i_44_1 ),
        .\iv[12]_i_9 (\sr[6]_i_12_2 ),
        .\iv[13]_i_15 (\sr_reg[6]_2 ),
        .\iv[13]_i_15_0 (\sr_reg[8]_96 ),
        .\iv[13]_i_2 (\iv[13]_i_2 ),
        .\iv[13]_i_2_0 (\sr[4]_i_20_1 ),
        .\iv[13]_i_5_0 (\iv[13]_i_25_n_0 ),
        .\iv[13]_i_5_1 (\tr[30]_i_3_0 ),
        .\iv[13]_i_5_2 (\iv[13]_i_31_n_0 ),
        .\iv[13]_i_5_3 (\iv[13]_i_32_n_0 ),
        .\iv[13]_i_5_4 (\sr[4]_i_45_1 ),
        .\iv[13]_i_6 (\sr[4]_i_45_0 ),
        .\iv[14]_i_19 (\abus_o[3] [0]),
        .\iv[14]_i_2 (\sr[4]_i_40 ),
        .\iv[14]_i_49 (\iv[14]_i_49 ),
        .\iv[14]_i_5_0 (\iv[14]_i_35_0 ),
        .\iv[14]_i_5_1 (\sr[4]_i_80_0 ),
        .\iv[14]_i_5_2 (\sr_reg[8]_27 ),
        .\iv[14]_i_5_3 (\sr[7]_i_7 ),
        .\iv[14]_i_5_4 (\iv[14]_i_5 ),
        .\iv[14]_i_6 (\sr_reg[8]_73 ),
        .\iv[15]_i_94 (\iv[15]_i_94 ),
        .\iv[1]_i_10_0 (\iv[1]_i_10 ),
        .\iv[1]_i_10_1 (\iv[1]_i_10_0 ),
        .\iv[1]_i_10_2 (\iv[1]_i_10_1 ),
        .\iv[1]_i_10_3 (\sr_reg[8]_84 ),
        .\iv[1]_i_15 (grn27_n_7),
        .\iv[1]_i_15_0 (\sr_reg[8]_61 ),
        .\iv[1]_i_20_0 (\sr_reg[8]_97 ),
        .\iv[1]_i_23_0 (\sr[4]_i_152 ),
        .\iv[1]_i_23_1 (\badr[14]_INST_0_i_1_0 ),
        .\iv[1]_i_32 (\iv[14]_i_64_n_0 ),
        .\iv[1]_i_3_0 (\iv[1]_i_18_n_0 ),
        .\iv[1]_i_9_0 (\iv[1]_i_25_n_0 ),
        .\iv[1]_i_9_1 (\tr[17]_i_3_1 ),
        .\iv[1]_i_9_2 (\tr[17]_i_3_2 ),
        .\iv[1]_i_9_3 (\sr_reg[8]_30 ),
        .\iv[1]_i_9_4 (\iv[1]_i_9 ),
        .\iv[2]_i_10_0 (\iv[10]_i_35_n_0 ),
        .\iv[2]_i_10_1 (\iv[2]_i_31_n_0 ),
        .\iv[2]_i_15 (grn27_n_10),
        .\iv[2]_i_15_0 (\sr_reg[8]_80 ),
        .\iv[2]_i_15_1 (\iv[10]_i_38_n_0 ),
        .\iv[2]_i_15_2 (\iv[10]_i_39_n_0 ),
        .\iv[2]_i_26 (grn27_n_11),
        .\iv[2]_i_3_0 (\iv[2]_i_17_n_0 ),
        .\iv[2]_i_9_0 (\tr[18]_i_3_1 ),
        .\iv[2]_i_9_1 (\sr_reg[8]_33 ),
        .\iv[2]_i_9_2 (\iv[2]_i_9 ),
        .\iv[3]_i_10_0 (\iv[3]_i_10 ),
        .\iv[3]_i_10_1 (\iv[3]_i_10_0 ),
        .\iv[3]_i_10_2 (\iv[3]_i_10_1 ),
        .\iv[3]_i_15 (\sr_reg[8]_59 ),
        .\iv[3]_i_15_0 (\iv[3]_i_15 ),
        .\iv[3]_i_20 (\iv[0]_i_19 ),
        .\iv[3]_i_3 (\iv[3]_i_18_n_0 ),
        .\iv[3]_i_3_0 (\sr[4]_i_21_3 ),
        .\iv[3]_i_9_0 (\tr[19]_i_3_2 ),
        .\iv[3]_i_9_1 (\sr_reg[8]_28 ),
        .\iv[3]_i_9_2 (\iv[3]_i_9 ),
        .\iv[4]_i_10_0 (\iv[12]_i_35_n_0 ),
        .\iv[4]_i_10_1 (\iv[0]_i_10_0 ),
        .\iv[4]_i_10_2 (\iv[4]_i_34_n_0 ),
        .\iv[4]_i_14 (\iv[13]_i_36_n_0 ),
        .\iv[4]_i_14_0 (\sr[4]_i_89_0 ),
        .\iv[4]_i_14_1 (\iv[4]_i_14 ),
        .\iv[4]_i_17_0 (\tr[20]_i_16_n_0 ),
        .\iv[4]_i_29 (grn27_n_22),
        .\iv[4]_i_3 (\iv[4]_i_18_n_0 ),
        .\iv[4]_i_9_0 (\tr[20]_i_3_1 ),
        .\iv[4]_i_9_1 (\iv[12]_i_27_0 ),
        .\iv[4]_i_9_2 (\iv[4]_i_9 ),
        .\iv[5]_i_10_0 (\iv[13]_i_37_n_0 ),
        .\iv[5]_i_10_1 (\sr_reg[8]_77 ),
        .\iv[5]_i_10_2 (\iv[5]_i_33_n_0 ),
        .\iv[5]_i_14 (\iv[5]_i_14 ),
        .\iv[5]_i_23 (\iv[5]_i_23 ),
        .\iv[5]_i_28 (grn27_n_20),
        .\iv[5]_i_3 (\iv[5]_i_18_n_0 ),
        .\iv[5]_i_3_0 (\sr[4]_i_16_0 ),
        .\iv[5]_i_7 (\tr_reg[5] ),
        .\iv[5]_i_9_0 (\tr[21]_i_3_2 ),
        .\iv[5]_i_9_1 (\iv[13]_i_29_0 ),
        .\iv[5]_i_9_2 (\iv[5]_i_9 ),
        .\iv[6]_i_10 (\iv[6]_i_10 ),
        .\iv[6]_i_10_0 (\iv[6]_i_10_0 ),
        .\iv[6]_i_10_1 (\iv[6]_i_10_1 ),
        .\iv[6]_i_15 (\sr_reg[8]_52 ),
        .\iv[6]_i_15_0 (\iv[6]_i_15 ),
        .\iv[6]_i_9 (\tr[16]_i_6_2 ),
        .\iv[6]_i_9_0 (\iv[6]_i_29_n_0 ),
        .\iv[6]_i_9_1 (\iv[6]_i_30_n_0 ),
        .\iv[6]_i_9_2 (\sr[4]_i_38_0 ),
        .\iv[7]_i_17 (\iv[7]_i_17 ),
        .\iv[7]_i_17_0 (\sr_reg[8]_55 ),
        .\iv[7]_i_17_1 (\iv[7]_i_17_0 ),
        .\iv[7]_i_25 (\iv[7]_i_25 ),
        .\iv[7]_i_3 (\iv[7]_i_3 ),
        .\iv[7]_i_33 (\iv[7]_i_33 ),
        .\iv[7]_i_3_0 (\iv[7]_i_3_0 ),
        .\iv[7]_i_3_1 (\iv[7]_i_3_1 ),
        .\iv[7]_i_7 ({\abus_o[7] [3],\abus_o[7] [1]}),
        .\iv[7]_i_7_0 (\iv[7]_i_7 ),
        .\iv[7]_i_7_1 (\iv[7]_i_7_0 ),
        .\iv[7]_i_7_2 (\iv[7]_i_7_1 ),
        .\iv[7]_i_9_0 (\iv[7]_i_37_n_0 ),
        .\iv[7]_i_9_1 (\iv[7]_i_38_n_0 ),
        .\iv[7]_i_9_2 (\tr[23]_i_3_0 ),
        .\iv[7]_i_9_3 (\iv[7]_i_9 ),
        .\iv[7]_i_9_4 (\sr[6]_i_11_0 ),
        .\iv[8]_i_10 (\sr_reg[8]_48 ),
        .\iv[8]_i_10_0 (\iv[0]_i_8 ),
        .\iv[8]_i_2 (\sr[4]_i_39 ),
        .\iv[8]_i_2_0 (\iv[8]_i_2 ),
        .\iv[8]_i_5_0 (\sr_reg[8]_1 ),
        .\iv[8]_i_5_1 (\iv[8]_i_26_n_0 ),
        .\iv[8]_i_5_2 (\iv[8]_i_27_n_0 ),
        .\iv[8]_i_5_3 (\tr[24]_i_3_0 ),
        .\iv[8]_i_5_4 (\iv[8]_i_30 ),
        .\iv[8]_i_5_5 (\iv[8]_i_5 ),
        .\iv[8]_i_6_0 (\sr_reg[8]_49 ),
        .\iv[8]_i_6_1 (\sr_reg[8]_91 ),
        .\iv[8]_i_9 (\tr[17]_i_3_0 ),
        .\iv[9]_i_11 (\iv[9]_i_11 ),
        .\iv[9]_i_11_0 (\iv[9]_i_11_0 ),
        .\iv[9]_i_2 (\sr[4]_i_37 ),
        .\iv[9]_i_2_0 (\sr[4]_i_16_3 ),
        .\iv[9]_i_2_1 (\iv[9]_i_2 ),
        .\iv[9]_i_36 (grn27_n_27),
        .\iv[9]_i_4_0 (\sr[4]_i_36 ),
        .\iv[9]_i_4_1 (\sr_reg[8]_3 ),
        .\iv[9]_i_4_2 (\sr[4]_i_36_0 ),
        .\iv[9]_i_4_3 (\tr[30]_i_3_4 ),
        .\iv[9]_i_5_0 (\tr[26]_i_3_0 ),
        .\iv[9]_i_5_1 (\iv[9]_i_28_n_0 ),
        .\iv[9]_i_5_2 (\tr[25]_i_3_0 ),
        .\iv[9]_i_5_3 (\sr_reg[8]_29 ),
        .\iv[9]_i_5_4 (\iv[9]_i_5 ),
        .\niho_dsp_a[15]_INST_0_i_3 (\niho_dsp_a[15]_INST_0_i_3 ),
        .\niho_dsp_a[32] (\niho_dsp_a[16] [3:2]),
        .\niho_dsp_a[32]_0 (\niho_dsp_a[32] ),
        .\niho_dsp_a[32]_1 (\niho_dsp_a[32]_0 ),
        .\niho_dsp_a[32]_2 (\niho_dsp_a[32]_1 ),
        .p_0_in(p_0_in[15]),
        .p_1_in(p_1_in[15]),
        .\sr[4]_i_114 (\sr[7]_i_36_n_0 ),
        .\sr[4]_i_114_0 (\badr[14]_INST_0_i_1 ),
        .\sr[4]_i_135 (\badr[0]_INST_0_i_1 ),
        .\sr[4]_i_135_0 (\iv[14]_i_48_n_0 ),
        .\sr[4]_i_135_1 (\iv[14]_i_46_n_0 ),
        .\sr[4]_i_135_2 (\iv[14]_i_47_n_0 ),
        .\sr[4]_i_146 (\tr_reg[0] ),
        .\sr[4]_i_146_0 (\sr[7]_i_41_n_0 ),
        .\sr[4]_i_146_1 (\iv[14]_i_45_n_0 ),
        .\sr[4]_i_19 (\sr[4]_i_19_0 ),
        .\sr[4]_i_21 (\sr[4]_i_21_5 ),
        .\sr[4]_i_31 (\tr[21]_i_3_1 ),
        .\sr[4]_i_31_0 (\tr[20]_i_3_0 ),
        .\sr[4]_i_31_1 (\sr_reg[8]_76 ),
        .\sr[4]_i_33 (\tr[21]_i_3_0 ),
        .\sr[4]_i_33_0 (\sr[4]_i_33_0 ),
        .\sr[4]_i_33_1 (\iv[5]_i_28_n_0 ),
        .\sr[4]_i_46 (\iv[3]_i_30_n_0 ),
        .\sr[4]_i_46_0 (\tr[19]_i_3_0 ),
        .\sr[4]_i_46_1 (\tr[19]_i_3_1 ),
        .\sr[4]_i_47 (\tr[18]_i_3_0 ),
        .\sr[4]_i_47_0 (\iv[2]_i_26_n_0 ),
        .\sr[4]_i_82 (\iv[13]_i_17_0 ),
        .\sr[4]_i_88 (\sr[4]_i_88 ),
        .\sr[4]_i_88_0 (\iv[7]_i_43_n_0 ),
        .\sr[7]_i_20 (grn27_n_3),
        .\sr_reg[6] (grn27_n_58),
        .\sr_reg[6]_0 (\sr_reg[6]_10 ),
        .\sr_reg[6]_1 (\sr_reg[6]_9 ),
        .\sr_reg[6]_2 (\sr_reg[6]_11 ),
        .\sr_reg[6]_3 (\sr_reg[6]_6 ),
        .\sr_reg[8] (\sr_reg[8]_2 ),
        .\sr_reg[8]_0 (\sr_reg[8]_5 ),
        .\sr_reg[8]_1 (\sr_reg[8]_7 ),
        .\sr_reg[8]_10 (\sr_reg[8]_14 ),
        .\sr_reg[8]_11 (\sr_reg[8]_16 ),
        .\sr_reg[8]_12 (\sr_reg[8]_18 ),
        .\sr_reg[8]_13 (\sr_reg[8]_19 ),
        .\sr_reg[8]_14 (\sr_reg[8]_20 ),
        .\sr_reg[8]_15 (\sr_reg[8]_21 ),
        .\sr_reg[8]_16 (\sr_reg[8]_23 ),
        .\sr_reg[8]_17 (\sr_reg[8]_24 ),
        .\sr_reg[8]_18 (grn27_n_30),
        .\sr_reg[8]_19 (\sr_reg[8]_37 ),
        .\sr_reg[8]_2 (\sr_reg[8]_8 ),
        .\sr_reg[8]_20 (\sr_reg[8]_38 ),
        .\sr_reg[8]_21 (grn27_n_33),
        .\sr_reg[8]_22 (\sr_reg[8]_43 ),
        .\sr_reg[8]_23 (\sr_reg[8]_56 ),
        .\sr_reg[8]_24 (\sr_reg[8]_57 ),
        .\sr_reg[8]_25 (\sr_reg[8]_58 ),
        .\sr_reg[8]_26 (\sr_reg[8]_60 ),
        .\sr_reg[8]_27 (\sr_reg[8]_62 ),
        .\sr_reg[8]_28 (\sr_reg[8]_63 ),
        .\sr_reg[8]_29 (\sr_reg[8]_64 ),
        .\sr_reg[8]_3 (grn27_n_8),
        .\sr_reg[8]_30 (\sr_reg[8]_26 ),
        .\sr_reg[8]_31 (\sr_reg[8]_66 ),
        .\sr_reg[8]_32 (\sr_reg[8]_68 ),
        .\sr_reg[8]_33 (\sr_reg[8]_69 ),
        .\sr_reg[8]_34 (\sr_reg[8]_70 ),
        .\sr_reg[8]_35 (\sr_reg[8]_75 ),
        .\sr_reg[8]_36 (\sr_reg[8]_82 ),
        .\sr_reg[8]_37 (\sr_reg[8]_40 ),
        .\sr_reg[8]_38 (\sr_reg[8]_94 ),
        .\sr_reg[8]_39 (grn27_n_57),
        .\sr_reg[8]_4 (\sr_reg[8]_10 ),
        .\sr_reg[8]_40 (\sr_reg[8]_101 ),
        .\sr_reg[8]_41 (\sr_reg[8]_104 ),
        .\sr_reg[8]_42 (\sr_reg[8]_106 ),
        .\sr_reg[8]_43 (\sr_reg[8]_108 ),
        .\sr_reg[8]_44 (\sr_reg[8]_109 ),
        .\sr_reg[8]_45 (\sr_reg[8]_85 ),
        .\sr_reg[8]_46 (\sr_reg[8]_120 ),
        .\sr_reg[8]_47 (\sr_reg[8]_128 ),
        .\sr_reg[8]_48 (\sr_reg[8]_129 ),
        .\sr_reg[8]_49 (\sr_reg[8]_130 ),
        .\sr_reg[8]_5 (\sr_reg[8]_9 ),
        .\sr_reg[8]_50 (\sr_reg[8]_42 ),
        .\sr_reg[8]_6 (grn27_n_13),
        .\sr_reg[8]_7 (\sr_reg[8]_11 ),
        .\sr_reg[8]_8 (grn27_n_15),
        .\sr_reg[8]_9 (\sr_reg[8]_12 ),
        .\tr[17]_i_9 (\badr[0]_INST_0_i_1_0 ),
        .\tr[23]_i_10 (\sr_reg[8]_4 ),
        .\tr[25]_i_7 (\sr_reg[8]_50 ),
        .\tr[25]_i_7_0 (\sr_reg[8]_72 ),
        .\tr_reg[1] (\tr_reg[1] ),
        .\tr_reg[1]_0 (\tr_reg[1]_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4F4F4FFF4F)) 
    \iv[0]_i_10 
       (.I0(\iv[0]_i_3 ),
        .I1(\iv[0]_i_21_n_0 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(\iv[0]_i_22_n_0 ),
        .I4(\iv[0]_i_23_n_0 ),
        .I5(\iv[0]_i_3_0 ),
        .O(\sr_reg[8]_15 ));
  LUT6 #(
    .INIT(64'hF505F3F3F5050303)) 
    \iv[0]_i_14 
       (.I0(\sr_reg[8]_47 ),
        .I1(\sr_reg[8]_48 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\iv[0]_i_8 ),
        .I4(\iv[0]_i_10_0 ),
        .I5(\iv[0]_i_8_0 ),
        .O(\sr_reg[8]_67 ));
  LUT6 #(
    .INIT(64'h888AAA8A00022202)) 
    \iv[0]_i_16 
       (.I0(\sr[4]_i_36_0 ),
        .I1(\sr_reg[8]_3 ),
        .I2(\sr_reg[8]_48 ),
        .I3(\iv[0]_i_10_0 ),
        .I4(\sr_reg[8]_47 ),
        .I5(\sr[4]_i_36 ),
        .O(\sr_reg[8]_125 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[0]_i_17 
       (.I0(\sr_reg[8]_47 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_48 ),
        .O(\iv[0]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFF000000FF47FF47)) 
    \iv[0]_i_18 
       (.I0(\sr_reg[8]_47 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_48 ),
        .I3(\iv[13]_i_17_0 ),
        .I4(\niho_dsp_a[16] [2]),
        .I5(\sr_reg[8]_1 ),
        .O(\iv[0]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \iv[0]_i_21 
       (.I0(\iv[0]_i_10_2 ),
        .I1(\sr_reg[8]_48 ),
        .I2(\iv[0]_i_10_0 ),
        .I3(\sr_reg[8]_47 ),
        .I4(\sr_reg[8]_3 ),
        .I5(\iv[0]_i_10_3 ),
        .O(\iv[0]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFFFFF)) 
    \iv[0]_i_22 
       (.I0(\sr_reg[8]_50 ),
        .I1(\iv[0]_i_10_0 ),
        .I2(\iv[0]_i_30_n_0 ),
        .I3(\iv[13]_i_17_0 ),
        .I4(\sr_reg[8]_3 ),
        .O(\iv[0]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hAAAB)) 
    \iv[0]_i_23 
       (.I0(\tr_reg[5] ),
        .I1(\iv[0]_i_10_1 ),
        .I2(\iv[13]_i_17_0 ),
        .I3(\sr_reg[8]_3 ),
        .O(\iv[0]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_28 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr[7]_i_36_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\badr[14]_INST_0_i_1 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr_reg[6]_0 ),
        .O(\sr_reg[8]_92 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_30 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr[7]_i_36_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\badr[14]_INST_0_i_1 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[0]_i_22_0 ),
        .O(\iv[0]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0000B0B0000000FF)) 
    \iv[0]_i_9 
       (.I0(\sr_reg[8]_9 ),
        .I1(\iv[0]_i_17_n_0 ),
        .I2(\iv[0]_i_18_n_0 ),
        .I3(\iv[0]_i_3_1 ),
        .I4(\niho_dsp_a[16] [3]),
        .I5(bbus_0[1]),
        .O(\sr_reg[8]_46 ));
  LUT6 #(
    .INIT(64'hFFFF0000FEAEFEAE)) 
    \iv[10]_i_21 
       (.I0(\iv[0]_i_19 ),
        .I1(\iv[14]_i_48_n_0 ),
        .I2(\sr_reg[8]_93 ),
        .I3(\badr[0]_INST_0_i_1 ),
        .I4(\sr_reg[8]_84 ),
        .I5(\sr[4]_i_89_0 ),
        .O(\sr_reg[8]_17 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[10]_i_22 
       (.I0(\iv[0]_i_19 ),
        .I1(\iv[10]_i_38_n_0 ),
        .I2(\iv[10]_i_39_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\iv[10]_i_10_0 ),
        .O(\sr_reg[8]_41 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_24 
       (.I0(\sr_reg[8]_84 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_99 ),
        .O(\iv[10]_i_24_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[10]_i_27 
       (.I0(\iv[15]_i_149_n_0 ),
        .I1(\iv[15]_i_150_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[10]_i_13 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\badr[15]_INST_0_i_1 ),
        .O(\sr_reg[8]_81 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \iv[10]_i_30 
       (.I0(\iv[0]_i_19 ),
        .I1(\iv[10]_i_38_n_0 ),
        .I2(\iv[10]_i_45_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr[4]_i_64 ),
        .O(\sr_reg[8]_32 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[10]_i_33 
       (.I0(\iv[14]_i_46_n_0 ),
        .I1(\iv[14]_i_47_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_42_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_43_n_0 ),
        .O(\sr_reg[8]_84 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[10]_i_34 
       (.I0(\iv[14]_i_61_n_0 ),
        .I1(\iv[14]_i_62_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_59_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_60_n_0 ),
        .O(\sr_reg[8]_61 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[10]_i_35 
       (.I0(\iv[0]_i_19 ),
        .I1(\iv[10]_i_38_n_0 ),
        .I2(\sr_reg[6]_11 ),
        .O(\iv[10]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_38 
       (.I0(\iv[15]_i_149_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[15]_i_150_n_0 ),
        .O(\iv[10]_i_38_n_0 ));
  LUT3 #(
    .INIT(8'hC5)) 
    \iv[10]_i_39 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(\iv[10]_i_22_0 ),
        .I2(\sr_reg[8]_93 ),
        .O(\iv[10]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[10]_i_42 
       (.I0(\iv[2]_i_24 ),
        .I1(\iv[0]_i_19 ),
        .I2(\sr_reg[6]_0 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\iv[14]_i_48_n_0 ),
        .O(\sr_reg[8]_99 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[10]_i_43 
       (.I0(\sr[7]_i_36_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\badr[14]_INST_0_i_1 ),
        .I3(\iv[0]_i_19 ),
        .I4(\iv[10]_i_25 ),
        .O(\sr_reg[8]_119 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[10]_i_45 
       (.I0(\tr[18]_i_3_2 ),
        .I1(\tr_reg[0] ),
        .I2(\tr[17]_i_3_0 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\badr[15]_INST_0_i_1 ),
        .O(\iv[10]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \iv[10]_i_9 
       (.I0(\sr_reg[8]_17 ),
        .I1(\tr[30]_i_3_4 ),
        .I2(\sr[4]_i_36_0 ),
        .I3(\sr[4]_i_36 ),
        .I4(\sr_reg[8]_40 ),
        .I5(\sr_reg[8]_41 ),
        .O(\sr_reg[8]_39 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_26 
       (.I0(\sr_reg[8]_45 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_44 ),
        .O(\iv[11]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[11]_i_28 
       (.I0(\iv[11]_i_13 ),
        .I1(\badr[16]_INST_0_i_1 ),
        .I2(\iv[0]_i_19 ),
        .I3(\badr[14]_INST_0_i_1_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_63_n_0 ),
        .O(\sr_reg[8]_79 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \iv[11]_i_30 
       (.I0(\iv[0]_i_19 ),
        .I1(\tr[27]_i_6_0 ),
        .I2(\sr_reg[6]_7 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_80 ),
        .O(\iv[11]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[11]_i_31 
       (.I0(\iv[7]_i_43_n_0 ),
        .I1(\iv[0]_i_19 ),
        .I2(\sr_reg[8]_109 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\tr[28]_i_6_0 ),
        .O(\iv[11]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[11]_i_33 
       (.I0(\sr[7]_i_42_n_0 ),
        .I1(\sr[7]_i_43_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr[7]_i_34_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr[7]_i_35_n_0 ),
        .O(\sr_reg[8]_45 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[11]_i_38 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\iv[15]_i_154_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_151_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[15]_i_152_n_0 ),
        .O(\sr_reg[8]_80 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \iv[11]_i_43 
       (.I0(\iv[11]_i_25 ),
        .I1(\iv[0]_i_19 ),
        .I2(\iv[14]_i_45_n_0 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\tr[16]_i_32_n_0 ),
        .O(\sr_reg[8]_114 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \iv[11]_i_44 
       (.I0(\badr[0]_INST_0_i_1_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\sr[7]_i_41_n_0 ),
        .I3(\iv[0]_i_19 ),
        .I4(\iv[3]_i_31 ),
        .O(\sr_reg[8]_44 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[12]_i_25 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr_reg[8]_115 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\sr_reg[8]_116 ),
        .I4(\sr[4]_i_98_0 ),
        .O(\iv[12]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[12]_i_27 
       (.I0(\iv[12]_i_13 ),
        .I1(\iv[0]_i_19 ),
        .I2(\badr[15]_INST_0_i_1 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\iv[15]_i_149_n_0 ),
        .O(\sr_reg[8]_74 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_29 
       (.I0(\sr_reg[8]_110 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_59 ),
        .O(\iv[12]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_30 
       (.I0(\sr_reg[8]_74 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\tr[29]_i_8_0 ),
        .O(\iv[12]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[12]_i_33 
       (.I0(\iv[14]_i_43_n_0 ),
        .I1(\iv[14]_i_44_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_47_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_42_n_0 ),
        .O(\sr_reg[8]_115 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[12]_i_34 
       (.I0(\iv[14]_i_64_n_0 ),
        .I1(\iv[14]_i_61_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_62_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_59_n_0 ),
        .O(\sr_reg[8]_59 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_35 
       (.I0(\iv[12]_i_50_n_0 ),
        .I1(\iv[0]_i_19 ),
        .I2(\sr_reg[8]_94 ),
        .O(\iv[12]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[12]_i_49 
       (.I0(\iv[14]_i_60_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\sr_reg[6]_3 ),
        .I3(\iv[0]_i_19 ),
        .I4(\iv[4]_i_31 ),
        .O(\sr_reg[8]_110 ));
  LUT5 #(
    .INIT(32'hF044F077)) 
    \iv[12]_i_50 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\iv[14]_i_60_n_0 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\niho_dsp_a[16] [2]),
        .O(\iv[12]_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[13]_i_23 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr_reg[8]_76 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\sr_reg[8]_96 ),
        .I4(\sr_reg[8]_106 ),
        .O(\sr_reg[8]_13 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[13]_i_25 
       (.I0(\sr_reg[8]_76 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[6]_1 ),
        .I3(\iv[0]_i_19 ),
        .I4(\sr_reg[8]_96 ),
        .O(\iv[13]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \iv[13]_i_29 
       (.I0(\badr[16]_INST_0_i_1 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\badr[14]_INST_0_i_1_0 ),
        .I3(\iv[0]_i_19 ),
        .I4(\iv[13]_i_13 ),
        .O(\sr_reg[8]_78 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_31 
       (.I0(\sr_reg[8]_78 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\tr[30]_i_9_0 ),
        .O(\iv[13]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_32 
       (.I0(\sr_reg[8]_95 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\iv[13]_i_36_n_0 ),
        .O(\iv[13]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[13]_i_35 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr[7]_i_36_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr[7]_i_43_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr[7]_i_34_n_0 ),
        .O(\sr_reg[8]_76 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[13]_i_36 
       (.I0(\iv[15]_i_150_n_0 ),
        .I1(\iv[15]_i_151_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_152_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[15]_i_153_n_0 ),
        .O(\iv[13]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[13]_i_37 
       (.I0(\iv[15]_i_154_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[15]_i_155_n_0 ),
        .I3(\iv[0]_i_19 ),
        .I4(\sr_reg[6]_9 ),
        .O(\iv[13]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h5500C3FF55FFC3FF)) 
    \iv[13]_i_39 
       (.I0(\tr_reg[5] ),
        .I1(DI[1]),
        .I2(bbus_0[3]),
        .I3(\iv[13]_i_17 ),
        .I4(\iv[13]_i_17_0 ),
        .I5(\iv[13]_i_17_1 ),
        .O(\badr[21]_INST_0_i_1 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[13]_i_41 
       (.I0(\sr[4]_i_36 ),
        .I1(\tr_reg[0] ),
        .I2(\niho_dsp_a[16] [2]),
        .I3(\sr_reg[8]_93 ),
        .I4(\badr[0]_INST_0_i_1_0 ),
        .O(\sr_reg[6]_1 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[13]_i_44 
       (.I0(\tr[16]_i_32_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[13]_i_26 ),
        .I3(\iv[0]_i_19 ),
        .I4(\iv[13]_i_26_0 ),
        .O(\sr_reg[8]_105 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[13]_i_46 
       (.I0(DI[1]),
        .I1(\tr_reg[0] ),
        .I2(DI[2]),
        .O(\badr[14]_INST_0_i_1_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[13]_i_50 
       (.I0(\iv[15]_i_154_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[15]_i_155_n_0 ),
        .I3(\iv[0]_i_19 ),
        .I4(\iv[5]_i_30 ),
        .O(\sr_reg[8]_95 ));
  LUT4 #(
    .INIT(16'h60CC)) 
    \iv[14]_i_15 
       (.I0(\tr_reg[5] ),
        .I1(bbus_0[1]),
        .I2(\niho_dsp_a[16] [3]),
        .I3(\sr[6]_i_12_2 ),
        .O(\sr_reg[8]_3 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_16 
       (.I0(\sr_reg[8]_73 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[6]_4 ),
        .O(\iv[14]_i_35_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[14]_i_24 
       (.I0(\iv[14]_i_42_n_0 ),
        .I1(\iv[14]_i_43_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_44_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_45_n_0 ),
        .O(\sr_reg[8]_73 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[14]_i_32 
       (.I0(\sr_reg[8]_100 ),
        .I1(\iv[0]_i_19 ),
        .I2(\iv[14]_i_57_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_77 ),
        .O(\sr_reg[8]_27 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[14]_i_35 
       (.I0(\sr_reg[6]_0 ),
        .I1(\iv[14]_i_48_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_46_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_47_n_0 ),
        .O(\sr_reg[6]_4 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_38 
       (.I0(\iv[14]_i_59_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[14]_i_60_n_0 ),
        .O(\sr_reg[8]_100 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[14]_i_39 
       (.I0(\iv[14]_i_61_n_0 ),
        .I1(\iv[14]_i_62_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_63_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_64_n_0 ),
        .O(\sr_reg[8]_77 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_42 
       (.I0(\abus_o[11] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [3]),
        .O(\iv[14]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_43 
       (.I0(\abus_o[11] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [1]),
        .O(\iv[14]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_44 
       (.I0(DI[0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [3]),
        .O(\iv[14]_i_44_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[14]_i_45 
       (.I0(DI[1]),
        .I1(\tr_reg[0] ),
        .I2(DI[2]),
        .O(\iv[14]_i_45_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_46 
       (.I0(\abus_o[7] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [3]),
        .O(\iv[14]_i_46_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[14]_i_47 
       (.I0(\abus_o[7] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [2]),
        .O(\iv[14]_i_47_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_48 
       (.I0(\abus_o[3] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [1]),
        .O(\iv[14]_i_48_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_54 
       (.I0(DI[2]),
        .I1(\tr_reg[0] ),
        .I2(DI[3]),
        .O(\badr[15]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h470047CC473347FF)) 
    \iv[14]_i_57 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\niho_dsp_a[16] [2]),
        .I3(\sr_reg[8]_93 ),
        .I4(\sr[4]_i_36 ),
        .I5(\iv[14]_i_32_0 ),
        .O(\iv[14]_i_57_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \iv[14]_i_58 
       (.I0(\abus_o[3] [0]),
        .I1(\niho_dsp_a[16] [2]),
        .I2(\tr_reg[0] ),
        .O(\sr_reg[6]_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_59 
       (.I0(\abus_o[3] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [0]),
        .O(\iv[14]_i_59_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_60 
       (.I0(\abus_o[3] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [2]),
        .O(\iv[14]_i_60_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_61 
       (.I0(\abus_o[7] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [0]),
        .O(\iv[14]_i_61_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_62 
       (.I0(\abus_o[7] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [2]),
        .O(\iv[14]_i_62_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_63 
       (.I0(\abus_o[11] [3]),
        .I1(\tr_reg[0] ),
        .I2(DI[0]),
        .O(\iv[14]_i_63_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[14]_i_64 
       (.I0(\abus_o[11] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [2]),
        .O(\iv[14]_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_103 
       (.I0(\iv[15]_i_149_n_0 ),
        .I1(\iv[15]_i_150_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_151_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[15]_i_152_n_0 ),
        .O(\sr_reg[8]_52 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_104 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\iv[15]_i_154_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_155_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[15]_i_60_0 ),
        .O(\iv[15]_i_104_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_106 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\iv[15]_i_154_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_155_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[15]_i_157_n_0 ),
        .O(\iv[15]_i_106_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_110 
       (.I0(\abus_o[7] [3]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_6 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_148 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(\tr[17]_i_3_0 ),
        .O(\badr[16]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_149 
       (.I0(DI[0]),
        .I1(\tr_reg[0] ),
        .I2(DI[1]),
        .O(\iv[15]_i_149_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_150 
       (.I0(\abus_o[11] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [3]),
        .O(\iv[15]_i_150_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_151 
       (.I0(\abus_o[11] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [1]),
        .O(\iv[15]_i_151_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_152 
       (.I0(\abus_o[7] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [3]),
        .O(\iv[15]_i_152_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_153 
       (.I0(\abus_o[7] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [1]),
        .O(\iv[15]_i_153_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_154 
       (.I0(\abus_o[3] [2]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [3]),
        .O(\iv[15]_i_154_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \iv[15]_i_155 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [1]),
        .O(\iv[15]_i_155_n_0 ));
  LUT3 #(
    .INIT(8'h35)) 
    \iv[15]_i_157 
       (.I0(DI[3]),
        .I1(\niho_dsp_a[16] [2]),
        .I2(\tr_reg[0] ),
        .O(\iv[15]_i_157_n_0 ));
  LUT6 #(
    .INIT(64'h4F4F4F4F4F4F4F44)) 
    \iv[15]_i_22 
       (.I0(\iv[15]_i_55_n_0 ),
        .I1(\iv[15]_i_8 ),
        .I2(\iv[15]_i_8_0 ),
        .I3(\iv[15]_i_8_1 ),
        .I4(\iv[15]_i_8_2 ),
        .I5(\iv[15]_i_60_n_0 ),
        .O(\sr_reg[8]_34 ));
  LUT5 #(
    .INIT(32'h0000202A)) 
    \iv[15]_i_53 
       (.I0(\sr_reg[8]_35 ),
        .I1(\sr_reg[8]_65 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\sr_reg[8]_4 ),
        .I4(\sr_reg[8]_1 ),
        .O(\sr_reg[8]_88 ));
  LUT6 #(
    .INIT(64'hFF00B8B8FFFFB8B8)) 
    \iv[15]_i_55 
       (.I0(\sr_reg[8]_65 ),
        .I1(\iv[0]_i_10_0 ),
        .I2(\sr_reg[8]_4 ),
        .I3(\iv[15]_i_22_0 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\iv[13]_i_17_0 ),
        .O(\iv[15]_i_55_n_0 ));
  LUT5 #(
    .INIT(32'h00088808)) 
    \iv[15]_i_60 
       (.I0(\iv[13]_i_17_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\sr_reg[8]_52 ),
        .I3(\iv[0]_i_10_0 ),
        .I4(\iv[15]_i_104_n_0 ),
        .O(\iv[15]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'h0000000D0D0D000D)) 
    \iv[15]_i_61 
       (.I0(\sr_reg[8]_1 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(bbus_0[1]),
        .I3(\sr_reg[8]_4 ),
        .I4(\iv[0]_i_10_0 ),
        .I5(\sr_reg[8]_65 ),
        .O(\sr_reg[8]_87 ));
  LUT5 #(
    .INIT(32'h00B80000)) 
    \iv[15]_i_64 
       (.I0(\iv[15]_i_106_n_0 ),
        .I1(\iv[0]_i_10_0 ),
        .I2(\sr_reg[8]_52 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\iv[13]_i_17_0 ),
        .O(\sr_reg[8]_51 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[1]_i_18 
       (.I0(\sr[4]_i_85_0 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\sr_reg[8]_61 ),
        .I4(\iv[0]_i_10_0 ),
        .I5(\sr_reg[8]_83 ),
        .O(\iv[1]_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[1]_i_25 
       (.I0(\sr_reg[8]_97 ),
        .I1(\iv[0]_i_19 ),
        .I2(\sr_reg[8]_103 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_84 ),
        .O(\iv[1]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[1]_i_29 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr_reg[8]_61 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\sr_reg[8]_108 ),
        .I4(\iv[9]_i_51_n_0 ),
        .O(\sr_reg[8]_30 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[2]_i_17 
       (.I0(\sr[4]_i_108_0 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\sr_reg[8]_80 ),
        .I4(\iv[0]_i_10_0 ),
        .I5(\sr_reg[8]_81 ),
        .O(\iv[2]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[2]_i_26 
       (.I0(\sr_reg[8]_119 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_45 ),
        .O(\iv[2]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[2]_i_29 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr_reg[8]_80 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\iv[10]_i_38_n_0 ),
        .I4(\iv[10]_i_45_n_0 ),
        .O(\sr_reg[8]_33 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[2]_i_31 
       (.I0(\iv[13]_i_17_0 ),
        .I1(\abus_o[3] [1]),
        .I2(\niho_dsp_a[16] [3]),
        .I3(\sr_reg[8]_1 ),
        .O(\iv[2]_i_31_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[3]_i_18 
       (.I0(\sr[4]_i_104_0 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\sr_reg[8]_59 ),
        .I4(\iv[0]_i_10_0 ),
        .I5(\sr_reg[8]_79 ),
        .O(\iv[3]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[3]_i_30 
       (.I0(\sr_reg[8]_114 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_115 ),
        .O(\iv[3]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_34 
       (.I0(\sr_reg[8]_59 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\iv[7]_i_43_n_0 ),
        .I3(\iv[0]_i_19 ),
        .I4(\sr_reg[8]_109 ),
        .O(\sr_reg[8]_28 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[4]_i_18 
       (.I0(\sr[4]_i_53_0 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\iv[13]_i_36_n_0 ),
        .I4(\iv[0]_i_10_0 ),
        .I5(\sr_reg[8]_74 ),
        .O(\iv[4]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_23 
       (.I0(\iv[14]_i_48_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[14]_i_46_n_0 ),
        .O(\sr_reg[8]_116 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[4]_i_24 
       (.I0(\tr_reg[0] ),
        .I1(\abus_o[3] [0]),
        .O(\badr[0]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_32 
       (.I0(\iv[13]_i_36_n_0 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_74 ),
        .O(\iv[12]_i_27_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[4]_i_34 
       (.I0(\iv[13]_i_17_0 ),
        .I1(\abus_o[3] [3]),
        .I2(\niho_dsp_a[16] [3]),
        .I3(\sr_reg[8]_1 ),
        .O(\iv[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[5]_i_18 
       (.I0(\sr[4]_i_58_0 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\sr_reg[8]_77 ),
        .I4(\iv[0]_i_10_0 ),
        .I5(\sr_reg[8]_78 ),
        .O(\iv[5]_i_18_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_24 
       (.I0(\sr[7]_i_41_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\sr[7]_i_42_n_0 ),
        .O(\sr_reg[8]_96 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_28 
       (.I0(\sr_reg[8]_105 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_73 ),
        .O(\iv[5]_i_28_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_31 
       (.I0(\sr_reg[8]_77 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_78 ),
        .O(\iv[13]_i_29_0 ));
  LUT4 #(
    .INIT(16'hF7F0)) 
    \iv[5]_i_33 
       (.I0(\iv[13]_i_17_0 ),
        .I1(\abus_o[7] [0]),
        .I2(\niho_dsp_a[16] [3]),
        .I3(\sr_reg[8]_1 ),
        .O(\iv[5]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[6]_i_29 
       (.I0(\tr[22]_i_8_0 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_100 ),
        .I3(\iv[0]_i_19 ),
        .I4(\iv[14]_i_57_n_0 ),
        .O(\iv[6]_i_29_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[6]_i_30 
       (.I0(\sr_reg[8]_52 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\tr[23]_i_6_0 ),
        .O(\iv[6]_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[7]_i_37 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr[4]_i_89_1 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\iv[7]_i_46_n_0 ),
        .I4(\sr_reg[8]_113 ),
        .O(\iv[7]_i_37_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_38 
       (.I0(\sr_reg[8]_4 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\tr[23]_i_7_0 ),
        .O(\iv[7]_i_38_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[7]_i_41 
       (.I0(\badr[14]_INST_0_i_1_0 ),
        .I1(\iv[14]_i_63_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_64_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_61_n_0 ),
        .O(\sr_reg[8]_55 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \iv[7]_i_43 
       (.I0(\tr[18]_i_3_2 ),
        .I1(\tr_reg[0] ),
        .I2(\tr[19]_i_3_3 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\badr[16]_INST_0_i_1 ),
        .O(\iv[7]_i_43_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_44 
       (.I0(\iv[14]_i_43_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[14]_i_44_n_0 ),
        .O(\sr_reg[8]_113 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_45 
       (.I0(\iv[15]_i_153_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[15]_i_154_n_0 ),
        .O(\sr_reg[8]_118 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_46 
       (.I0(\iv[14]_i_45_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\tr[16]_i_32_n_0 ),
        .O(\iv[7]_i_46_n_0 ));
  LUT5 #(
    .INIT(32'h00FF4747)) 
    \iv[8]_i_26 
       (.I0(\sr_reg[8]_91 ),
        .I1(\iv[0]_i_19 ),
        .I2(\iv[8]_i_41_n_0 ),
        .I3(\sr[4]_i_76_0 ),
        .I4(\sr[4]_i_89_0 ),
        .O(\iv[8]_i_26_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_27 
       (.I0(\sr_reg[8]_49 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\tr[24]_i_10_1 ),
        .O(\iv[8]_i_27_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[8]_i_29 
       (.I0(\badr[15]_INST_0_i_1 ),
        .I1(\iv[15]_i_149_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_150_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[15]_i_151_n_0 ),
        .O(\sr_reg[8]_48 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_32 
       (.I0(\sr_reg[8]_48 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr[4]_i_75 ),
        .O(\iv[8]_i_30 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[8]_i_35 
       (.I0(\iv[14]_i_48_n_0 ),
        .I1(\iv[14]_i_46_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_47_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_42_n_0 ),
        .O(\sr_reg[8]_49 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_36 
       (.I0(\sr[7]_i_35_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\sr[7]_i_36_n_0 ),
        .O(\sr_reg[8]_91 ));
  LUT5 #(
    .INIT(32'h88B8B8B8)) 
    \iv[8]_i_37 
       (.I0(\badr[14]_INST_0_i_1 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\badr[0]_INST_0_i_1 ),
        .I3(\niho_dsp_a[16] [2]),
        .I4(\tr_reg[0] ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[8]_i_38 
       (.I0(\iv[14]_i_62_n_0 ),
        .I1(\iv[14]_i_59_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_60_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr_reg[6]_3 ),
        .O(\sr_reg[8]_112 ));
  LUT5 #(
    .INIT(32'h888BBB8B)) 
    \iv[8]_i_41 
       (.I0(\badr[14]_INST_0_i_1 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\tr[18]_i_3_2 ),
        .I3(\tr_reg[0] ),
        .I4(\tr[17]_i_3_0 ),
        .O(\iv[8]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[8]_i_42 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\niho_dsp_a[16] [2]),
        .O(\sr_reg[6]_3 ));
  LUT4 #(
    .INIT(16'h60CC)) 
    \iv[9]_i_16 
       (.I0(\tr_reg[5] ),
        .I1(bbus_0[1]),
        .I2(\niho_dsp_a[16] [3]),
        .I3(\sr[6]_i_12_2 ),
        .O(\sr_reg[8]_1 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_28 
       (.I0(\sr_reg[8]_50 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\tr[25]_i_10_0 ),
        .O(\iv[9]_i_28_n_0 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[9]_i_30 
       (.I0(\iv[14]_i_63_n_0 ),
        .I1(\iv[14]_i_64_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\badr[16]_INST_0_i_1 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\badr[14]_INST_0_i_1_0 ),
        .O(\sr_reg[8]_83 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \iv[9]_i_33 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr_reg[8]_108 ),
        .I2(\iv[9]_i_51_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr[4]_i_67 ),
        .O(\sr_reg[8]_29 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_35 
       (.I0(\sr[7]_i_41_n_0 ),
        .I1(\sr[7]_i_42_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr[7]_i_43_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr[7]_i_34_n_0 ),
        .O(\sr_reg[8]_50 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[9]_i_36 
       (.I0(\iv[0]_i_19 ),
        .I1(\badr[0]_INST_0_i_1_0 ),
        .I2(\sr_reg[8]_93 ),
        .O(\sr_reg[8]_72 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_37 
       (.I0(\iv[14]_i_44_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[14]_i_45_n_0 ),
        .O(\sr_reg[8]_97 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[9]_i_38 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(\niho_dsp_a[16] [2]),
        .I3(\sr_reg[8]_93 ),
        .I4(\badr[0]_INST_0_i_1_0 ),
        .O(\sr_reg[6]_2 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_41 
       (.I0(\iv[15]_i_152_n_0 ),
        .I1(\iv[15]_i_153_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_154_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[15]_i_155_n_0 ),
        .O(\sr_reg[8]_47 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[9]_i_43 
       (.I0(\abus_o[3] [1]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_8 ));
  LUT5 #(
    .INIT(32'h888BBB8B)) 
    \iv[9]_i_48 
       (.I0(\tr[16]_i_32_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\tr[19]_i_3_3 ),
        .I3(\tr_reg[0] ),
        .I4(\tr[18]_i_3_2 ),
        .O(\sr_reg[8]_103 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_51 
       (.I0(\badr[16]_INST_0_i_1 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\badr[14]_INST_0_i_1_0 ),
        .O(\iv[9]_i_51_n_0 ));
  CARRY4 \iv_reg[3]_i_11 
       (.CI(\<const0> ),
        .CO({\iv_reg[3]_i_11_n_0 ,\iv_reg[3]_i_11_n_1 ,\iv_reg[3]_i_11_n_2 ,\iv_reg[3]_i_11_n_3 }),
        .CYINIT(\iv[0]_i_6 ),
        .DI(\abus_o[3] ),
        .O(\sr_reg[6]_8 ),
        .S({\iv[0]_i_6_0 ,\art/add/iv[3]_i_26_n_0 }));
  CARRY4 \iv_reg[7]_i_12 
       (.CI(\iv_reg[3]_i_11_n_0 ),
        .CO({\iv_reg[7]_i_12_n_0 ,\iv_reg[7]_i_12_n_1 ,\iv_reg[7]_i_12_n_2 ,\iv_reg[7]_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\abus_o[7] ),
        .O(\art/add/iv[7]_i_32 ),
        .S({\iv[4]_i_6 [2:1],\art/add/iv[7]_i_31_n_0 ,\iv[4]_i_6 [0]}));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[16]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[0]),
        .O(niho_dsp_a[0]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[17]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[1]),
        .O(niho_dsp_a[1]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[18]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[2]),
        .O(niho_dsp_a[2]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[19]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[3]),
        .O(niho_dsp_a[3]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[20]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[4]),
        .O(niho_dsp_a[4]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[21]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[5]),
        .O(niho_dsp_a[5]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[22]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[6]),
        .O(niho_dsp_a[6]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[23]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[7]),
        .O(niho_dsp_a[7]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[24]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[8]),
        .O(niho_dsp_a[8]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[25]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[9]),
        .O(niho_dsp_a[9]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[26]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[10]),
        .O(niho_dsp_a[10]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[27]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[11]),
        .O(niho_dsp_a[11]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[28]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[12]),
        .O(niho_dsp_a[12]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[29]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[13]),
        .O(niho_dsp_a[13]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[30]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[14]),
        .O(niho_dsp_a[14]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[31]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[15]),
        .O(niho_dsp_a[15]));
  LUT5 #(
    .INIT(32'hF8888888)) 
    \niho_dsp_a[32]_INST_0 
       (.I0(\niho_dsp_a[16]_0 ),
        .I1(\sr_reg[8]_120 ),
        .I2(\niho_dsp_a[16] [3]),
        .I3(mul_rslt),
        .I4(mul_a[16]),
        .O(niho_dsp_a[16]));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_101 
       (.I0(\iv[15]_i_8 ),
        .I1(\sr[4]_i_45_1 ),
        .I2(\iv[13]_i_32_n_0 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\iv[13]_i_31_n_0 ),
        .I5(\tr[16]_i_6_2 ),
        .O(\sr[4]_i_101_n_0 ));
  LUT6 #(
    .INIT(64'h530053005300530F)) 
    \sr[4]_i_102 
       (.I0(\tr[30]_i_3_0 ),
        .I1(\iv[13]_i_25_n_0 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\iv[13]_i_17_0 ),
        .I4(\sr_reg[8]_13 ),
        .I5(\tr_reg[5] ),
        .O(\sr[4]_i_102_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_104 
       (.I0(\iv[3]_i_18_n_0 ),
        .I1(bbus_0[1]),
        .O(\sr[4]_i_104_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_106 
       (.I0(\tr_reg[5] ),
        .I1(\iv[3]_i_18_n_0 ),
        .O(\sr[4]_i_106_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F000F0D0F08)) 
    \sr[4]_i_107 
       (.I0(\iv[0]_i_10_0 ),
        .I1(\sr_reg[8]_80 ),
        .I2(\sr[4]_i_45_2 ),
        .I3(\iv[2]_i_31_n_0 ),
        .I4(\iv[10]_i_35_n_0 ),
        .I5(\sr_reg[8]_9 ),
        .O(\sr[4]_i_107_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_108 
       (.I0(\iv[2]_i_17_n_0 ),
        .I1(bbus_0[1]),
        .O(\sr[4]_i_108_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_110 
       (.I0(\tr_reg[5] ),
        .I1(\iv[2]_i_17_n_0 ),
        .O(\sr[4]_i_110_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_113 
       (.I0(\sr_reg[6]_8 [2]),
        .I1(\art/add/sr[5]_i_18 [0]),
        .I2(\art/add/iv[7]_i_32 [0]),
        .I3(\art/add/sr[5]_i_18 [1]),
        .O(\sr[4]_i_113_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[4]_i_114 
       (.I0(\sr_reg[8]_84 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(grn27_n_57),
        .I3(\iv[0]_i_19 ),
        .I4(grn27_n_58),
        .O(\sr[4]_i_114_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \sr[4]_i_116 
       (.I0(\sr_reg[8]_1 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_72 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_50 ),
        .O(\sr_reg[8]_25 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \sr[4]_i_118 
       (.I0(\sr_reg[8]_1 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\tr[25]_i_10_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_50 ),
        .O(\sr[4]_i_118_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_12 
       (.I0(\tr[23]_i_3_n_0 ),
        .I1(\tr[17]_i_9_0 ),
        .I2(\tr[24]_i_10_0 ),
        .I3(\tr[30]_i_10_0 ),
        .O(\sr[4]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[4]_i_122 
       (.I0(\sr_reg[6]_4 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_65 ),
        .O(\sr[4]_i_122_n_0 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \sr[4]_i_127 
       (.I0(\sr_reg[8]_1 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\tr[24]_i_10_1 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_49 ),
        .O(\sr[4]_i_127_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \sr[4]_i_13 
       (.I0(\tr[20]_i_9_0 ),
        .I1(\tr[21]_i_3_n_0 ),
        .I2(\tr[22]_i_9_0 ),
        .O(\sr[4]_i_13_n_0 ));
  LUT5 #(
    .INIT(32'hFFFEEEFE)) 
    \sr[4]_i_132 
       (.I0(\sr_reg[8]_3 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr[4]_i_159_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_73 ),
        .O(\sr_reg[8]_22 ));
  LUT3 #(
    .INIT(8'h08)) 
    \sr[4]_i_134 
       (.I0(\iv[13]_i_17_0 ),
        .I1(\sr_reg[8]_3 ),
        .I2(\sr[4]_i_80_0 ),
        .O(\sr[4]_i_134_n_0 ));
  LUT6 #(
    .INIT(64'h0050F0500050F350)) 
    \sr[4]_i_138 
       (.I0(\sr[4]_i_162_n_0 ),
        .I1(\sr_reg[8]_3 ),
        .I2(\iv[13]_i_17_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_4 ),
        .I5(bbus_0[1]),
        .O(\sr_reg[8]_86 ));
  LUT4 #(
    .INIT(16'h0004)) 
    \sr[4]_i_14 
       (.I0(\sr_reg[8]_31 ),
        .I1(\tr[19]_i_3_n_0 ),
        .I2(\tr[27]_i_3_n_0 ),
        .I3(\tr[28]_i_3_n_0 ),
        .O(\sr[4]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFF47FFFF)) 
    \sr[4]_i_140 
       (.I0(\sr_reg[8]_55 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\iv[15]_i_106_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\iv[13]_i_17_0 ),
        .O(\sr_reg[8]_54 ));
  LUT6 #(
    .INIT(64'h0010301000103310)) 
    \sr[4]_i_142 
       (.I0(\tr[23]_i_7_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\iv[13]_i_17_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_4 ),
        .I5(\tr_reg[5] ),
        .O(\sr[4]_i_142_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFEEEEEFFFE)) 
    \sr[4]_i_147 
       (.I0(\sr_reg[8]_3 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_85 ),
        .I3(\iv[0]_i_19 ),
        .I4(\sr[4]_i_89_0 ),
        .I5(\sr_reg[8]_45 ),
        .O(\sr_reg[8]_6 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \sr[4]_i_149 
       (.I0(\sr_reg[8]_1 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_44 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_45 ),
        .O(\sr[4]_i_149_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_15 
       (.I0(\tr[18]_i_9_0 ),
        .I1(\sr[4]_i_4_0 ),
        .I2(\tr[26]_i_9_0 ),
        .I3(\tr[29]_i_3_n_0 ),
        .O(\sr[4]_i_15_n_0 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \sr[4]_i_153 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr_reg[8]_115 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\sr_reg[8]_116 ),
        .I4(\sr_reg[6] ),
        .O(\sr_reg[8]_132 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \sr[4]_i_154 
       (.I0(\iv[0]_i_19 ),
        .I1(\sr_reg[8]_76 ),
        .I2(\sr[4]_i_89_0 ),
        .I3(\sr_reg[8]_96 ),
        .I4(\sr_reg[6]_2 ),
        .O(\sr_reg[8]_131 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \sr[4]_i_156 
       (.I0(\iv[14]_i_63_n_0 ),
        .I1(\iv[14]_i_64_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[15]_i_157_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\badr[14]_INST_0_i_1_0 ),
        .O(\sr_reg[8]_102 ));
  LUT6 #(
    .INIT(64'hF5050303F505F3F3)) 
    \sr[4]_i_158 
       (.I0(\iv[14]_i_63_n_0 ),
        .I1(\iv[14]_i_64_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr[4]_i_152 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\badr[14]_INST_0_i_1_0 ),
        .O(\sr_reg[8]_107 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \sr[4]_i_159 
       (.I0(\iv[14]_i_46_n_0 ),
        .I1(\iv[14]_i_47_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\badr[0]_INST_0_i_1 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_48_n_0 ),
        .O(\sr[4]_i_159_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDCFC00000000)) 
    \sr[4]_i_16 
       (.I0(\sr[4]_i_31_n_0 ),
        .I1(\sr[4]_i_32_n_0 ),
        .I2(\tr_reg[1]_0 ),
        .I3(\sr[4]_i_33_n_0 ),
        .I4(\sr[4]_i_34_n_0 ),
        .I5(\tr_reg[1] ),
        .O(\sr[4]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_160 
       (.I0(\iv[14]_i_59_n_0 ),
        .I1(\iv[14]_i_60_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr_reg[6]_3 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\badr[15]_INST_0_i_1 ),
        .O(\sr_reg[8]_98 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_162 
       (.I0(\iv[14]_i_43_n_0 ),
        .I1(\iv[14]_i_44_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_45_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr[4]_i_168_n_0 ),
        .O(\sr[4]_i_162_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_165 
       (.I0(\iv[15]_i_155_n_0 ),
        .I1(\iv[15]_i_157_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\badr[14]_INST_0_i_1_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_63_n_0 ),
        .O(\sr_reg[6]_5 ));
  LUT6 #(
    .INIT(64'hF505F3F3F5050303)) 
    \sr[4]_i_167 
       (.I0(\badr[14]_INST_0_i_1_0 ),
        .I1(\iv[14]_i_63_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr[4]_i_152_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr[4]_i_152 ),
        .O(\sr_reg[8]_111 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[4]_i_168 
       (.I0(\niho_dsp_a[16] [2]),
        .I1(\tr_reg[0] ),
        .I2(DI[3]),
        .O(\sr[4]_i_168_n_0 ));
  LUT6 #(
    .INIT(64'hFBF0FFF0FFF0FFF0)) 
    \sr[4]_i_19 
       (.I0(grn27_n_7),
        .I1(\sr[4]_i_41_n_0 ),
        .I2(\sr[4]_i_5_0 ),
        .I3(\tr_reg[1] ),
        .I4(\sr[4]_i_5_1 ),
        .I5(\sr[4]_i_5_2 ),
        .O(\sr[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDCFC00000000)) 
    \sr[4]_i_20 
       (.I0(\sr[4]_i_44_n_0 ),
        .I1(\sr[4]_i_5_4 ),
        .I2(\tr_reg[1]_0 ),
        .I3(\sr[4]_i_45_n_0 ),
        .I4(\sr[4]_i_5_5 ),
        .I5(\tr_reg[1] ),
        .O(\sr[4]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFDCFC00000000)) 
    \sr[4]_i_21 
       (.I0(\sr[4]_i_46_n_0 ),
        .I1(\sr[4]_i_5_3 ),
        .I2(\tr_reg[1]_0 ),
        .I3(\sr[4]_i_47_n_0 ),
        .I4(grn27_n_10),
        .I5(\tr_reg[1] ),
        .O(\sr[4]_i_21_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_29 
       (.I0(\sr[4]_i_50_n_0 ),
        .I1(\art/add/iv[7]_i_32 [1]),
        .I2(\art/add/sr[5]_i_14 [3]),
        .I3(\sr_reg[6]_8 [0]),
        .I4(\art/add/sr[5]_i_14 [0]),
        .I5(\sr[4]_i_51_n_0 ),
        .O(\sr[4]_i_51_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_31 
       (.I0(\sr[4]_i_52_n_0 ),
        .I1(\sr[4]_i_53_n_0 ),
        .I2(grn27_n_44),
        .I3(\sr[4]_i_16_2 ),
        .I4(\sr[4]_i_55_n_0 ),
        .I5(grn27_n_22),
        .O(\sr[4]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_32 
       (.I0(\sr[4]_i_16_3 ),
        .I1(\sr[4]_i_56_n_0 ),
        .I2(\sr[4]_i_16_5 ),
        .O(\sr[4]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_33 
       (.I0(\sr[4]_i_57_n_0 ),
        .I1(\sr[4]_i_58_n_0 ),
        .I2(\sr[4]_i_16_0 ),
        .I3(\sr[4]_i_16_1 ),
        .I4(\sr[4]_i_60_n_0 ),
        .I5(grn27_n_20),
        .O(\sr[4]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \sr[4]_i_34 
       (.I0(\sr[4]_i_16_3 ),
        .I1(\sr[4]_i_61_n_0 ),
        .I2(\sr[4]_i_16_4 ),
        .O(\sr[4]_i_34_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0EEE0EEEE)) 
    \sr[4]_i_35 
       (.I0(\sr[4]_i_62_n_0 ),
        .I1(\sr[4]_i_63_n_0 ),
        .I2(\sr[4]_i_17 ),
        .I3(\sr[4]_i_17_0 ),
        .I4(\tr_reg[5] ),
        .I5(\sr[4]_i_65_n_0 ),
        .O(\sr[4]_i_65_0 ));
  LUT6 #(
    .INIT(64'hF1F1F100FFFFFFFF)) 
    \sr[4]_i_38 
       (.I0(\sr[4]_i_18 ),
        .I1(\sr[4]_i_70_n_0 ),
        .I2(\sr[4]_i_71_n_0 ),
        .I3(\sr[4]_i_72_n_0 ),
        .I4(\sr[4]_i_18_0 ),
        .I5(\tr_reg[1]_0 ),
        .O(\sr_reg[8]_122 ));
  LUT6 #(
    .INIT(64'h00000100FFFFFFFF)) 
    \sr[4]_i_4 
       (.I0(\sr_reg[8] ),
        .I1(\sr[4]_i_12_n_0 ),
        .I2(\sr[4]_i_13_n_0 ),
        .I3(\sr[4]_i_14_n_0 ),
        .I4(\sr[4]_i_15_n_0 ),
        .I5(\niho_dsp_a[16] [3]),
        .O(\sr_reg[8]_121 ));
  LUT6 #(
    .INIT(64'hF1F1F100FFFFFFFF)) 
    \sr[4]_i_41 
       (.I0(\sr[4]_i_82_n_0 ),
        .I1(\sr[4]_i_83_n_0 ),
        .I2(\sr[4]_i_19_1 ),
        .I3(\sr[4]_i_85_n_0 ),
        .I4(\sr[4]_i_19_2 ),
        .I5(\tr_reg[1]_0 ),
        .O(\sr[4]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0EEE0EEEE)) 
    \sr[4]_i_44 
       (.I0(\sr[4]_i_95_n_0 ),
        .I1(\sr[4]_i_20_2 ),
        .I2(\sr[4]_i_97_n_0 ),
        .I3(\sr[4]_i_20_3 ),
        .I4(\tr_reg[5] ),
        .I5(\sr[4]_i_98_n_0 ),
        .O(\sr[4]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'hE0E0E0E0EEE0EEEE)) 
    \sr[4]_i_45 
       (.I0(\sr[4]_i_99_n_0 ),
        .I1(\sr[4]_i_20_0 ),
        .I2(\sr[4]_i_101_n_0 ),
        .I3(\sr[4]_i_20_1 ),
        .I4(\tr_reg[5] ),
        .I5(\sr[4]_i_102_n_0 ),
        .O(\sr[4]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_46 
       (.I0(\sr[4]_i_21_2 ),
        .I1(\sr[4]_i_104_n_0 ),
        .I2(\sr[4]_i_21_3 ),
        .I3(\sr[4]_i_21_4 ),
        .I4(\sr[4]_i_106_n_0 ),
        .I5(grn27_n_15),
        .O(\sr[4]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAE00AE00AE00AEAE)) 
    \sr[4]_i_47 
       (.I0(\sr[4]_i_107_n_0 ),
        .I1(\sr[4]_i_108_n_0 ),
        .I2(grn27_n_37),
        .I3(\sr[4]_i_21_1 ),
        .I4(\sr[4]_i_110_n_0 ),
        .I5(grn27_n_11),
        .O(\sr[4]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \sr[4]_i_5 
       (.I0(\sr[4]_i_16_n_0 ),
        .I1(\sr_reg[4] ),
        .I2(\sr_reg[4]_0 ),
        .I3(\sr[4]_i_19_n_0 ),
        .I4(\sr[4]_i_20_n_0 ),
        .I5(\sr[4]_i_21_n_0 ),
        .O(\sr[4]_i_21_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_50 
       (.I0(\sr_reg[6]_8 [1]),
        .I1(\art/add/iv[7]_i_32 [2]),
        .I2(\art/add/sr[5]_i_18 [2]),
        .I3(\art/add/sr[5]_i_14 [1]),
        .O(\sr[4]_i_50_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[4]_i_51 
       (.I0(\art/add/sr[5]_i_18 [3]),
        .I1(\art/add/iv[7]_i_32 [3]),
        .I2(\art/add/sr[5]_i_14 [2]),
        .I3(\sr_reg[6]_8 [3]),
        .I4(\sr[4]_i_113_n_0 ),
        .O(\sr[4]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F000F0D0F08)) 
    \sr[4]_i_52 
       (.I0(\iv[0]_i_10_0 ),
        .I1(\iv[13]_i_36_n_0 ),
        .I2(\sr[4]_i_45_2 ),
        .I3(\iv[4]_i_34_n_0 ),
        .I4(\iv[12]_i_35_n_0 ),
        .I5(\sr_reg[8]_9 ),
        .O(\sr[4]_i_52_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_53 
       (.I0(\iv[4]_i_18_n_0 ),
        .I1(bbus_0[1]),
        .O(\sr[4]_i_53_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_55 
       (.I0(\tr_reg[5] ),
        .I1(\iv[4]_i_18_n_0 ),
        .O(\sr[4]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \sr[4]_i_56 
       (.I0(\sr[4]_i_36_0 ),
        .I1(\sr[4]_i_36 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\sr_reg[8]_42 ),
        .I4(\tr[20]_i_16_n_0 ),
        .I5(\tr[30]_i_3_4 ),
        .O(\sr[4]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h0F000F000F0D0F08)) 
    \sr[4]_i_57 
       (.I0(\iv[0]_i_10_0 ),
        .I1(\sr_reg[8]_77 ),
        .I2(\sr[4]_i_45_2 ),
        .I3(\iv[5]_i_33_n_0 ),
        .I4(\iv[13]_i_37_n_0 ),
        .I5(\sr_reg[8]_9 ),
        .O(\sr[4]_i_57_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[4]_i_58 
       (.I0(\iv[5]_i_18_n_0 ),
        .I1(bbus_0[1]),
        .O(\sr[4]_i_58_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_60 
       (.I0(\tr_reg[5] ),
        .I1(\iv[5]_i_18_n_0 ),
        .O(\sr[4]_i_60_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \sr[4]_i_61 
       (.I0(\tr[21]_i_15_n_0 ),
        .I1(\tr[30]_i_3_4 ),
        .I2(\sr[4]_i_36_0 ),
        .I3(\sr[4]_i_36 ),
        .I4(\sr_reg[8]_3 ),
        .I5(\iv[5]_i_23 ),
        .O(\sr[4]_i_61_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_62 
       (.I0(\sr[4]_i_45_2 ),
        .I1(\sr[4]_i_35_0 ),
        .I2(\iv[10]_i_35_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_61 ),
        .I5(\sr_reg[8]_9 ),
        .O(\sr[4]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_63 
       (.I0(\sr[4]_i_17_0 ),
        .I1(bbus_0[1]),
        .I2(\sr_reg[8]_17 ),
        .I3(\iv[13]_i_17_0 ),
        .I4(\sr_reg[8]_3 ),
        .I5(\sr[4]_i_114_n_0 ),
        .O(\sr[4]_i_63_n_0 ));
  LUT6 #(
    .INIT(64'h0001F00100F1F0F1)) 
    \sr[4]_i_65 
       (.I0(\sr_reg[8]_17 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[13]_i_17_0 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\tr[27]_i_3_0 ),
        .I5(\iv[10]_i_24_n_0 ),
        .O(\sr[4]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hDFDDCFCCDFDDFFFF)) 
    \sr[4]_i_68 
       (.I0(\sr[4]_i_37 ),
        .I1(\sr[4]_i_118_n_0 ),
        .I2(\tr[26]_i_3_0 ),
        .I3(grn27_n_13),
        .I4(\tr_reg[5] ),
        .I5(\sr_reg[8]_25 ),
        .O(\sr[4]_i_116_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_70 
       (.I0(\tr_reg[5] ),
        .I1(\sr[4]_i_38_1 ),
        .O(\sr[4]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_71 
       (.I0(\iv[15]_i_8 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\iv[6]_i_30_n_0 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\iv[6]_i_29_n_0 ),
        .I5(\tr[16]_i_6_2 ),
        .O(\sr[4]_i_71_n_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \sr[4]_i_72 
       (.I0(\sr[4]_i_38_1 ),
        .I1(bbus_0[1]),
        .I2(\tr[22]_i_3_0 ),
        .I3(\iv[13]_i_17_0 ),
        .I4(\sr_reg[8]_3 ),
        .I5(\sr[4]_i_122_n_0 ),
        .O(\sr[4]_i_72_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFF47FF47FF47)) 
    \sr[4]_i_76 
       (.I0(\sr[4]_i_39 ),
        .I1(\tr_reg[5] ),
        .I2(\sr[4]_i_39_0 ),
        .I3(\sr[4]_i_127_n_0 ),
        .I4(\iv[8]_i_26_n_0 ),
        .I5(grn27_n_13),
        .O(\iv[13]_i_27 ));
  LUT6 #(
    .INIT(64'hFF47FF47FF47FFFF)) 
    \sr[4]_i_80 
       (.I0(\sr[4]_i_40 ),
        .I1(\tr_reg[5] ),
        .I2(\sr_reg[8]_22 ),
        .I3(\sr[4]_i_134_n_0 ),
        .I4(\iv[14]_i_35_0 ),
        .I5(\sr_reg[8]_9 ),
        .O(\iv[8]_i_20 ));
  LUT6 #(
    .INIT(64'h111F111FFFFF111F)) 
    \sr[4]_i_82 
       (.I0(grn27_n_8),
        .I1(\tr_reg[5] ),
        .I2(\sr_reg[8]_9 ),
        .I3(\tr[17]_i_3_1 ),
        .I4(grn27_n_13),
        .I5(\iv[1]_i_25_n_0 ),
        .O(\sr[4]_i_82_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_83 
       (.I0(\tr_reg[5] ),
        .I1(\iv[1]_i_18_n_0 ),
        .O(\sr[4]_i_83_n_0 ));
  LUT4 #(
    .INIT(16'h00B8)) 
    \sr[4]_i_85 
       (.I0(\iv[1]_i_18_n_0 ),
        .I1(bbus_0[1]),
        .I2(grn27_n_8),
        .I3(\sr[4]_i_41_0 ),
        .O(\sr[4]_i_85_n_0 ));
  LUT5 #(
    .INIT(32'hF4F4FFF4)) 
    \sr[4]_i_89 
       (.I0(\sr[4]_i_42 ),
        .I1(\tr_reg[5] ),
        .I2(\sr[4]_i_142_n_0 ),
        .I3(grn27_n_13),
        .I4(\iv[7]_i_37_n_0 ),
        .O(\iv[7]_i_37_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_92 
       (.I0(\iv[15]_i_8 ),
        .I1(\sr[4]_i_43_1 ),
        .I2(\iv[11]_i_31_n_0 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\iv[11]_i_30_n_0 ),
        .I5(\tr[16]_i_6_2 ),
        .O(\sr_reg[8]_124 ));
  LUT6 #(
    .INIT(64'hDFDDCFCCDFDDFFFF)) 
    \sr[4]_i_93 
       (.I0(\sr[4]_i_43 ),
        .I1(\sr[4]_i_149_n_0 ),
        .I2(\sr[4]_i_43_0 ),
        .I3(grn27_n_13),
        .I4(\tr_reg[5] ),
        .I5(\sr_reg[8]_6 ),
        .O(\sr[4]_i_147_0 ));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_95 
       (.I0(\sr[4]_i_45_2 ),
        .I1(\sr[4]_i_44_1 ),
        .I2(\iv[12]_i_35_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_59 ),
        .I5(\sr_reg[8]_9 ),
        .O(\sr[4]_i_95_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_97 
       (.I0(\iv[15]_i_8 ),
        .I1(\sr[4]_i_44_2 ),
        .I2(\iv[12]_i_30_n_0 ),
        .I3(\sr_reg[8]_3 ),
        .I4(\iv[12]_i_29_n_0 ),
        .I5(\tr[16]_i_6_2 ),
        .O(\sr[4]_i_97_n_0 ));
  LUT6 #(
    .INIT(64'h350035003500350F)) 
    \sr[4]_i_98 
       (.I0(\iv[12]_i_25_n_0 ),
        .I1(\tr[29]_i_3_0 ),
        .I2(\sr_reg[8]_3 ),
        .I3(\iv[13]_i_17_0 ),
        .I4(\sr[4]_i_44_0 ),
        .I5(\tr_reg[5] ),
        .O(\sr[4]_i_98_n_0 ));
  LUT6 #(
    .INIT(64'h4444444454555444)) 
    \sr[4]_i_99 
       (.I0(\sr[4]_i_45_2 ),
        .I1(\sr[4]_i_45_0 ),
        .I2(\iv[13]_i_37_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\iv[13]_i_36_n_0 ),
        .I5(\sr_reg[8]_9 ),
        .O(\sr[4]_i_99_n_0 ));
  LUT6 #(
    .INIT(64'h08080F080D0D0F08)) 
    \sr[6]_i_10 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr[6]_i_4 ),
        .I2(\tr[24]_i_3_2 ),
        .I3(\sr[6]_i_27_n_0 ),
        .I4(\iv[13]_i_17_0 ),
        .I5(\sr[6]_i_28_n_0 ),
        .O(\sr_reg[8]_126 ));
  LUT6 #(
    .INIT(64'h000F0E0E000F000E)) 
    \sr[6]_i_12 
       (.I0(\sr_reg[8]_3 ),
        .I1(\sr[6]_i_27_n_0 ),
        .I2(\tr[16]_i_12_n_0 ),
        .I3(\tr[16]_i_13_n_0 ),
        .I4(\iv[13]_i_17_0 ),
        .I5(\sr[4]_i_36 ),
        .O(\sr_reg[8]_53 ));
  LUT5 #(
    .INIT(32'h11113111)) 
    \sr[6]_i_27 
       (.I0(\sr[6]_i_35_n_0 ),
        .I1(\sr_reg[8]_3 ),
        .I2(\sr[6]_i_12_0 ),
        .I3(\sr[6]_i_12_1 ),
        .I4(\sr[6]_i_12_2 ),
        .O(\sr[6]_i_27_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_28 
       (.I0(\sr_reg[8]_112 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_55 ),
        .O(\sr[6]_i_28_n_0 ));
  LUT4 #(
    .INIT(16'h444F)) 
    \sr[6]_i_30 
       (.I0(\tr[16]_i_28_n_0 ),
        .I1(\sr_reg[8]_3 ),
        .I2(\sr[6]_i_11 ),
        .I3(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_71 ));
  LUT5 #(
    .INIT(32'hB800B8FF)) 
    \sr[6]_i_34 
       (.I0(\tr[19]_i_3_3 ),
        .I1(\tr_reg[0] ),
        .I2(\tr[18]_i_3_2 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\badr[16]_INST_0_i_1 ),
        .O(\sr_reg[8]_117 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[6]_i_35 
       (.I0(\sr[6]_i_39_n_0 ),
        .I1(\iv[0]_i_19 ),
        .I2(\sr[6]_i_40_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_55 ),
        .O(\sr[6]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_39 
       (.I0(\iv[14]_i_62_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[14]_i_59_n_0 ),
        .O(\sr[6]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF077)) 
    \sr[6]_i_40 
       (.I0(\abus_o[3] [0]),
        .I1(\tr_reg[0] ),
        .I2(\iv[14]_i_60_n_0 ),
        .I3(\sr_reg[8]_93 ),
        .O(\sr[6]_i_40_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \sr[7]_i_10 
       (.I0(\tr[24]_i_3_2 ),
        .I1(\sr[7]_i_17_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\sr[7]_i_7 ),
        .O(\sr_reg[8]_123 ));
  LUT4 #(
    .INIT(16'hB800)) 
    \sr[7]_i_11 
       (.I0(\sr_reg[8]_65 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_4 ),
        .I3(\sr_reg[8]_36 ),
        .O(\sr_reg[8]_127 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[7]_i_17 
       (.I0(\sr_reg[8]_118 ),
        .I1(\iv[0]_i_19 ),
        .I2(\sr_reg[6]_7 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_52 ),
        .O(\sr[7]_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[7]_i_19 
       (.I0(\sr[7]_i_34_n_0 ),
        .I1(\sr[7]_i_35_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr[7]_i_36_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\badr[14]_INST_0_i_1 ),
        .O(\sr_reg[8]_65 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[7]_i_21 
       (.I0(\badr[0]_INST_0_i_1_0 ),
        .I1(\sr[7]_i_41_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\sr[7]_i_42_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\sr[7]_i_43_n_0 ),
        .O(\sr_reg[8]_4 ));
  LUT3 #(
    .INIT(8'h20)) 
    \sr[7]_i_22 
       (.I0(bbus_0[1]),
        .I1(\tr_reg[5] ),
        .I2(\niho_dsp_a[16] [3]),
        .O(\sr_reg[8]_36 ));
  LUT2 #(
    .INIT(4'hB)) 
    \sr[7]_i_24 
       (.I0(\sr_reg[8]_1 ),
        .I1(\sr[6]_i_12_0 ),
        .O(\sr_reg[8]_89 ));
  LUT4 #(
    .INIT(16'h8FFF)) 
    \sr[7]_i_25 
       (.I0(\sr_reg[8]_1 ),
        .I1(\sr[4]_i_36 ),
        .I2(\sr[4]_i_36_0 ),
        .I3(\sr[6]_i_12_1 ),
        .O(\sr_reg[8]_90 ));
  LUT5 #(
    .INIT(32'h88BB8B8B)) 
    \sr[7]_i_33 
       (.I0(\iv[15]_i_155_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\sr[4]_i_36 ),
        .I3(\niho_dsp_a[16] [2]),
        .I4(\tr_reg[0] ),
        .O(\sr_reg[6]_7 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_34 
       (.I0(\abus_o[11] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [0]),
        .O(\sr[7]_i_34_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_35 
       (.I0(\abus_o[11] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[11] [2]),
        .O(\sr[7]_i_35_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_36 
       (.I0(DI[1]),
        .I1(\tr_reg[0] ),
        .I2(DI[0]),
        .O(\sr[7]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'h57DFA820)) 
    \sr[7]_i_37 
       (.I0(\tr_reg[0] ),
        .I1(\niho_dsp_a[16] [3]),
        .I2(bbus_0[1]),
        .I3(\tr_reg[5] ),
        .I4(bbus_0[0]),
        .O(\sr_reg[8]_93 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_38 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(DI[2]),
        .O(\badr[14]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_40 
       (.I0(\abus_o[3] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [0]),
        .O(\badr[0]_INST_0_i_1_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_41 
       (.I0(\abus_o[3] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[3] [2]),
        .O(\sr[7]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_42 
       (.I0(\abus_o[7] [1]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [0]),
        .O(\sr[7]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h1D)) 
    \sr[7]_i_43 
       (.I0(\abus_o[7] [3]),
        .I1(\tr_reg[0] ),
        .I2(\abus_o[7] [2]),
        .O(\sr[7]_i_43_n_0 ));
  CARRY4 \sr_reg[5]_i_10 
       (.CI(\iv_reg[7]_i_12_n_0 ),
        .CO({\sr_reg[5]_i_10_n_0 ,\sr_reg[5]_i_10_n_1 ,\sr_reg[5]_i_10_n_2 ,\sr_reg[5]_i_10_n_3 }),
        .CYINIT(\<const0> ),
        .DI(\abus_o[11] ),
        .O(\art/add/sr[5]_i_18 ),
        .S(\iv[8]_i_8 ));
  CARRY4 \sr_reg[5]_i_5 
       (.CI(\sr_reg[5]_i_10_n_0 ),
        .CO({CO,\sr_reg[5]_i_5_n_1 ,\sr_reg[5]_i_5_n_2 ,\sr_reg[5]_i_5_n_3 }),
        .CYINIT(\<const0> ),
        .DI(DI),
        .O(\art/add/sr[5]_i_14 ),
        .S(S));
  LUT3 #(
    .INIT(8'h53)) 
    \tr[16]_i_10 
       (.I0(\tr_reg[5] ),
        .I1(bbus_0[1]),
        .I2(\niho_dsp_a[16] [3]),
        .O(\sr_reg[8]_35 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[16]_i_12 
       (.I0(\sr[6]_i_28_n_0 ),
        .I1(\sr_reg[8]_9 ),
        .O(\tr[16]_i_12_n_0 ));
  LUT3 #(
    .INIT(8'h70)) 
    \tr[16]_i_13 
       (.I0(\iv[13]_i_17_0 ),
        .I1(DI[3]),
        .I2(\sr_reg[8]_3 ),
        .O(\tr[16]_i_13_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \tr[16]_i_15 
       (.I0(\tr[16]_i_26_n_0 ),
        .I1(\iv[13]_i_17_0 ),
        .I2(\sr_reg[8]_0 ),
        .O(\tr[16]_i_9_0 ));
  LUT6 #(
    .INIT(64'hAA88AF88FA88FF88)) 
    \tr[16]_i_16 
       (.I0(\tr_reg[5] ),
        .I1(\tr[16]_i_6_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\iv[13]_i_17_0 ),
        .I4(\tr[16]_i_28_n_0 ),
        .I5(\tr[16]_i_6_1 ),
        .O(\tr[16]_i_16_n_0 ));
  LUT5 #(
    .INIT(32'h0000EEFE)) 
    \tr[16]_i_17 
       (.I0(\tr[16]_i_6_0 ),
        .I1(\tr[16]_i_6_2 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\sr[6]_i_28_n_0 ),
        .I4(\tr[16]_i_6_3 ),
        .O(\tr[16]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \tr[16]_i_2 
       (.I0(\tr_reg[1] ),
        .I1(\tr_reg[16] ),
        .I2(\tr[16]_i_5_n_0 ),
        .I3(\tr[16]_i_6_n_0 ),
        .I4(\tr_reg[1]_0 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \tr[16]_i_24 
       (.I0(\iv[14]_i_45_n_0 ),
        .I1(\tr[16]_i_32_n_0 ),
        .I2(\iv[0]_i_19 ),
        .I3(\iv[14]_i_43_n_0 ),
        .I4(\sr_reg[8]_93 ),
        .I5(\iv[14]_i_44_n_0 ),
        .O(\tr[16]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \tr[16]_i_26 
       (.I0(\sr_reg[8]_113 ),
        .I1(\iv[0]_i_19 ),
        .I2(\sr_reg[6]_6 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_49 ),
        .O(\tr[16]_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hE4FFE400)) 
    \tr[16]_i_28 
       (.I0(\iv[0]_i_19 ),
        .I1(\iv[7]_i_46_n_0 ),
        .I2(\sr_reg[8]_113 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_49 ),
        .O(\tr[16]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[16]_i_31 
       (.I0(\abus_o[11] [0]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_5 ));
  LUT3 #(
    .INIT(8'h47)) 
    \tr[16]_i_32 
       (.I0(DI[3]),
        .I1(\tr_reg[0] ),
        .I2(\tr[17]_i_3_0 ),
        .O(\tr[16]_i_32_n_0 ));
  LUT6 #(
    .INIT(64'h00001010000000FF)) 
    \tr[16]_i_5 
       (.I0(\tr[16]_i_12_n_0 ),
        .I1(\tr[16]_i_13_n_0 ),
        .I2(\tr[16]_i_2_0 ),
        .I3(\tr[16]_i_9_0 ),
        .I4(\niho_dsp_a[16] [3]),
        .I5(bbus_0[1]),
        .O(\tr[16]_i_5_n_0 ));
  LUT6 #(
    .INIT(64'h55FF55FF545454FF)) 
    \tr[16]_i_6 
       (.I0(\tr[16]_i_16_n_0 ),
        .I1(\sr_reg[8]_0 ),
        .I2(\iv[13]_i_17_0 ),
        .I3(\tr[16]_i_17_n_0 ),
        .I4(\niho_dsp_a[16] [3]),
        .I5(\tr_reg[5] ),
        .O(\tr[16]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \tr[16]_i_9 
       (.I0(\iv[0]_i_10_1 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[16]_i_24_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_49 ),
        .O(\sr_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \tr[17]_i_16 
       (.I0(\sr_reg[8]_91 ),
        .I1(\iv[0]_i_19 ),
        .I2(\iv[8]_i_41_n_0 ),
        .I3(\sr[4]_i_89_0 ),
        .I4(\sr_reg[8]_50 ),
        .O(\tr[17]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[17]_i_17 
       (.I0(\abus_o[11] [1]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_4 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[17]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[17]_i_6_n_0 ),
        .I2(\tr[17]_i_7_n_0 ),
        .I3(\tr[17]_i_2 ),
        .I4(\tr[17]_i_9_n_0 ),
        .O(\tr[17]_i_9_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47FF47FF)) 
    \tr[17]_i_6 
       (.I0(\iv[0]_i_17_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[17]_i_3_2 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[17]_i_3_0 ),
        .I5(\tr[24]_i_3_2 ),
        .O(\tr[17]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[17]_i_7 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\tr[17]_i_3_1 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\tr[17]_i_16_n_0 ),
        .O(\tr[17]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \tr[17]_i_9 
       (.I0(\sr_reg[8]_35 ),
        .I1(grn27_n_30),
        .I2(\tr[17]_i_16_n_0 ),
        .I3(\tr[19]_i_3_4 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\tr[17]_i_3_3 ),
        .O(\tr[17]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[18]_i_16 
       (.I0(\abus_o[11] [2]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_3 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[18]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[18]_i_2 ),
        .I2(\tr[18]_i_7_n_0 ),
        .I3(\tr[18]_i_8_n_0 ),
        .I4(\tr[18]_i_9_n_0 ),
        .O(\tr[18]_i_9_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \tr[18]_i_7 
       (.I0(\sr_reg[8]_35 ),
        .I1(grn27_n_33),
        .I2(\iv[1]_i_25_n_0 ),
        .I3(\tr[19]_i_3_4 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\tr[18]_i_3_3 ),
        .O(\tr[18]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[18]_i_8 
       (.I0(\sr_reg[8]_30 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[18]_i_3_1 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[18]_i_3_2 ),
        .I5(\tr[24]_i_3_2 ),
        .O(\tr[18]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[18]_i_9 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\tr[18]_i_3_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\iv[1]_i_25_n_0 ),
        .O(\tr[18]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[19]_i_15 
       (.I0(\abus_o[11] [3]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_2 ));
  LUT5 #(
    .INIT(32'hFFFFFF75)) 
    \tr[19]_i_2 
       (.I0(\tr[19]_i_3_n_0 ),
        .I1(\tr_reg[27] ),
        .I2(niho_dsp_c[0]),
        .I3(\tr_reg[19] ),
        .I4(\tr_reg[19]_0 ),
        .O(p_2_in[0]));
  LUT5 #(
    .INIT(32'hDDD0FFFF)) 
    \tr[19]_i_3 
       (.I0(\tr[19]_i_6_n_0 ),
        .I1(\tr[19]_i_7_n_0 ),
        .I2(\tr[19]_i_2_0 ),
        .I3(\tr[19]_i_9_n_0 ),
        .I4(\tr_reg[1] ),
        .O(\tr[19]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47FF47FF)) 
    \tr[19]_i_6 
       (.I0(\sr_reg[8]_33 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[19]_i_3_2 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[19]_i_3_3 ),
        .I5(\tr[24]_i_3_2 ),
        .O(\tr[19]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[19]_i_7 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\tr[19]_i_3_1 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\iv[2]_i_26_n_0 ),
        .O(\tr[19]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h88FFA0A088FFA0FF)) 
    \tr[19]_i_9 
       (.I0(\sr_reg[8]_35 ),
        .I1(\tr[19]_i_3_0 ),
        .I2(\iv[2]_i_26_n_0 ),
        .I3(\tr[19]_i_3_4 ),
        .I4(\sr_reg[8]_1 ),
        .I5(\tr[19]_i_3_5 ),
        .O(\tr[19]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hBBB888B8FFFFFFFF)) 
    \tr[20]_i_16 
       (.I0(\tr[20]_i_19_n_0 ),
        .I1(\iv[0]_i_19 ),
        .I2(\iv[14]_i_46_n_0 ),
        .I3(\sr_reg[8]_93 ),
        .I4(\iv[14]_i_48_n_0 ),
        .I5(\sr[4]_i_89_0 ),
        .O(\tr[20]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[20]_i_18 
       (.I0(DI[0]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_1 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \tr[20]_i_19 
       (.I0(bbus_0[0]),
        .I1(\abus_o[3] [0]),
        .I2(\tr_reg[0] ),
        .O(\tr[20]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[20]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[20]_i_2 ),
        .I2(\tr[20]_i_7_n_0 ),
        .I3(\tr[20]_i_8_n_0 ),
        .I4(\tr[20]_i_9_n_0 ),
        .O(\tr[20]_i_9_0 ));
  LUT5 #(
    .INIT(32'hFFFFA280)) 
    \tr[20]_i_7 
       (.I0(\sr_reg[8]_35 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[20]_i_16_n_0 ),
        .I3(\iv[3]_i_30_n_0 ),
        .I4(\tr[20]_i_3_3 ),
        .O(\tr[20]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000B800FF00B800)) 
    \tr[20]_i_8 
       (.I0(\sr_reg[8]_28 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[20]_i_3_1 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_2 ),
        .I5(\tr[20]_i_3_2 ),
        .O(\tr[20]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[20]_i_9 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\tr[20]_i_3_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\iv[3]_i_30_n_0 ),
        .O(\tr[20]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hEFECE3E0FFFFFFFF)) 
    \tr[21]_i_15 
       (.I0(\badr[0]_INST_0_i_1_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\sr[4]_i_61_0 ),
        .I3(\sr[7]_i_42_n_0 ),
        .I4(\sr[7]_i_41_n_0 ),
        .I5(\sr[4]_i_89_0 ),
        .O(\tr[21]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[21]_i_17 
       (.I0(DI[1]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[21]_i_2 
       (.I0(\tr[21]_i_3_n_0 ),
        .I1(\tr_reg[27] ),
        .I2(niho_dsp_c[1]),
        .I3(\tr_reg[21] ),
        .I4(\tr_reg[21]_0 ),
        .O(p_2_in[1]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[21]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[21]_i_2_0 ),
        .I2(\tr[21]_i_7_n_0 ),
        .I3(\tr[21]_i_8_n_0 ),
        .I4(\tr[21]_i_9_n_0 ),
        .O(\tr[21]_i_3_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA280)) 
    \tr[21]_i_7 
       (.I0(\sr_reg[8]_35 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[21]_i_15_n_0 ),
        .I3(\tr[21]_i_3_1 ),
        .I4(\tr[21]_i_3_4 ),
        .O(\tr[21]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[21]_i_8 
       (.I0(\iv[12]_i_27_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[21]_i_3_2 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[21]_i_3_3 ),
        .I5(\tr[24]_i_3_2 ),
        .O(\tr[21]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[21]_i_9 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\tr[21]_i_3_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\tr[21]_i_3_1 ),
        .O(\tr[21]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[22]_i_17 
       (.I0(DI[2]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[22]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[22]_i_6_n_0 ),
        .I2(\tr[22]_i_2 ),
        .I3(\tr[22]_i_8_n_0 ),
        .I4(\tr[22]_i_9_n_0 ),
        .O(\tr[22]_i_9_0 ));
  LUT5 #(
    .INIT(32'h11511555)) 
    \tr[22]_i_6 
       (.I0(\tr[26]_i_3_3 ),
        .I1(\sr_reg[8]_35 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\tr[22]_i_3_0 ),
        .I4(\iv[5]_i_28_n_0 ),
        .O(\tr[22]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[22]_i_8 
       (.I0(\iv[13]_i_29_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\iv[6]_i_29_n_0 ),
        .I3(\tr_reg[5] ),
        .I4(\iv[13]_i_17_1 ),
        .I5(\tr[24]_i_3_2 ),
        .O(\tr[22]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[22]_i_9 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\tr[22]_i_3_1 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\iv[5]_i_28_n_0 ),
        .O(\tr[22]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hEEEEE000)) 
    \tr[23]_i_10 
       (.I0(\tr[23]_i_3_2 ),
        .I1(\sr_reg[8]_1 ),
        .I2(grn27_n_3),
        .I3(\sr_reg[8]_35 ),
        .I4(\tr[30]_i_3_4 ),
        .O(\tr[23]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFBAFFFF)) 
    \tr[23]_i_2 
       (.I0(\tr[23]_i_3_n_0 ),
        .I1(\tr_reg[27] ),
        .I2(niho_dsp_c[2]),
        .I3(\tr_reg[23] ),
        .I4(\tr_reg[23]_0 ),
        .O(p_2_in[2]));
  LUT6 #(
    .INIT(64'h08080808080808AA)) 
    \tr[23]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[23]_i_6_n_0 ),
        .I2(\tr[23]_i_7_n_0 ),
        .I3(\tr[23]_i_2_0 ),
        .I4(\tr[23]_i_2_1 ),
        .I5(\tr[23]_i_10_n_0 ),
        .O(\tr[23]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47FF47FF)) 
    \tr[23]_i_6 
       (.I0(\iv[6]_i_30_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[23]_i_3_0 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[23]_i_3_1 ),
        .I5(\tr[24]_i_3_2 ),
        .O(\tr[23]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[23]_i_7 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[7]_i_38_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\tr[23]_i_3_2 ),
        .O(\tr[23]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[24]_i_10 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[8]_i_27_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\iv[7]_i_37_n_0 ),
        .O(\tr[24]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h000800080008AAAA)) 
    \tr[24]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[24]_i_6_n_0 ),
        .I2(\tr[24]_i_7_n_0 ),
        .I3(\tr[24]_i_2 ),
        .I4(\tr[24]_i_9_n_0 ),
        .I5(\tr[24]_i_10_n_0 ),
        .O(\tr[24]_i_10_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \tr[24]_i_6 
       (.I0(\sr_reg[8]_1 ),
        .I1(\tr[24]_i_3_3 ),
        .I2(\tr[19]_i_3_4 ),
        .O(\tr[24]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFB00FB00FB00)) 
    \tr[24]_i_7 
       (.I0(\tr[24]_i_3_4 ),
        .I1(\sr[4]_i_89_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\tr[24]_i_3_5 ),
        .I4(\tr[30]_i_3_4 ),
        .I5(\iv[7]_i_37_n_0 ),
        .O(\tr[24]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000FF00B800B800)) 
    \tr[24]_i_9 
       (.I0(\sr_reg[8]_26 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[24]_i_3_0 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_1 ),
        .I5(\tr[24]_i_3_2 ),
        .O(\tr[24]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'hFFC5)) 
    \tr[25]_i_10 
       (.I0(\iv[8]_i_26_n_0 ),
        .I1(\iv[9]_i_28_n_0 ),
        .I2(\sr_reg[8]_1 ),
        .I3(\tr_reg[5] ),
        .O(\tr[25]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h08AA080808AA08AA)) 
    \tr[25]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[25]_i_6_n_0 ),
        .I2(\tr[25]_i_7_n_0 ),
        .I3(\tr[25]_i_2 ),
        .I4(\tr[25]_i_9_n_0 ),
        .I5(\tr[25]_i_10_n_0 ),
        .O(\sr_reg[8]_31 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \tr[25]_i_6 
       (.I0(\tr[19]_i_3_4 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[25]_i_3_2 ),
        .O(\tr[25]_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFF8F8FFF8)) 
    \tr[25]_i_7 
       (.I0(\sr_reg[8]_36 ),
        .I1(grn27_n_27),
        .I2(\tr[26]_i_3_3 ),
        .I3(\tr[30]_i_3_4 ),
        .I4(\iv[8]_i_26_n_0 ),
        .I5(\tr[25]_i_3_3 ),
        .O(\tr[25]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFF001D0000001D00)) 
    \tr[25]_i_9 
       (.I0(\tr[25]_i_3_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\iv[8]_i_30 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_2 ),
        .I5(\tr[25]_i_3_1 ),
        .O(\tr[25]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[26]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[26]_i_6_n_0 ),
        .I2(\tr[26]_i_7_n_0 ),
        .I3(\tr[26]_i_2 ),
        .I4(\tr[26]_i_9_n_0 ),
        .O(\tr[26]_i_9_0 ));
  LUT6 #(
    .INIT(64'hFFFF47FF00FF47FF)) 
    \tr[26]_i_6 
       (.I0(\sr_reg[8]_29 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[26]_i_3_1 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_2 ),
        .I5(\tr[26]_i_3_2 ),
        .O(\tr[26]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[26]_i_7 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[10]_i_24_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\tr[26]_i_3_0 ),
        .O(\tr[26]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \tr[26]_i_9 
       (.I0(\sr_reg[8]_36 ),
        .I1(\sr_reg[8]_17 ),
        .I2(\tr[26]_i_3_3 ),
        .I3(\tr[26]_i_3_0 ),
        .I4(\tr[30]_i_3_4 ),
        .I5(\tr[26]_i_3_4 ),
        .O(\tr[26]_i_9_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[27]_i_17 
       (.I0(\abus_o[3] [3]),
        .I1(\tr[22]_i_11 ),
        .O(\iv[15]_i_108_7 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[27]_i_2 
       (.I0(\tr[27]_i_3_n_0 ),
        .I1(\tr_reg[27] ),
        .I2(niho_dsp_c[3]),
        .I3(\tr_reg[27]_0 ),
        .I4(\tr_reg[27]_1 ),
        .O(p_2_in[3]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[27]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[27]_i_6_n_0 ),
        .I2(\tr[27]_i_7_n_0 ),
        .I3(\tr[27]_i_2_0 ),
        .I4(\tr[27]_i_9_n_0 ),
        .O(\tr[27]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF47FF00FF47FF)) 
    \tr[27]_i_6 
       (.I0(\sr_reg[8]_32 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\iv[11]_i_30_n_0 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_2 ),
        .I5(\tr[27]_i_3_1 ),
        .O(\tr[27]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[27]_i_7 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[11]_i_26_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\tr[27]_i_3_0 ),
        .O(\tr[27]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8F8F8)) 
    \tr[27]_i_9 
       (.I0(\sr_reg[8]_36 ),
        .I1(\sr_reg[8]_7 ),
        .I2(\tr[26]_i_3_3 ),
        .I3(\tr[27]_i_3_0 ),
        .I4(\tr[30]_i_3_4 ),
        .I5(\tr[27]_i_3_2 ),
        .O(\tr[27]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[28]_i_2 
       (.I0(\tr[28]_i_3_n_0 ),
        .I1(\tr_reg[27] ),
        .I2(niho_dsp_c[4]),
        .I3(\tr_reg[28] ),
        .I4(\tr_reg[28]_0 ),
        .O(p_2_in[4]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[28]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[28]_i_6_n_0 ),
        .I2(\tr[28]_i_7_n_0 ),
        .I3(\tr[28]_i_2_0 ),
        .I4(\tr[28]_i_2_1 ),
        .O(\tr[28]_i_3_n_0 ));
  LUT6 #(
    .INIT(64'hFFFF47FF00FF47FF)) 
    \tr[28]_i_6 
       (.I0(\iv[11]_i_31_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\iv[12]_i_29_n_0 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_2 ),
        .I5(\tr[28]_i_3_0 ),
        .O(\tr[28]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[28]_i_7 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[12]_i_25_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\sr[4]_i_43_0 ),
        .O(\tr[28]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFBA)) 
    \tr[29]_i_2 
       (.I0(\tr[29]_i_3_n_0 ),
        .I1(\tr_reg[27] ),
        .I2(niho_dsp_c[5]),
        .I3(\tr_reg[29] ),
        .I4(\tr_reg[29]_0 ),
        .O(p_2_in[5]));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[29]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[29]_i_6_n_0 ),
        .I2(\tr[29]_i_7_n_0 ),
        .I3(\tr[29]_i_8_n_0 ),
        .I4(\tr[29]_i_9_n_0 ),
        .O(\tr[29]_i_3_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \tr[29]_i_6 
       (.I0(\tr[19]_i_3_4 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\tr[29]_i_3_2 ),
        .O(\tr[29]_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \tr[29]_i_7 
       (.I0(\tr[30]_i_3_4 ),
        .I1(\tr[29]_i_3_0 ),
        .I2(\tr[29]_i_3_3 ),
        .I3(\sr_reg[8]_36 ),
        .I4(\sr_reg[8]_13 ),
        .O(\tr[29]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'h0000B800FF00B800)) 
    \tr[29]_i_8 
       (.I0(\iv[12]_i_30_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\iv[13]_i_32_n_0 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_2 ),
        .I5(\tr[29]_i_3_1 ),
        .O(\tr[29]_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[29]_i_9 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[13]_i_25_n_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\tr[29]_i_3_0 ),
        .O(\tr[29]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hBABBBAAA)) 
    \tr[30]_i_10 
       (.I0(\tr[25]_i_2 ),
        .I1(\tr_reg[5] ),
        .I2(\iv[14]_i_35_0 ),
        .I3(\sr_reg[8]_1 ),
        .I4(\tr[30]_i_3_0 ),
        .O(\tr[30]_i_10_n_0 ));
  LUT5 #(
    .INIT(32'h080808AA)) 
    \tr[30]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\tr[30]_i_7_n_0 ),
        .I2(\tr[30]_i_8_n_0 ),
        .I3(\tr[30]_i_9_n_0 ),
        .I4(\tr[30]_i_10_n_0 ),
        .O(\tr[30]_i_10_0 ));
  LUT3 #(
    .INIT(8'hF4)) 
    \tr[30]_i_7 
       (.I0(\sr_reg[8]_1 ),
        .I1(\tr[30]_i_3_2 ),
        .I2(\tr[19]_i_3_4 ),
        .O(\tr[30]_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFF8F8F8)) 
    \tr[30]_i_8 
       (.I0(\sr_reg[8]_23 ),
        .I1(\sr_reg[8]_36 ),
        .I2(\tr[30]_i_3_3 ),
        .I3(\tr[30]_i_3_0 ),
        .I4(\tr[30]_i_3_4 ),
        .O(\tr[30]_i_8_n_0 ));
  LUT6 #(
    .INIT(64'h0000B800FF00B800)) 
    \tr[30]_i_9 
       (.I0(\iv[13]_i_31_n_0 ),
        .I1(\sr_reg[8]_1 ),
        .I2(\sr_reg[8]_27 ),
        .I3(\tr_reg[5] ),
        .I4(\tr[24]_i_3_2 ),
        .I5(\tr[30]_i_3_1 ),
        .O(\tr[30]_i_9_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank" *) 
module niho_rgf_bank_0
   (.out({gr21[15],gr21[14],gr21[13],gr21[12],gr21[11],gr21[10],gr21[9],gr21[8],gr21[7],gr21[6],gr21[5],gr21[4],gr21[3],gr21[2],gr21[1],gr21[0]}),
    .\grn_reg[15] ({gr22[15],gr22[14],gr22[13],gr22[12],gr22[11],gr22[10],gr22[9],gr22[8],gr22[7],gr22[6],gr22[5],gr22[4],gr22[3],gr22[2],gr22[1],gr22[0]}),
    .\grn_reg[15]_0 ({gr25[15],gr25[14],gr25[13],gr25[12],gr25[11],gr25[10],gr25[9],gr25[8],gr25[7],gr25[6],gr25[5],gr25[4],gr25[3],gr25[2],gr25[1],gr25[0]}),
    .\grn_reg[15]_1 ({gr26[15],gr26[14],gr26[13],gr26[12],gr26[11],gr26[10],gr26[9],gr26[8],gr26[7],gr26[6],gr26[5],gr26[4],gr26[3],gr26[2],gr26[1],gr26[0]}),
    SR,
    \grn_reg[15]_2 ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_3 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    \grn_reg[15]_4 ,
    \grn_reg[14]_1 ,
    \grn_reg[13]_1 ,
    \grn_reg[12]_1 ,
    \grn_reg[11]_1 ,
    \grn_reg[10]_1 ,
    \grn_reg[9]_1 ,
    \grn_reg[8]_1 ,
    \grn_reg[7]_1 ,
    \grn_reg[6]_1 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_1 ,
    \grn_reg[3]_1 ,
    \grn_reg[2]_1 ,
    \grn_reg[1]_1 ,
    \grn_reg[0]_1 ,
    \grn_reg[5]_2 ,
    \grn_reg[4]_2 ,
    \grn_reg[3]_2 ,
    \grn_reg[2]_2 ,
    \grn_reg[1]_2 ,
    \grn_reg[0]_2 ,
    \grn_reg[15]_5 ,
    \grn_reg[14]_2 ,
    \grn_reg[13]_2 ,
    \grn_reg[12]_2 ,
    \grn_reg[11]_2 ,
    \grn_reg[10]_2 ,
    \grn_reg[9]_2 ,
    \grn_reg[8]_2 ,
    \grn_reg[7]_2 ,
    \grn_reg[6]_2 ,
    \grn_reg[5]_3 ,
    \grn_reg[4]_3 ,
    \grn_reg[3]_3 ,
    \grn_reg[2]_3 ,
    \grn_reg[1]_3 ,
    \grn_reg[0]_3 ,
    \grn_reg[15]_6 ,
    \grn_reg[14]_3 ,
    \grn_reg[13]_3 ,
    \grn_reg[12]_3 ,
    \grn_reg[11]_3 ,
    \grn_reg[10]_3 ,
    \grn_reg[9]_3 ,
    \grn_reg[8]_3 ,
    \grn_reg[7]_3 ,
    \grn_reg[6]_3 ,
    \grn_reg[5]_4 ,
    \grn_reg[4]_4 ,
    \grn_reg[3]_4 ,
    \grn_reg[2]_4 ,
    \grn_reg[1]_4 ,
    \grn_reg[0]_4 ,
    \grn_reg[15]_7 ,
    \grn_reg[14]_4 ,
    \grn_reg[13]_4 ,
    \grn_reg[12]_4 ,
    \grn_reg[11]_4 ,
    \grn_reg[10]_4 ,
    \grn_reg[9]_4 ,
    \grn_reg[8]_4 ,
    \grn_reg[7]_4 ,
    \grn_reg[6]_4 ,
    \grn_reg[5]_5 ,
    \grn_reg[4]_5 ,
    \grn_reg[3]_5 ,
    \grn_reg[2]_5 ,
    \grn_reg[1]_5 ,
    \grn_reg[0]_5 ,
    \grn_reg[5]_6 ,
    \grn_reg[4]_6 ,
    \grn_reg[3]_6 ,
    \grn_reg[2]_6 ,
    \grn_reg[1]_6 ,
    \grn_reg[0]_6 ,
    \grn_reg[15]_8 ,
    \grn_reg[14]_5 ,
    \grn_reg[13]_5 ,
    \grn_reg[12]_5 ,
    \grn_reg[11]_5 ,
    \grn_reg[10]_5 ,
    \grn_reg[9]_5 ,
    \grn_reg[8]_5 ,
    \grn_reg[7]_5 ,
    \grn_reg[6]_5 ,
    \grn_reg[5]_7 ,
    \grn_reg[4]_7 ,
    \grn_reg[3]_7 ,
    \grn_reg[2]_7 ,
    \grn_reg[1]_7 ,
    \grn_reg[0]_7 ,
    \grn_reg[15]_9 ,
    \grn_reg[14]_6 ,
    \grn_reg[13]_6 ,
    \grn_reg[12]_6 ,
    \grn_reg[11]_6 ,
    \grn_reg[10]_6 ,
    \grn_reg[9]_6 ,
    \grn_reg[8]_6 ,
    \grn_reg[7]_6 ,
    \grn_reg[6]_6 ,
    \grn_reg[5]_8 ,
    \grn_reg[4]_8 ,
    \grn_reg[3]_8 ,
    \grn_reg[2]_8 ,
    \grn_reg[1]_8 ,
    \grn_reg[0]_8 ,
    \grn_reg[15]_10 ,
    \grn_reg[14]_7 ,
    \grn_reg[13]_7 ,
    \grn_reg[12]_7 ,
    \grn_reg[11]_7 ,
    \grn_reg[10]_7 ,
    \grn_reg[9]_7 ,
    \grn_reg[8]_7 ,
    \grn_reg[7]_7 ,
    \grn_reg[6]_7 ,
    \grn_reg[5]_9 ,
    \grn_reg[4]_9 ,
    \grn_reg[3]_9 ,
    \grn_reg[2]_9 ,
    \grn_reg[1]_9 ,
    \grn_reg[0]_9 ,
    \grn_reg[15]_11 ,
    \grn_reg[14]_8 ,
    \grn_reg[13]_8 ,
    \grn_reg[12]_8 ,
    \grn_reg[11]_8 ,
    \grn_reg[10]_8 ,
    \grn_reg[9]_8 ,
    \grn_reg[8]_8 ,
    \grn_reg[7]_8 ,
    \grn_reg[6]_8 ,
    \grn_reg[5]_10 ,
    \grn_reg[4]_10 ,
    \grn_reg[3]_10 ,
    \grn_reg[2]_10 ,
    \grn_reg[1]_10 ,
    \grn_reg[0]_10 ,
    rst_n,
    \i_/badr[15]_INST_0_i_20 ,
    abus_sel_0,
    \i_/badr[15]_INST_0_i_19 ,
    bbus_sel_0,
    \i_/bdatw[15]_INST_0_i_66 ,
    ctl_selb_rn,
    \i_/bdatw[15]_INST_0_i_66_0 ,
    \i_/bdatw[15]_INST_0_i_66_1 ,
    ctl_selb_0,
    \i_/bdatw[15]_INST_0_i_66_2 ,
    \i_/badr[15]_INST_0_i_17 ,
    \i_/bdatw[15]_INST_0_i_67 ,
    \i_/bdatw[15]_INST_0_i_27 ,
    \i_/bdatw[15]_INST_0_i_67_0 ,
    \i_/bdatw[15]_INST_0_i_27_0 ,
    \badr[31]_INST_0_i_1 ,
    \badr[30]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1 ,
    \badr[31]_INST_0_i_1_0 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1_0 ,
    \bdatw[31]_INST_0_i_5 ,
    \bdatw[30]_INST_0_i_3 ,
    \bdatw[29]_INST_0_i_3 ,
    \bdatw[28]_INST_0_i_3 ,
    \bdatw[27]_INST_0_i_3 ,
    \bdatw[26]_INST_0_i_3 ,
    \bdatw[25]_INST_0_i_3 ,
    \bdatw[24]_INST_0_i_3 ,
    \bdatw[23]_INST_0_i_3 ,
    \bdatw[22]_INST_0_i_3 ,
    \bdatw[21]_INST_0_i_3 ,
    \bdatw[20]_INST_0_i_3 ,
    \bdatw[19]_INST_0_i_3 ,
    \bdatw[18]_INST_0_i_3 ,
    \bdatw[17]_INST_0_i_3 ,
    \bdatw[16]_INST_0_i_3 ,
    \bdatw[31]_INST_0_i_5_0 ,
    \bdatw[30]_INST_0_i_3_0 ,
    \bdatw[29]_INST_0_i_3_0 ,
    \bdatw[28]_INST_0_i_3_0 ,
    \bdatw[27]_INST_0_i_3_0 ,
    \bdatw[26]_INST_0_i_3_0 ,
    \bdatw[25]_INST_0_i_3_0 ,
    \bdatw[24]_INST_0_i_3_0 ,
    \bdatw[23]_INST_0_i_3_0 ,
    \bdatw[22]_INST_0_i_3_0 ,
    \bdatw[21]_INST_0_i_3_0 ,
    \bdatw[20]_INST_0_i_3_0 ,
    \bdatw[19]_INST_0_i_3_0 ,
    \bdatw[18]_INST_0_i_3_0 ,
    \bdatw[17]_INST_0_i_3_0 ,
    \bdatw[16]_INST_0_i_3_0 ,
    \grn_reg[15]_12 ,
    cbus,
    clk,
    \grn_reg[15]_13 ,
    \grn_reg[15]_14 ,
    E,
    \grn_reg[15]_15 ,
    \grn_reg[0]_11 ,
    \grn_reg[15]_16 ,
    \grn_reg[15]_17 ,
    \grn_reg[15]_18 ,
    \grn_reg[15]_19 ,
    \grn_reg[15]_20 ,
    \grn_reg[15]_21 ,
    \grn_reg[0]_12 ,
    \grn_reg[15]_22 ,
    \grn_reg[0]_13 ,
    \grn_reg[15]_23 ,
    \grn_reg[15]_24 );
  output [0:0]SR;
  output \grn_reg[15]_2 ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_3 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  output \grn_reg[15]_4 ;
  output \grn_reg[14]_1 ;
  output \grn_reg[13]_1 ;
  output \grn_reg[12]_1 ;
  output \grn_reg[11]_1 ;
  output \grn_reg[10]_1 ;
  output \grn_reg[9]_1 ;
  output \grn_reg[8]_1 ;
  output \grn_reg[7]_1 ;
  output \grn_reg[6]_1 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_1 ;
  output \grn_reg[3]_1 ;
  output \grn_reg[2]_1 ;
  output \grn_reg[1]_1 ;
  output \grn_reg[0]_1 ;
  output \grn_reg[5]_2 ;
  output \grn_reg[4]_2 ;
  output \grn_reg[3]_2 ;
  output \grn_reg[2]_2 ;
  output \grn_reg[1]_2 ;
  output \grn_reg[0]_2 ;
  output \grn_reg[15]_5 ;
  output \grn_reg[14]_2 ;
  output \grn_reg[13]_2 ;
  output \grn_reg[12]_2 ;
  output \grn_reg[11]_2 ;
  output \grn_reg[10]_2 ;
  output \grn_reg[9]_2 ;
  output \grn_reg[8]_2 ;
  output \grn_reg[7]_2 ;
  output \grn_reg[6]_2 ;
  output \grn_reg[5]_3 ;
  output \grn_reg[4]_3 ;
  output \grn_reg[3]_3 ;
  output \grn_reg[2]_3 ;
  output \grn_reg[1]_3 ;
  output \grn_reg[0]_3 ;
  output \grn_reg[15]_6 ;
  output \grn_reg[14]_3 ;
  output \grn_reg[13]_3 ;
  output \grn_reg[12]_3 ;
  output \grn_reg[11]_3 ;
  output \grn_reg[10]_3 ;
  output \grn_reg[9]_3 ;
  output \grn_reg[8]_3 ;
  output \grn_reg[7]_3 ;
  output \grn_reg[6]_3 ;
  output \grn_reg[5]_4 ;
  output \grn_reg[4]_4 ;
  output \grn_reg[3]_4 ;
  output \grn_reg[2]_4 ;
  output \grn_reg[1]_4 ;
  output \grn_reg[0]_4 ;
  output \grn_reg[15]_7 ;
  output \grn_reg[14]_4 ;
  output \grn_reg[13]_4 ;
  output \grn_reg[12]_4 ;
  output \grn_reg[11]_4 ;
  output \grn_reg[10]_4 ;
  output \grn_reg[9]_4 ;
  output \grn_reg[8]_4 ;
  output \grn_reg[7]_4 ;
  output \grn_reg[6]_4 ;
  output \grn_reg[5]_5 ;
  output \grn_reg[4]_5 ;
  output \grn_reg[3]_5 ;
  output \grn_reg[2]_5 ;
  output \grn_reg[1]_5 ;
  output \grn_reg[0]_5 ;
  output \grn_reg[5]_6 ;
  output \grn_reg[4]_6 ;
  output \grn_reg[3]_6 ;
  output \grn_reg[2]_6 ;
  output \grn_reg[1]_6 ;
  output \grn_reg[0]_6 ;
  output \grn_reg[15]_8 ;
  output \grn_reg[14]_5 ;
  output \grn_reg[13]_5 ;
  output \grn_reg[12]_5 ;
  output \grn_reg[11]_5 ;
  output \grn_reg[10]_5 ;
  output \grn_reg[9]_5 ;
  output \grn_reg[8]_5 ;
  output \grn_reg[7]_5 ;
  output \grn_reg[6]_5 ;
  output \grn_reg[5]_7 ;
  output \grn_reg[4]_7 ;
  output \grn_reg[3]_7 ;
  output \grn_reg[2]_7 ;
  output \grn_reg[1]_7 ;
  output \grn_reg[0]_7 ;
  output \grn_reg[15]_9 ;
  output \grn_reg[14]_6 ;
  output \grn_reg[13]_6 ;
  output \grn_reg[12]_6 ;
  output \grn_reg[11]_6 ;
  output \grn_reg[10]_6 ;
  output \grn_reg[9]_6 ;
  output \grn_reg[8]_6 ;
  output \grn_reg[7]_6 ;
  output \grn_reg[6]_6 ;
  output \grn_reg[5]_8 ;
  output \grn_reg[4]_8 ;
  output \grn_reg[3]_8 ;
  output \grn_reg[2]_8 ;
  output \grn_reg[1]_8 ;
  output \grn_reg[0]_8 ;
  output \grn_reg[15]_10 ;
  output \grn_reg[14]_7 ;
  output \grn_reg[13]_7 ;
  output \grn_reg[12]_7 ;
  output \grn_reg[11]_7 ;
  output \grn_reg[10]_7 ;
  output \grn_reg[9]_7 ;
  output \grn_reg[8]_7 ;
  output \grn_reg[7]_7 ;
  output \grn_reg[6]_7 ;
  output \grn_reg[5]_9 ;
  output \grn_reg[4]_9 ;
  output \grn_reg[3]_9 ;
  output \grn_reg[2]_9 ;
  output \grn_reg[1]_9 ;
  output \grn_reg[0]_9 ;
  output \grn_reg[15]_11 ;
  output \grn_reg[14]_8 ;
  output \grn_reg[13]_8 ;
  output \grn_reg[12]_8 ;
  output \grn_reg[11]_8 ;
  output \grn_reg[10]_8 ;
  output \grn_reg[9]_8 ;
  output \grn_reg[8]_8 ;
  output \grn_reg[7]_8 ;
  output \grn_reg[6]_8 ;
  output \grn_reg[5]_10 ;
  output \grn_reg[4]_10 ;
  output \grn_reg[3]_10 ;
  output \grn_reg[2]_10 ;
  output \grn_reg[1]_10 ;
  output \grn_reg[0]_10 ;
  input rst_n;
  input [2:0]\i_/badr[15]_INST_0_i_20 ;
  input [7:0]abus_sel_0;
  input \i_/badr[15]_INST_0_i_19 ;
  input [5:0]bbus_sel_0;
  input \i_/bdatw[15]_INST_0_i_66 ;
  input [1:0]ctl_selb_rn;
  input \i_/bdatw[15]_INST_0_i_66_0 ;
  input \i_/bdatw[15]_INST_0_i_66_1 ;
  input [0:0]ctl_selb_0;
  input \i_/bdatw[15]_INST_0_i_66_2 ;
  input \i_/badr[15]_INST_0_i_17 ;
  input \i_/bdatw[15]_INST_0_i_67 ;
  input \i_/bdatw[15]_INST_0_i_27 ;
  input \i_/bdatw[15]_INST_0_i_67_0 ;
  input \i_/bdatw[15]_INST_0_i_27_0 ;
  input \badr[31]_INST_0_i_1 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1 ;
  input \badr[31]_INST_0_i_1_0 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1_0 ;
  input \bdatw[31]_INST_0_i_5 ;
  input \bdatw[30]_INST_0_i_3 ;
  input \bdatw[29]_INST_0_i_3 ;
  input \bdatw[28]_INST_0_i_3 ;
  input \bdatw[27]_INST_0_i_3 ;
  input \bdatw[26]_INST_0_i_3 ;
  input \bdatw[25]_INST_0_i_3 ;
  input \bdatw[24]_INST_0_i_3 ;
  input \bdatw[23]_INST_0_i_3 ;
  input \bdatw[22]_INST_0_i_3 ;
  input \bdatw[21]_INST_0_i_3 ;
  input \bdatw[20]_INST_0_i_3 ;
  input \bdatw[19]_INST_0_i_3 ;
  input \bdatw[18]_INST_0_i_3 ;
  input \bdatw[17]_INST_0_i_3 ;
  input \bdatw[16]_INST_0_i_3 ;
  input \bdatw[31]_INST_0_i_5_0 ;
  input \bdatw[30]_INST_0_i_3_0 ;
  input \bdatw[29]_INST_0_i_3_0 ;
  input \bdatw[28]_INST_0_i_3_0 ;
  input \bdatw[27]_INST_0_i_3_0 ;
  input \bdatw[26]_INST_0_i_3_0 ;
  input \bdatw[25]_INST_0_i_3_0 ;
  input \bdatw[24]_INST_0_i_3_0 ;
  input \bdatw[23]_INST_0_i_3_0 ;
  input \bdatw[22]_INST_0_i_3_0 ;
  input \bdatw[21]_INST_0_i_3_0 ;
  input \bdatw[20]_INST_0_i_3_0 ;
  input \bdatw[19]_INST_0_i_3_0 ;
  input \bdatw[18]_INST_0_i_3_0 ;
  input \bdatw[17]_INST_0_i_3_0 ;
  input \bdatw[16]_INST_0_i_3_0 ;
  input [0:0]\grn_reg[15]_12 ;
  input [15:0]cbus;
  input clk;
  input [0:0]\grn_reg[15]_13 ;
  input [0:0]\grn_reg[15]_14 ;
  input [0:0]E;
  input [0:0]\grn_reg[15]_15 ;
  input [0:0]\grn_reg[0]_11 ;
  input [0:0]\grn_reg[15]_16 ;
  input [0:0]\grn_reg[15]_17 ;
  input [0:0]\grn_reg[15]_18 ;
  input [15:0]\grn_reg[15]_19 ;
  input [0:0]\grn_reg[15]_20 ;
  input [0:0]\grn_reg[15]_21 ;
  input [0:0]\grn_reg[0]_12 ;
  input [0:0]\grn_reg[15]_22 ;
  input [0:0]\grn_reg[0]_13 ;
  input [0:0]\grn_reg[15]_23 ;
  input [0:0]\grn_reg[15]_24 ;
     output [15:0]gr21;
     output [15:0]gr22;
     output [15:0]gr25;
     output [15:0]gr26;

  wire [0:0]E;
  wire [0:0]SR;
  wire [7:0]abus_sel_0;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire \badr[31]_INST_0_i_1 ;
  wire \badr[31]_INST_0_i_1_0 ;
  wire [5:0]bbus_sel_0;
  wire \bdatw[16]_INST_0_i_3 ;
  wire \bdatw[16]_INST_0_i_3_0 ;
  wire \bdatw[17]_INST_0_i_3 ;
  wire \bdatw[17]_INST_0_i_3_0 ;
  wire \bdatw[18]_INST_0_i_3 ;
  wire \bdatw[18]_INST_0_i_3_0 ;
  wire \bdatw[19]_INST_0_i_3 ;
  wire \bdatw[19]_INST_0_i_3_0 ;
  wire \bdatw[20]_INST_0_i_3 ;
  wire \bdatw[20]_INST_0_i_3_0 ;
  wire \bdatw[21]_INST_0_i_3 ;
  wire \bdatw[21]_INST_0_i_3_0 ;
  wire \bdatw[22]_INST_0_i_3 ;
  wire \bdatw[22]_INST_0_i_3_0 ;
  wire \bdatw[23]_INST_0_i_3 ;
  wire \bdatw[23]_INST_0_i_3_0 ;
  wire \bdatw[24]_INST_0_i_3 ;
  wire \bdatw[24]_INST_0_i_3_0 ;
  wire \bdatw[25]_INST_0_i_3 ;
  wire \bdatw[25]_INST_0_i_3_0 ;
  wire \bdatw[26]_INST_0_i_3 ;
  wire \bdatw[26]_INST_0_i_3_0 ;
  wire \bdatw[27]_INST_0_i_3 ;
  wire \bdatw[27]_INST_0_i_3_0 ;
  wire \bdatw[28]_INST_0_i_3 ;
  wire \bdatw[28]_INST_0_i_3_0 ;
  wire \bdatw[29]_INST_0_i_3 ;
  wire \bdatw[29]_INST_0_i_3_0 ;
  wire \bdatw[30]_INST_0_i_3 ;
  wire \bdatw[30]_INST_0_i_3_0 ;
  wire \bdatw[31]_INST_0_i_5 ;
  wire \bdatw[31]_INST_0_i_5_0 ;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  (* DONT_TOUCH *) wire [15:0]gr00;
  (* DONT_TOUCH *) wire [15:0]gr01;
  (* DONT_TOUCH *) wire [15:0]gr02;
  (* DONT_TOUCH *) wire [15:0]gr03;
  (* DONT_TOUCH *) wire [15:0]gr04;
  (* DONT_TOUCH *) wire [15:0]gr05;
  (* DONT_TOUCH *) wire [15:0]gr06;
  (* DONT_TOUCH *) wire [15:0]gr07;
  (* DONT_TOUCH *) wire [15:0]gr20;
  (* DONT_TOUCH *) wire [15:0]gr21;
  (* DONT_TOUCH *) wire [15:0]gr22;
  (* DONT_TOUCH *) wire [15:0]gr23;
  (* DONT_TOUCH *) wire [15:0]gr24;
  (* DONT_TOUCH *) wire [15:0]gr25;
  (* DONT_TOUCH *) wire [15:0]gr26;
  (* DONT_TOUCH *) wire [15:0]gr27;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[0]_10 ;
  wire [0:0]\grn_reg[0]_11 ;
  wire [0:0]\grn_reg[0]_12 ;
  wire [0:0]\grn_reg[0]_13 ;
  wire \grn_reg[0]_2 ;
  wire \grn_reg[0]_3 ;
  wire \grn_reg[0]_4 ;
  wire \grn_reg[0]_5 ;
  wire \grn_reg[0]_6 ;
  wire \grn_reg[0]_7 ;
  wire \grn_reg[0]_8 ;
  wire \grn_reg[0]_9 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[10]_1 ;
  wire \grn_reg[10]_2 ;
  wire \grn_reg[10]_3 ;
  wire \grn_reg[10]_4 ;
  wire \grn_reg[10]_5 ;
  wire \grn_reg[10]_6 ;
  wire \grn_reg[10]_7 ;
  wire \grn_reg[10]_8 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[11]_1 ;
  wire \grn_reg[11]_2 ;
  wire \grn_reg[11]_3 ;
  wire \grn_reg[11]_4 ;
  wire \grn_reg[11]_5 ;
  wire \grn_reg[11]_6 ;
  wire \grn_reg[11]_7 ;
  wire \grn_reg[11]_8 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[12]_1 ;
  wire \grn_reg[12]_2 ;
  wire \grn_reg[12]_3 ;
  wire \grn_reg[12]_4 ;
  wire \grn_reg[12]_5 ;
  wire \grn_reg[12]_6 ;
  wire \grn_reg[12]_7 ;
  wire \grn_reg[12]_8 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[13]_1 ;
  wire \grn_reg[13]_2 ;
  wire \grn_reg[13]_3 ;
  wire \grn_reg[13]_4 ;
  wire \grn_reg[13]_5 ;
  wire \grn_reg[13]_6 ;
  wire \grn_reg[13]_7 ;
  wire \grn_reg[13]_8 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[14]_1 ;
  wire \grn_reg[14]_2 ;
  wire \grn_reg[14]_3 ;
  wire \grn_reg[14]_4 ;
  wire \grn_reg[14]_5 ;
  wire \grn_reg[14]_6 ;
  wire \grn_reg[14]_7 ;
  wire \grn_reg[14]_8 ;
  wire \grn_reg[15]_10 ;
  wire \grn_reg[15]_11 ;
  wire [0:0]\grn_reg[15]_12 ;
  wire [0:0]\grn_reg[15]_13 ;
  wire [0:0]\grn_reg[15]_14 ;
  wire [0:0]\grn_reg[15]_15 ;
  wire [0:0]\grn_reg[15]_16 ;
  wire [0:0]\grn_reg[15]_17 ;
  wire [0:0]\grn_reg[15]_18 ;
  wire [15:0]\grn_reg[15]_19 ;
  wire \grn_reg[15]_2 ;
  wire [0:0]\grn_reg[15]_20 ;
  wire [0:0]\grn_reg[15]_21 ;
  wire [0:0]\grn_reg[15]_22 ;
  wire [0:0]\grn_reg[15]_23 ;
  wire [0:0]\grn_reg[15]_24 ;
  wire \grn_reg[15]_3 ;
  wire \grn_reg[15]_4 ;
  wire \grn_reg[15]_5 ;
  wire \grn_reg[15]_6 ;
  wire \grn_reg[15]_7 ;
  wire \grn_reg[15]_8 ;
  wire \grn_reg[15]_9 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[1]_1 ;
  wire \grn_reg[1]_10 ;
  wire \grn_reg[1]_2 ;
  wire \grn_reg[1]_3 ;
  wire \grn_reg[1]_4 ;
  wire \grn_reg[1]_5 ;
  wire \grn_reg[1]_6 ;
  wire \grn_reg[1]_7 ;
  wire \grn_reg[1]_8 ;
  wire \grn_reg[1]_9 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[2]_1 ;
  wire \grn_reg[2]_10 ;
  wire \grn_reg[2]_2 ;
  wire \grn_reg[2]_3 ;
  wire \grn_reg[2]_4 ;
  wire \grn_reg[2]_5 ;
  wire \grn_reg[2]_6 ;
  wire \grn_reg[2]_7 ;
  wire \grn_reg[2]_8 ;
  wire \grn_reg[2]_9 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[3]_1 ;
  wire \grn_reg[3]_10 ;
  wire \grn_reg[3]_2 ;
  wire \grn_reg[3]_3 ;
  wire \grn_reg[3]_4 ;
  wire \grn_reg[3]_5 ;
  wire \grn_reg[3]_6 ;
  wire \grn_reg[3]_7 ;
  wire \grn_reg[3]_8 ;
  wire \grn_reg[3]_9 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[4]_1 ;
  wire \grn_reg[4]_10 ;
  wire \grn_reg[4]_2 ;
  wire \grn_reg[4]_3 ;
  wire \grn_reg[4]_4 ;
  wire \grn_reg[4]_5 ;
  wire \grn_reg[4]_6 ;
  wire \grn_reg[4]_7 ;
  wire \grn_reg[4]_8 ;
  wire \grn_reg[4]_9 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[5]_10 ;
  wire \grn_reg[5]_2 ;
  wire \grn_reg[5]_3 ;
  wire \grn_reg[5]_4 ;
  wire \grn_reg[5]_5 ;
  wire \grn_reg[5]_6 ;
  wire \grn_reg[5]_7 ;
  wire \grn_reg[5]_8 ;
  wire \grn_reg[5]_9 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[6]_1 ;
  wire \grn_reg[6]_2 ;
  wire \grn_reg[6]_3 ;
  wire \grn_reg[6]_4 ;
  wire \grn_reg[6]_5 ;
  wire \grn_reg[6]_6 ;
  wire \grn_reg[6]_7 ;
  wire \grn_reg[6]_8 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[7]_1 ;
  wire \grn_reg[7]_2 ;
  wire \grn_reg[7]_3 ;
  wire \grn_reg[7]_4 ;
  wire \grn_reg[7]_5 ;
  wire \grn_reg[7]_6 ;
  wire \grn_reg[7]_7 ;
  wire \grn_reg[7]_8 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[8]_1 ;
  wire \grn_reg[8]_2 ;
  wire \grn_reg[8]_3 ;
  wire \grn_reg[8]_4 ;
  wire \grn_reg[8]_5 ;
  wire \grn_reg[8]_6 ;
  wire \grn_reg[8]_7 ;
  wire \grn_reg[8]_8 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \grn_reg[9]_1 ;
  wire \grn_reg[9]_2 ;
  wire \grn_reg[9]_3 ;
  wire \grn_reg[9]_4 ;
  wire \grn_reg[9]_5 ;
  wire \grn_reg[9]_6 ;
  wire \grn_reg[9]_7 ;
  wire \grn_reg[9]_8 ;
  wire \i_/badr[15]_INST_0_i_17 ;
  wire \i_/badr[15]_INST_0_i_19 ;
  wire [2:0]\i_/badr[15]_INST_0_i_20 ;
  wire \i_/bdatw[15]_INST_0_i_27 ;
  wire \i_/bdatw[15]_INST_0_i_27_0 ;
  wire \i_/bdatw[15]_INST_0_i_66 ;
  wire \i_/bdatw[15]_INST_0_i_66_0 ;
  wire \i_/bdatw[15]_INST_0_i_66_1 ;
  wire \i_/bdatw[15]_INST_0_i_66_2 ;
  wire \i_/bdatw[15]_INST_0_i_67 ;
  wire \i_/bdatw[15]_INST_0_i_67_0 ;
  wire rst_n;

  niho_rgf_bank_bus abuso
       (.abus_sel_0(abus_sel_0),
        .\badr[15]_INST_0_i_5 (gr04),
        .\badr[15]_INST_0_i_5_0 (gr07),
        .\badr[15]_INST_0_i_5_1 (gr00),
        .\grn_reg[0] (\grn_reg[0] ),
        .\grn_reg[0]_0 (\grn_reg[0]_0 ),
        .\grn_reg[10] (\grn_reg[10] ),
        .\grn_reg[10]_0 (\grn_reg[10]_0 ),
        .\grn_reg[11] (\grn_reg[11] ),
        .\grn_reg[11]_0 (\grn_reg[11]_0 ),
        .\grn_reg[12] (\grn_reg[12] ),
        .\grn_reg[12]_0 (\grn_reg[12]_0 ),
        .\grn_reg[13] (\grn_reg[13] ),
        .\grn_reg[13]_0 (\grn_reg[13]_0 ),
        .\grn_reg[14] (\grn_reg[14] ),
        .\grn_reg[14]_0 (\grn_reg[14]_0 ),
        .\grn_reg[15] (\grn_reg[15]_2 ),
        .\grn_reg[15]_0 (\grn_reg[15]_3 ),
        .\grn_reg[1] (\grn_reg[1] ),
        .\grn_reg[1]_0 (\grn_reg[1]_0 ),
        .\grn_reg[2] (\grn_reg[2] ),
        .\grn_reg[2]_0 (\grn_reg[2]_0 ),
        .\grn_reg[3] (\grn_reg[3] ),
        .\grn_reg[3]_0 (\grn_reg[3]_0 ),
        .\grn_reg[4] (\grn_reg[4] ),
        .\grn_reg[4]_0 (\grn_reg[4]_0 ),
        .\grn_reg[5] (\grn_reg[5] ),
        .\grn_reg[5]_0 (\grn_reg[5]_0 ),
        .\grn_reg[6] (\grn_reg[6] ),
        .\grn_reg[6]_0 (\grn_reg[6]_0 ),
        .\grn_reg[7] (\grn_reg[7] ),
        .\grn_reg[7]_0 (\grn_reg[7]_0 ),
        .\grn_reg[8] (\grn_reg[8] ),
        .\grn_reg[8]_0 (\grn_reg[8]_0 ),
        .\grn_reg[9] (\grn_reg[9] ),
        .\grn_reg[9]_0 (\grn_reg[9]_0 ),
        .\i_/badr[15]_INST_0_i_19_0 (gr06),
        .\i_/badr[15]_INST_0_i_19_1 (gr05),
        .\i_/badr[15]_INST_0_i_19_2 (\i_/badr[15]_INST_0_i_19 ),
        .\i_/badr[15]_INST_0_i_20_0 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/badr[15]_INST_0_i_20_1 (gr02),
        .\i_/badr[15]_INST_0_i_20_2 (gr01),
        .out(gr03));
  niho_rgf_bank_bus_2 abuso2h
       (.abus_sel_0({abus_sel_0[7],abus_sel_0[4:3],abus_sel_0[0]}),
        .\badr[16]_INST_0_i_1 (\badr[16]_INST_0_i_1 ),
        .\badr[16]_INST_0_i_1_0 (\badr[16]_INST_0_i_1_0 ),
        .\badr[17]_INST_0_i_1 (\badr[17]_INST_0_i_1 ),
        .\badr[17]_INST_0_i_1_0 (\badr[17]_INST_0_i_1_0 ),
        .\badr[18]_INST_0_i_1 (\badr[18]_INST_0_i_1 ),
        .\badr[18]_INST_0_i_1_0 (\badr[18]_INST_0_i_1_0 ),
        .\badr[19]_INST_0_i_1 (\badr[19]_INST_0_i_1 ),
        .\badr[19]_INST_0_i_1_0 (\badr[19]_INST_0_i_1_0 ),
        .\badr[20]_INST_0_i_1 (\badr[20]_INST_0_i_1 ),
        .\badr[20]_INST_0_i_1_0 (\badr[20]_INST_0_i_1_0 ),
        .\badr[21]_INST_0_i_1 (\badr[21]_INST_0_i_1 ),
        .\badr[21]_INST_0_i_1_0 (\badr[21]_INST_0_i_1_0 ),
        .\badr[22]_INST_0_i_1 (\badr[22]_INST_0_i_1 ),
        .\badr[22]_INST_0_i_1_0 (\badr[22]_INST_0_i_1_0 ),
        .\badr[23]_INST_0_i_1 (\badr[23]_INST_0_i_1 ),
        .\badr[23]_INST_0_i_1_0 (\badr[23]_INST_0_i_1_0 ),
        .\badr[24]_INST_0_i_1 (\badr[24]_INST_0_i_1 ),
        .\badr[24]_INST_0_i_1_0 (\badr[24]_INST_0_i_1_0 ),
        .\badr[25]_INST_0_i_1 (\badr[25]_INST_0_i_1 ),
        .\badr[25]_INST_0_i_1_0 (\badr[25]_INST_0_i_1_0 ),
        .\badr[26]_INST_0_i_1 (\badr[26]_INST_0_i_1 ),
        .\badr[26]_INST_0_i_1_0 (\badr[26]_INST_0_i_1_0 ),
        .\badr[27]_INST_0_i_1 (\badr[27]_INST_0_i_1 ),
        .\badr[27]_INST_0_i_1_0 (\badr[27]_INST_0_i_1_0 ),
        .\badr[28]_INST_0_i_1 (\badr[28]_INST_0_i_1 ),
        .\badr[28]_INST_0_i_1_0 (\badr[28]_INST_0_i_1_0 ),
        .\badr[29]_INST_0_i_1 (\badr[29]_INST_0_i_1 ),
        .\badr[29]_INST_0_i_1_0 (\badr[29]_INST_0_i_1_0 ),
        .\badr[30]_INST_0_i_1 (\badr[30]_INST_0_i_1 ),
        .\badr[30]_INST_0_i_1_0 (\badr[30]_INST_0_i_1_0 ),
        .\badr[31]_INST_0_i_1 (gr20),
        .\badr[31]_INST_0_i_1_0 (\badr[31]_INST_0_i_1 ),
        .\badr[31]_INST_0_i_1_1 (gr23),
        .\badr[31]_INST_0_i_1_2 (gr24),
        .\badr[31]_INST_0_i_1_3 (\badr[31]_INST_0_i_1_0 ),
        .\grn_reg[0] (\grn_reg[0]_7 ),
        .\grn_reg[0]_0 (\grn_reg[0]_8 ),
        .\grn_reg[10] (\grn_reg[10]_5 ),
        .\grn_reg[10]_0 (\grn_reg[10]_6 ),
        .\grn_reg[11] (\grn_reg[11]_5 ),
        .\grn_reg[11]_0 (\grn_reg[11]_6 ),
        .\grn_reg[12] (\grn_reg[12]_5 ),
        .\grn_reg[12]_0 (\grn_reg[12]_6 ),
        .\grn_reg[13] (\grn_reg[13]_5 ),
        .\grn_reg[13]_0 (\grn_reg[13]_6 ),
        .\grn_reg[14] (\grn_reg[14]_5 ),
        .\grn_reg[14]_0 (\grn_reg[14]_6 ),
        .\grn_reg[15] (\grn_reg[15]_8 ),
        .\grn_reg[15]_0 (\grn_reg[15]_9 ),
        .\grn_reg[1] (\grn_reg[1]_7 ),
        .\grn_reg[1]_0 (\grn_reg[1]_8 ),
        .\grn_reg[2] (\grn_reg[2]_7 ),
        .\grn_reg[2]_0 (\grn_reg[2]_8 ),
        .\grn_reg[3] (\grn_reg[3]_7 ),
        .\grn_reg[3]_0 (\grn_reg[3]_8 ),
        .\grn_reg[4] (\grn_reg[4]_7 ),
        .\grn_reg[4]_0 (\grn_reg[4]_8 ),
        .\grn_reg[5] (\grn_reg[5]_7 ),
        .\grn_reg[5]_0 (\grn_reg[5]_8 ),
        .\grn_reg[6] (\grn_reg[6]_5 ),
        .\grn_reg[6]_0 (\grn_reg[6]_6 ),
        .\grn_reg[7] (\grn_reg[7]_5 ),
        .\grn_reg[7]_0 (\grn_reg[7]_6 ),
        .\grn_reg[8] (\grn_reg[8]_5 ),
        .\grn_reg[8]_0 (\grn_reg[8]_6 ),
        .\grn_reg[9] (\grn_reg[9]_5 ),
        .\grn_reg[9]_0 (\grn_reg[9]_6 ),
        .\i_/badr[31]_INST_0_i_7_0 ({\i_/badr[15]_INST_0_i_20 [2],\i_/badr[15]_INST_0_i_20 [0]}),
        .out(gr27));
  niho_rgf_bank_bus_3 abuso2l
       (.abus_sel_0(abus_sel_0),
        .\badr[15]_INST_0_i_5 (gr20),
        .\badr[15]_INST_0_i_5_0 (gr23),
        .\badr[15]_INST_0_i_5_1 (gr24),
        .\grn_reg[0] (\grn_reg[0]_3 ),
        .\grn_reg[0]_0 (\grn_reg[0]_4 ),
        .\grn_reg[10] (\grn_reg[10]_2 ),
        .\grn_reg[10]_0 (\grn_reg[10]_3 ),
        .\grn_reg[11] (\grn_reg[11]_2 ),
        .\grn_reg[11]_0 (\grn_reg[11]_3 ),
        .\grn_reg[12] (\grn_reg[12]_2 ),
        .\grn_reg[12]_0 (\grn_reg[12]_3 ),
        .\grn_reg[13] (\grn_reg[13]_2 ),
        .\grn_reg[13]_0 (\grn_reg[13]_3 ),
        .\grn_reg[14] (\grn_reg[14]_2 ),
        .\grn_reg[14]_0 (\grn_reg[14]_3 ),
        .\grn_reg[15] (\grn_reg[15]_5 ),
        .\grn_reg[15]_0 (\grn_reg[15]_6 ),
        .\grn_reg[1] (\grn_reg[1]_3 ),
        .\grn_reg[1]_0 (\grn_reg[1]_4 ),
        .\grn_reg[2] (\grn_reg[2]_3 ),
        .\grn_reg[2]_0 (\grn_reg[2]_4 ),
        .\grn_reg[3] (\grn_reg[3]_3 ),
        .\grn_reg[3]_0 (\grn_reg[3]_4 ),
        .\grn_reg[4] (\grn_reg[4]_3 ),
        .\grn_reg[4]_0 (\grn_reg[4]_4 ),
        .\grn_reg[5] (\grn_reg[5]_3 ),
        .\grn_reg[5]_0 (\grn_reg[5]_4 ),
        .\grn_reg[6] (\grn_reg[6]_2 ),
        .\grn_reg[6]_0 (\grn_reg[6]_3 ),
        .\grn_reg[7] (\grn_reg[7]_2 ),
        .\grn_reg[7]_0 (\grn_reg[7]_3 ),
        .\grn_reg[8] (\grn_reg[8]_2 ),
        .\grn_reg[8]_0 (\grn_reg[8]_3 ),
        .\grn_reg[9] (\grn_reg[9]_2 ),
        .\grn_reg[9]_0 (\grn_reg[9]_3 ),
        .\i_/badr[15]_INST_0_i_17_0 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/badr[15]_INST_0_i_17_1 (gr26),
        .\i_/badr[15]_INST_0_i_17_2 (gr25),
        .\i_/badr[15]_INST_0_i_17_3 (\i_/badr[15]_INST_0_i_17 ),
        .\i_/badr[15]_INST_0_i_18_0 (gr22),
        .\i_/badr[15]_INST_0_i_18_1 (gr21),
        .out(gr27));
  niho_rgf_bank_bus_4 bbuso
       (.bbus_sel_0(bbus_sel_0),
        .\bdatw[15]_INST_0_i_9 (gr03),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .\grn_reg[0] (\grn_reg[0]_1 ),
        .\grn_reg[0]_0 (\grn_reg[0]_2 ),
        .\grn_reg[10] (\grn_reg[10]_1 ),
        .\grn_reg[11] (\grn_reg[11]_1 ),
        .\grn_reg[12] (\grn_reg[12]_1 ),
        .\grn_reg[13] (\grn_reg[13]_1 ),
        .\grn_reg[14] (\grn_reg[14]_1 ),
        .\grn_reg[15] (\grn_reg[15]_4 ),
        .\grn_reg[1] (\grn_reg[1]_1 ),
        .\grn_reg[1]_0 (\grn_reg[1]_2 ),
        .\grn_reg[2] (\grn_reg[2]_1 ),
        .\grn_reg[2]_0 (\grn_reg[2]_2 ),
        .\grn_reg[3] (\grn_reg[3]_1 ),
        .\grn_reg[3]_0 (\grn_reg[3]_2 ),
        .\grn_reg[4] (\grn_reg[4]_1 ),
        .\grn_reg[4]_0 (\grn_reg[4]_2 ),
        .\grn_reg[5] (\grn_reg[5]_1 ),
        .\grn_reg[5]_0 (\grn_reg[5]_2 ),
        .\grn_reg[6] (\grn_reg[6]_1 ),
        .\grn_reg[7] (\grn_reg[7]_1 ),
        .\grn_reg[8] (\grn_reg[8]_1 ),
        .\grn_reg[9] (\grn_reg[9]_1 ),
        .\i_/bdatw[15]_INST_0_i_26_0 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/bdatw[15]_INST_0_i_26_1 (gr07),
        .\i_/bdatw[15]_INST_0_i_26_2 (gr00),
        .\i_/bdatw[15]_INST_0_i_26_3 (gr02),
        .\i_/bdatw[15]_INST_0_i_26_4 (gr01),
        .\i_/bdatw[15]_INST_0_i_50_0 (gr06),
        .\i_/bdatw[15]_INST_0_i_50_1 (gr05),
        .\i_/bdatw[15]_INST_0_i_66_0 (\i_/badr[15]_INST_0_i_19 ),
        .\i_/bdatw[15]_INST_0_i_66_1 (\i_/bdatw[15]_INST_0_i_66 ),
        .\i_/bdatw[15]_INST_0_i_66_2 (\i_/bdatw[15]_INST_0_i_66_0 ),
        .\i_/bdatw[15]_INST_0_i_66_3 (\i_/bdatw[15]_INST_0_i_66_1 ),
        .\i_/bdatw[15]_INST_0_i_66_4 (\i_/bdatw[15]_INST_0_i_66_2 ),
        .out(gr04));
  niho_rgf_bank_bus_5 bbuso2h
       (.bbus_sel_0({bbus_sel_0[5:3],bbus_sel_0[0]}),
        .\bdatw[16]_INST_0_i_3 (\bdatw[16]_INST_0_i_3 ),
        .\bdatw[16]_INST_0_i_3_0 (\bdatw[16]_INST_0_i_3_0 ),
        .\bdatw[17]_INST_0_i_3 (\bdatw[17]_INST_0_i_3 ),
        .\bdatw[17]_INST_0_i_3_0 (\bdatw[17]_INST_0_i_3_0 ),
        .\bdatw[18]_INST_0_i_3 (\bdatw[18]_INST_0_i_3 ),
        .\bdatw[18]_INST_0_i_3_0 (\bdatw[18]_INST_0_i_3_0 ),
        .\bdatw[19]_INST_0_i_3 (\bdatw[19]_INST_0_i_3 ),
        .\bdatw[19]_INST_0_i_3_0 (\bdatw[19]_INST_0_i_3_0 ),
        .\bdatw[20]_INST_0_i_3 (\bdatw[20]_INST_0_i_3 ),
        .\bdatw[20]_INST_0_i_3_0 (\bdatw[20]_INST_0_i_3_0 ),
        .\bdatw[21]_INST_0_i_3 (\bdatw[21]_INST_0_i_3 ),
        .\bdatw[21]_INST_0_i_3_0 (\bdatw[21]_INST_0_i_3_0 ),
        .\bdatw[22]_INST_0_i_3 (\bdatw[22]_INST_0_i_3 ),
        .\bdatw[22]_INST_0_i_3_0 (\bdatw[22]_INST_0_i_3_0 ),
        .\bdatw[23]_INST_0_i_3 (\bdatw[23]_INST_0_i_3 ),
        .\bdatw[23]_INST_0_i_3_0 (\bdatw[23]_INST_0_i_3_0 ),
        .\bdatw[24]_INST_0_i_3 (\bdatw[24]_INST_0_i_3 ),
        .\bdatw[24]_INST_0_i_3_0 (\bdatw[24]_INST_0_i_3_0 ),
        .\bdatw[25]_INST_0_i_3 (\bdatw[25]_INST_0_i_3 ),
        .\bdatw[25]_INST_0_i_3_0 (\bdatw[25]_INST_0_i_3_0 ),
        .\bdatw[26]_INST_0_i_3 (\bdatw[26]_INST_0_i_3 ),
        .\bdatw[26]_INST_0_i_3_0 (\bdatw[26]_INST_0_i_3_0 ),
        .\bdatw[27]_INST_0_i_3 (\bdatw[27]_INST_0_i_3 ),
        .\bdatw[27]_INST_0_i_3_0 (\bdatw[27]_INST_0_i_3_0 ),
        .\bdatw[28]_INST_0_i_3 (\bdatw[28]_INST_0_i_3 ),
        .\bdatw[28]_INST_0_i_3_0 (\bdatw[28]_INST_0_i_3_0 ),
        .\bdatw[29]_INST_0_i_3 (\bdatw[29]_INST_0_i_3 ),
        .\bdatw[29]_INST_0_i_3_0 (\bdatw[29]_INST_0_i_3_0 ),
        .\bdatw[30]_INST_0_i_3 (\bdatw[30]_INST_0_i_3 ),
        .\bdatw[30]_INST_0_i_3_0 (\bdatw[30]_INST_0_i_3_0 ),
        .\bdatw[31]_INST_0_i_5 (gr20),
        .\bdatw[31]_INST_0_i_5_0 (\bdatw[31]_INST_0_i_5 ),
        .\bdatw[31]_INST_0_i_5_1 (gr23),
        .\bdatw[31]_INST_0_i_5_2 (gr24),
        .\bdatw[31]_INST_0_i_5_3 (\bdatw[31]_INST_0_i_5_0 ),
        .\grn_reg[0] (\grn_reg[0]_9 ),
        .\grn_reg[0]_0 (\grn_reg[0]_10 ),
        .\grn_reg[10] (\grn_reg[10]_7 ),
        .\grn_reg[10]_0 (\grn_reg[10]_8 ),
        .\grn_reg[11] (\grn_reg[11]_7 ),
        .\grn_reg[11]_0 (\grn_reg[11]_8 ),
        .\grn_reg[12] (\grn_reg[12]_7 ),
        .\grn_reg[12]_0 (\grn_reg[12]_8 ),
        .\grn_reg[13] (\grn_reg[13]_7 ),
        .\grn_reg[13]_0 (\grn_reg[13]_8 ),
        .\grn_reg[14] (\grn_reg[14]_7 ),
        .\grn_reg[14]_0 (\grn_reg[14]_8 ),
        .\grn_reg[15] (\grn_reg[15]_10 ),
        .\grn_reg[15]_0 (\grn_reg[15]_11 ),
        .\grn_reg[1] (\grn_reg[1]_9 ),
        .\grn_reg[1]_0 (\grn_reg[1]_10 ),
        .\grn_reg[2] (\grn_reg[2]_9 ),
        .\grn_reg[2]_0 (\grn_reg[2]_10 ),
        .\grn_reg[3] (\grn_reg[3]_9 ),
        .\grn_reg[3]_0 (\grn_reg[3]_10 ),
        .\grn_reg[4] (\grn_reg[4]_9 ),
        .\grn_reg[4]_0 (\grn_reg[4]_10 ),
        .\grn_reg[5] (\grn_reg[5]_9 ),
        .\grn_reg[5]_0 (\grn_reg[5]_10 ),
        .\grn_reg[6] (\grn_reg[6]_7 ),
        .\grn_reg[6]_0 (\grn_reg[6]_8 ),
        .\grn_reg[7] (\grn_reg[7]_7 ),
        .\grn_reg[7]_0 (\grn_reg[7]_8 ),
        .\grn_reg[8] (\grn_reg[8]_7 ),
        .\grn_reg[8]_0 (\grn_reg[8]_8 ),
        .\grn_reg[9] (\grn_reg[9]_7 ),
        .\grn_reg[9]_0 (\grn_reg[9]_8 ),
        .\i_/bdatw[31]_INST_0_i_17_0 ({\i_/badr[15]_INST_0_i_20 [2],\i_/badr[15]_INST_0_i_20 [0]}),
        .out(gr27));
  niho_rgf_bank_bus_6 bbuso2l
       (.bbus_sel_0(bbus_sel_0[2:1]),
        .\bdatw[15]_INST_0_i_9 (gr27),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .\grn_reg[0] (\grn_reg[0]_5 ),
        .\grn_reg[0]_0 (\grn_reg[0]_6 ),
        .\grn_reg[10] (\grn_reg[10]_4 ),
        .\grn_reg[11] (\grn_reg[11]_4 ),
        .\grn_reg[12] (\grn_reg[12]_4 ),
        .\grn_reg[13] (\grn_reg[13]_4 ),
        .\grn_reg[14] (\grn_reg[14]_4 ),
        .\grn_reg[15] (\grn_reg[15]_7 ),
        .\grn_reg[1] (\grn_reg[1]_5 ),
        .\grn_reg[1]_0 (\grn_reg[1]_6 ),
        .\grn_reg[2] (\grn_reg[2]_5 ),
        .\grn_reg[2]_0 (\grn_reg[2]_6 ),
        .\grn_reg[3] (\grn_reg[3]_5 ),
        .\grn_reg[3]_0 (\grn_reg[3]_6 ),
        .\grn_reg[4] (\grn_reg[4]_5 ),
        .\grn_reg[4]_0 (\grn_reg[4]_6 ),
        .\grn_reg[5] (\grn_reg[5]_5 ),
        .\grn_reg[5]_0 (\grn_reg[5]_6 ),
        .\grn_reg[6] (\grn_reg[6]_4 ),
        .\grn_reg[7] (\grn_reg[7]_4 ),
        .\grn_reg[8] (\grn_reg[8]_4 ),
        .\grn_reg[9] (\grn_reg[9]_4 ),
        .\i_/bdatw[15]_INST_0_i_27_0 (\i_/badr[15]_INST_0_i_17 ),
        .\i_/bdatw[15]_INST_0_i_27_1 (\i_/bdatw[15]_INST_0_i_66_0 ),
        .\i_/bdatw[15]_INST_0_i_27_2 (\i_/bdatw[15]_INST_0_i_66_1 ),
        .\i_/bdatw[15]_INST_0_i_27_3 (\i_/bdatw[15]_INST_0_i_27 ),
        .\i_/bdatw[15]_INST_0_i_27_4 (gr26),
        .\i_/bdatw[15]_INST_0_i_27_5 (gr25),
        .\i_/bdatw[15]_INST_0_i_27_6 (gr21),
        .\i_/bdatw[15]_INST_0_i_27_7 (gr22),
        .\i_/bdatw[15]_INST_0_i_27_8 (\i_/bdatw[15]_INST_0_i_27_0 ),
        .\i_/bdatw[15]_INST_0_i_52_0 (\i_/bdatw[15]_INST_0_i_66 ),
        .\i_/bdatw[15]_INST_0_i_52_1 (\i_/bdatw[15]_INST_0_i_66_2 ),
        .\i_/bdatw[15]_INST_0_i_53_0 (gr24),
        .\i_/bdatw[15]_INST_0_i_53_1 (gr23),
        .\i_/bdatw[15]_INST_0_i_53_2 (\i_/badr[15]_INST_0_i_20 ),
        .\i_/bdatw[15]_INST_0_i_67_0 (\i_/bdatw[15]_INST_0_i_67 ),
        .\i_/bdatw[15]_INST_0_i_67_1 (\i_/bdatw[15]_INST_0_i_67_0 ),
        .out(gr20));
  niho_rgf_grn grn00
       (.Q(gr00),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_12 ));
  niho_rgf_grn_7 grn01
       (.Q(gr01),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_13 ));
  niho_rgf_grn_8 grn02
       (.Q(gr02),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_14 ));
  niho_rgf_grn_9 grn03
       (.E(E),
        .Q(gr03),
        .SR(SR),
        .cbus(cbus),
        .clk(clk));
  niho_rgf_grn_10 grn04
       (.Q(gr04),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_15 ));
  niho_rgf_grn_11 grn05
       (.Q(gr05),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_11 ));
  niho_rgf_grn_12 grn06
       (.Q(gr06),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_16 ));
  niho_rgf_grn_13 grn07
       (.Q(gr07),
        .SR(SR),
        .cbus(cbus),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_17 ));
  niho_rgf_grn_14 grn20
       (.Q(gr20),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_18 ),
        .\grn_reg[15]_1 (\grn_reg[15]_19 ));
  niho_rgf_grn_15 grn21
       (.Q(gr21),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_20 ),
        .\grn_reg[15]_1 (\grn_reg[15]_19 ));
  niho_rgf_grn_16 grn22
       (.Q(gr22),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_21 ),
        .\grn_reg[15]_1 (\grn_reg[15]_19 ));
  niho_rgf_grn_17 grn23
       (.Q(gr23),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_12 ),
        .\grn_reg[15]_0 (\grn_reg[15]_19 ));
  niho_rgf_grn_18 grn24
       (.Q(gr24),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_22 ),
        .\grn_reg[15]_1 (\grn_reg[15]_19 ));
  niho_rgf_grn_19 grn25
       (.Q(gr25),
        .SR(SR),
        .clk(clk),
        .\grn_reg[0]_0 (\grn_reg[0]_13 ),
        .\grn_reg[15]_0 (\grn_reg[15]_19 ));
  niho_rgf_grn_20 grn26
       (.Q(gr26),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_23 ),
        .\grn_reg[15]_1 (\grn_reg[15]_19 ));
  niho_rgf_grn_21 grn27
       (.Q(gr27),
        .SR(SR),
        .clk(clk),
        .\grn_reg[15]_0 (\grn_reg[15]_24 ),
        .\grn_reg[15]_1 (\grn_reg[15]_19 ),
        .rst_n(rst_n));
endmodule

module niho_rgf_bank_bus
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[15]_INST_0_i_5 ,
    \i_/badr[15]_INST_0_i_20_0 ,
    abus_sel_0,
    \badr[15]_INST_0_i_5_0 ,
    \badr[15]_INST_0_i_5_1 ,
    \i_/badr[15]_INST_0_i_19_0 ,
    \i_/badr[15]_INST_0_i_19_1 ,
    \i_/badr[15]_INST_0_i_19_2 ,
    \i_/badr[15]_INST_0_i_20_1 ,
    \i_/badr[15]_INST_0_i_20_2 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_5 ;
  input [2:0]\i_/badr[15]_INST_0_i_20_0 ;
  input [7:0]abus_sel_0;
  input [15:0]\badr[15]_INST_0_i_5_0 ;
  input [15:0]\badr[15]_INST_0_i_5_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_19_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_19_1 ;
  input \i_/badr[15]_INST_0_i_19_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_20_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_20_2 ;

  wire [7:0]abus_sel_0;
  wire [15:0]\badr[15]_INST_0_i_5 ;
  wire [15:0]\badr[15]_INST_0_i_5_0 ;
  wire [15:0]\badr[15]_INST_0_i_5_1 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_19_n_0 ;
  wire \i_/badr[0]_INST_0_i_20_n_0 ;
  wire \i_/badr[10]_INST_0_i_19_n_0 ;
  wire \i_/badr[10]_INST_0_i_20_n_0 ;
  wire \i_/badr[11]_INST_0_i_19_n_0 ;
  wire \i_/badr[11]_INST_0_i_20_n_0 ;
  wire \i_/badr[12]_INST_0_i_20_n_0 ;
  wire \i_/badr[12]_INST_0_i_21_n_0 ;
  wire \i_/badr[13]_INST_0_i_19_n_0 ;
  wire \i_/badr[13]_INST_0_i_20_n_0 ;
  wire \i_/badr[14]_INST_0_i_19_n_0 ;
  wire \i_/badr[14]_INST_0_i_20_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_19_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_19_1 ;
  wire \i_/badr[15]_INST_0_i_19_2 ;
  wire [2:0]\i_/badr[15]_INST_0_i_20_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_20_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_20_2 ;
  wire \i_/badr[15]_INST_0_i_40_n_0 ;
  wire \i_/badr[15]_INST_0_i_43_n_0 ;
  wire \i_/badr[1]_INST_0_i_19_n_0 ;
  wire \i_/badr[1]_INST_0_i_20_n_0 ;
  wire \i_/badr[2]_INST_0_i_19_n_0 ;
  wire \i_/badr[2]_INST_0_i_20_n_0 ;
  wire \i_/badr[3]_INST_0_i_19_n_0 ;
  wire \i_/badr[3]_INST_0_i_20_n_0 ;
  wire \i_/badr[4]_INST_0_i_20_n_0 ;
  wire \i_/badr[4]_INST_0_i_21_n_0 ;
  wire \i_/badr[5]_INST_0_i_19_n_0 ;
  wire \i_/badr[5]_INST_0_i_20_n_0 ;
  wire \i_/badr[6]_INST_0_i_19_n_0 ;
  wire \i_/badr[6]_INST_0_i_20_n_0 ;
  wire \i_/badr[7]_INST_0_i_19_n_0 ;
  wire \i_/badr[7]_INST_0_i_20_n_0 ;
  wire \i_/badr[8]_INST_0_i_20_n_0 ;
  wire \i_/badr[8]_INST_0_i_21_n_0 ;
  wire \i_/badr[9]_INST_0_i_19_n_0 ;
  wire \i_/badr[9]_INST_0_i_20_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [0]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_19_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[0]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [0]),
        .I4(\i_/badr[0]_INST_0_i_20_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[0]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [0]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [0]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[0]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[0]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [0]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [0]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[0]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [10]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_19_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[10]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [10]),
        .I4(\i_/badr[10]_INST_0_i_20_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[10]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [10]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [10]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[10]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[10]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [10]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [10]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[10]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [11]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_19_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[11]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [11]),
        .I4(\i_/badr[11]_INST_0_i_20_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[11]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [11]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [11]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[11]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[11]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [11]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [11]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[11]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [12]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_20_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[12]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [12]),
        .I4(\i_/badr[12]_INST_0_i_21_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[12]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [12]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [12]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[12]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[12]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [12]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [12]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[12]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [13]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_19_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[13]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [13]),
        .I4(\i_/badr[13]_INST_0_i_20_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[13]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [13]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [13]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[13]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[13]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [13]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [13]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[13]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [14]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_19_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[14]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [14]),
        .I4(\i_/badr[14]_INST_0_i_20_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[14]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [14]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [14]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[14]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[14]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [14]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [14]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[14]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [15]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_40_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(out[15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [15]),
        .I4(\i_/badr[15]_INST_0_i_43_n_0 ),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/badr[15]_INST_0_i_38 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I3(abus_sel_0[7]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/badr[15]_INST_0_i_39 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I3(abus_sel_0[0]),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[15]_INST_0_i_40 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [15]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [15]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[15]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/badr[15]_INST_0_i_41 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I3(abus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/badr[15]_INST_0_i_42 
       (.I0(\i_/badr[15]_INST_0_i_20_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_20_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_20_0 [0]),
        .I3(abus_sel_0[4]),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[15]_INST_0_i_43 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [15]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [15]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[15]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [1]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_19_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[1]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [1]),
        .I4(\i_/badr[1]_INST_0_i_20_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[1]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [1]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [1]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[1]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[1]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [1]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [1]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[1]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [2]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_19_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[2]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [2]),
        .I4(\i_/badr[2]_INST_0_i_20_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[2]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [2]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [2]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[2]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[2]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [2]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [2]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[2]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [3]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_19_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[3]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [3]),
        .I4(\i_/badr[3]_INST_0_i_20_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[3]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [3]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [3]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[3]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[3]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [3]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [3]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[3]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [4]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_20_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[4]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [4]),
        .I4(\i_/badr[4]_INST_0_i_21_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[4]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [4]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [4]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[4]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[4]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [4]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [4]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[4]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [5]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_19_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[5]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [5]),
        .I4(\i_/badr[5]_INST_0_i_20_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[5]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [5]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [5]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[5]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[5]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [5]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [5]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[5]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [6]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_19_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[6]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [6]),
        .I4(\i_/badr[6]_INST_0_i_20_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[6]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [6]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [6]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[6]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[6]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [6]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [6]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[6]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [7]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_19_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[7]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [7]),
        .I4(\i_/badr[7]_INST_0_i_20_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[7]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [7]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [7]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[7]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[7]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [7]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [7]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[7]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [8]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_20_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[8]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [8]),
        .I4(\i_/badr[8]_INST_0_i_21_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[8]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [8]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [8]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[8]_INST_0_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[8]_INST_0_i_21 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [8]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [8]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[8]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [9]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_19_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(out[9]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5 [9]),
        .I4(\i_/badr[9]_INST_0_i_20_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[9]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_19_0 [9]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_19_1 [9]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[9]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[9]_INST_0_i_20 
       (.I0(\i_/badr[15]_INST_0_i_20_1 [9]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_20_2 [9]),
        .I3(\i_/badr[15]_INST_0_i_19_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[9]_INST_0_i_20_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_2
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[31]_INST_0_i_1 ,
    \badr[31]_INST_0_i_1_0 ,
    \badr[30]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1 ,
    \badr[31]_INST_0_i_1_1 ,
    \badr[31]_INST_0_i_1_2 ,
    \badr[31]_INST_0_i_1_3 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1_0 ,
    \i_/badr[31]_INST_0_i_7_0 ,
    abus_sel_0);
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[31]_INST_0_i_1 ;
  input \badr[31]_INST_0_i_1_0 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1 ;
  input [15:0]\badr[31]_INST_0_i_1_1 ;
  input [15:0]\badr[31]_INST_0_i_1_2 ;
  input \badr[31]_INST_0_i_1_3 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1_0 ;
  input [1:0]\i_/badr[31]_INST_0_i_7_0 ;
  input [3:0]abus_sel_0;

  wire [3:0]abus_sel_0;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire [15:0]\badr[31]_INST_0_i_1 ;
  wire \badr[31]_INST_0_i_1_0 ;
  wire [15:0]\badr[31]_INST_0_i_1_1 ;
  wire [15:0]\badr[31]_INST_0_i_1_2 ;
  wire \badr[31]_INST_0_i_1_3 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire [1:0]\i_/badr[31]_INST_0_i_7_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[16]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [0]),
        .I4(\badr[16]_INST_0_i_1 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[16]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [0]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [0]),
        .I4(\badr[16]_INST_0_i_1_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[17]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [1]),
        .I4(\badr[17]_INST_0_i_1 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[17]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [1]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [1]),
        .I4(\badr[17]_INST_0_i_1_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[18]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [2]),
        .I4(\badr[18]_INST_0_i_1 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[18]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [2]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [2]),
        .I4(\badr[18]_INST_0_i_1_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[19]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [3]),
        .I4(\badr[19]_INST_0_i_1 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[19]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [3]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [3]),
        .I4(\badr[19]_INST_0_i_1_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[20]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [4]),
        .I4(\badr[20]_INST_0_i_1 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[20]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [4]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [4]),
        .I4(\badr[20]_INST_0_i_1_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[21]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [5]),
        .I4(\badr[21]_INST_0_i_1 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[21]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [5]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [5]),
        .I4(\badr[21]_INST_0_i_1_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[22]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [6]),
        .I4(\badr[22]_INST_0_i_1 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[22]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [6]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [6]),
        .I4(\badr[22]_INST_0_i_1_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[23]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [7]),
        .I4(\badr[23]_INST_0_i_1 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[23]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [7]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [7]),
        .I4(\badr[23]_INST_0_i_1_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[24]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [8]),
        .I4(\badr[24]_INST_0_i_1 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[24]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [8]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [8]),
        .I4(\badr[24]_INST_0_i_1_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[25]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [9]),
        .I4(\badr[25]_INST_0_i_1 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[25]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [9]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [9]),
        .I4(\badr[25]_INST_0_i_1_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[26]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [10]),
        .I4(\badr[26]_INST_0_i_1 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[26]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [10]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [10]),
        .I4(\badr[26]_INST_0_i_1_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[27]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [11]),
        .I4(\badr[27]_INST_0_i_1 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[27]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [11]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [11]),
        .I4(\badr[27]_INST_0_i_1_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[28]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [12]),
        .I4(\badr[28]_INST_0_i_1 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[28]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [12]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [12]),
        .I4(\badr[28]_INST_0_i_1_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[29]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [13]),
        .I4(\badr[29]_INST_0_i_1 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[29]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [13]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [13]),
        .I4(\badr[29]_INST_0_i_1_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[30]_INST_0_i_5 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [14]),
        .I4(\badr[30]_INST_0_i_1 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[30]_INST_0_i_6 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [14]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [14]),
        .I4(\badr[30]_INST_0_i_1_0 ),
        .O(\grn_reg[14]_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[31]_INST_0_i_20 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_7_0 [1]),
        .I2(abus_sel_0[3]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[31]_INST_0_i_21 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_7_0 [1]),
        .I2(abus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[31]_INST_0_i_23 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_7_0 [1]),
        .I2(abus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/badr[31]_INST_0_i_24 
       (.I0(\i_/badr[31]_INST_0_i_7_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_7_0 [1]),
        .I2(abus_sel_0[2]),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[31]_INST_0_i_6 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [15]),
        .I4(\badr[31]_INST_0_i_1_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[31]_INST_0_i_7 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [15]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [15]),
        .I4(\badr[31]_INST_0_i_1_3 ),
        .O(\grn_reg[15]_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_22
   (p_1_in,
    out,
    \mul_a_reg[15] ,
    \i_/badr[15]_INST_0_i_3_0 ,
    \i_/badr[15]_INST_0_i_3_1 ,
    \i_/badr[15]_INST_0_i_10_0 ,
    abus_sel_0,
    \i_/badr[15]_INST_0_i_3_2 ,
    \i_/badr[15]_INST_0_i_3_3 ,
    \i_/badr[15]_INST_0_i_11_0 ,
    \i_/badr[15]_INST_0_i_11_1 ,
    bank_sel);
  output [15:0]p_1_in;
  input [15:0]out;
  input [15:0]\mul_a_reg[15] ;
  input [15:0]\i_/badr[15]_INST_0_i_3_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_3_1 ;
  input [2:0]\i_/badr[15]_INST_0_i_10_0 ;
  input [7:0]abus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_3_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_3_3 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_11_1 ;
  input [0:0]bank_sel;

  wire [7:0]abus_sel_0;
  wire [0:0]bank_sel;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \i_/badr[0]_INST_0_i_15_n_0 ;
  wire \i_/badr[0]_INST_0_i_7_n_0 ;
  wire \i_/badr[0]_INST_0_i_8_n_0 ;
  wire \i_/badr[10]_INST_0_i_15_n_0 ;
  wire \i_/badr[10]_INST_0_i_7_n_0 ;
  wire \i_/badr[10]_INST_0_i_8_n_0 ;
  wire \i_/badr[11]_INST_0_i_15_n_0 ;
  wire \i_/badr[11]_INST_0_i_7_n_0 ;
  wire \i_/badr[11]_INST_0_i_8_n_0 ;
  wire \i_/badr[12]_INST_0_i_16_n_0 ;
  wire \i_/badr[12]_INST_0_i_7_n_0 ;
  wire \i_/badr[12]_INST_0_i_8_n_0 ;
  wire \i_/badr[13]_INST_0_i_15_n_0 ;
  wire \i_/badr[13]_INST_0_i_7_n_0 ;
  wire \i_/badr[13]_INST_0_i_8_n_0 ;
  wire \i_/badr[14]_INST_0_i_15_n_0 ;
  wire \i_/badr[14]_INST_0_i_7_n_0 ;
  wire \i_/badr[14]_INST_0_i_8_n_0 ;
  wire [2:0]\i_/badr[15]_INST_0_i_10_0 ;
  wire \i_/badr[15]_INST_0_i_10_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_11_1 ;
  wire \i_/badr[15]_INST_0_i_11_n_0 ;
  wire \i_/badr[15]_INST_0_i_26_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_3_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_3_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_3_2 ;
  wire [15:0]\i_/badr[15]_INST_0_i_3_3 ;
  wire \i_/badr[1]_INST_0_i_15_n_0 ;
  wire \i_/badr[1]_INST_0_i_7_n_0 ;
  wire \i_/badr[1]_INST_0_i_8_n_0 ;
  wire \i_/badr[2]_INST_0_i_15_n_0 ;
  wire \i_/badr[2]_INST_0_i_7_n_0 ;
  wire \i_/badr[2]_INST_0_i_8_n_0 ;
  wire \i_/badr[3]_INST_0_i_15_n_0 ;
  wire \i_/badr[3]_INST_0_i_7_n_0 ;
  wire \i_/badr[3]_INST_0_i_8_n_0 ;
  wire \i_/badr[4]_INST_0_i_16_n_0 ;
  wire \i_/badr[4]_INST_0_i_7_n_0 ;
  wire \i_/badr[4]_INST_0_i_8_n_0 ;
  wire \i_/badr[5]_INST_0_i_15_n_0 ;
  wire \i_/badr[5]_INST_0_i_7_n_0 ;
  wire \i_/badr[5]_INST_0_i_8_n_0 ;
  wire \i_/badr[6]_INST_0_i_15_n_0 ;
  wire \i_/badr[6]_INST_0_i_7_n_0 ;
  wire \i_/badr[6]_INST_0_i_8_n_0 ;
  wire \i_/badr[7]_INST_0_i_15_n_0 ;
  wire \i_/badr[7]_INST_0_i_7_n_0 ;
  wire \i_/badr[7]_INST_0_i_8_n_0 ;
  wire \i_/badr[8]_INST_0_i_16_n_0 ;
  wire \i_/badr[8]_INST_0_i_7_n_0 ;
  wire \i_/badr[8]_INST_0_i_8_n_0 ;
  wire \i_/badr[9]_INST_0_i_15_n_0 ;
  wire \i_/badr[9]_INST_0_i_7_n_0 ;
  wire \i_/badr[9]_INST_0_i_8_n_0 ;
  wire [15:0]\mul_a_reg[15] ;
  wire [15:0]out;
  wire [15:0]p_1_in;

  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[0]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [0]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [0]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[0]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_3 
       (.I0(out[0]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [0]),
        .I3(gr5_bus1),
        .I4(\i_/badr[0]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[0]_INST_0_i_8_n_0 ),
        .O(p_1_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [0]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [0]),
        .I4(\i_/badr[0]_INST_0_i_15_n_0 ),
        .O(\i_/badr[0]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[10]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [10]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [10]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[10]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_3 
       (.I0(out[10]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [10]),
        .I3(gr5_bus1),
        .I4(\i_/badr[10]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[10]_INST_0_i_8_n_0 ),
        .O(p_1_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [10]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [10]),
        .I4(\i_/badr[10]_INST_0_i_15_n_0 ),
        .O(\i_/badr[10]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[11]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [11]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [11]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[11]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_3 
       (.I0(out[11]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [11]),
        .I3(gr5_bus1),
        .I4(\i_/badr[11]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[11]_INST_0_i_8_n_0 ),
        .O(p_1_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [11]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [11]),
        .I4(\i_/badr[11]_INST_0_i_15_n_0 ),
        .O(\i_/badr[11]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[12]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [12]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [12]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[12]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_3 
       (.I0(out[12]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [12]),
        .I3(gr5_bus1),
        .I4(\i_/badr[12]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[12]_INST_0_i_8_n_0 ),
        .O(p_1_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [12]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [12]),
        .I4(\i_/badr[12]_INST_0_i_16_n_0 ),
        .O(\i_/badr[12]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[13]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [13]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [13]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[13]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_3 
       (.I0(out[13]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [13]),
        .I3(gr5_bus1),
        .I4(\i_/badr[13]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[13]_INST_0_i_8_n_0 ),
        .O(p_1_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [13]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [13]),
        .I4(\i_/badr[13]_INST_0_i_15_n_0 ),
        .O(\i_/badr[13]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[14]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [14]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [14]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[14]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_3 
       (.I0(out[14]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [14]),
        .I3(gr5_bus1),
        .I4(\i_/badr[14]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[14]_INST_0_i_8_n_0 ),
        .O(p_1_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [14]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [14]),
        .I4(\i_/badr[14]_INST_0_i_15_n_0 ),
        .O(\i_/badr[14]_INST_0_i_8_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_10 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [15]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [15]),
        .I4(\i_/badr[15]_INST_0_i_26_n_0 ),
        .O(\i_/badr[15]_INST_0_i_11_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/badr[15]_INST_0_i_22 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(abus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/badr[15]_INST_0_i_23 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(abus_sel_0[7]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/badr[15]_INST_0_i_24 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(abus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/badr[15]_INST_0_i_25 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(abus_sel_0[4]),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[15]_INST_0_i_26 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [15]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [15]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[15]_INST_0_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_3 
       (.I0(out[15]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [15]),
        .I3(gr5_bus1),
        .I4(\i_/badr[15]_INST_0_i_10_n_0 ),
        .I5(\i_/badr[15]_INST_0_i_11_n_0 ),
        .O(p_1_in[15]));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/badr[15]_INST_0_i_8 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(abus_sel_0[6]),
        .O(gr6_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/badr[15]_INST_0_i_9 
       (.I0(\i_/badr[15]_INST_0_i_10_0 [1]),
        .I1(\i_/badr[15]_INST_0_i_10_0 [2]),
        .I2(\i_/badr[15]_INST_0_i_10_0 [0]),
        .I3(abus_sel_0[5]),
        .O(gr5_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[1]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [1]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [1]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[1]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_3 
       (.I0(out[1]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [1]),
        .I3(gr5_bus1),
        .I4(\i_/badr[1]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[1]_INST_0_i_8_n_0 ),
        .O(p_1_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [1]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [1]),
        .I4(\i_/badr[1]_INST_0_i_15_n_0 ),
        .O(\i_/badr[1]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[2]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [2]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [2]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[2]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_3 
       (.I0(out[2]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [2]),
        .I3(gr5_bus1),
        .I4(\i_/badr[2]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[2]_INST_0_i_8_n_0 ),
        .O(p_1_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [2]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [2]),
        .I4(\i_/badr[2]_INST_0_i_15_n_0 ),
        .O(\i_/badr[2]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[3]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [3]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [3]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[3]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_3 
       (.I0(out[3]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [3]),
        .I3(gr5_bus1),
        .I4(\i_/badr[3]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[3]_INST_0_i_8_n_0 ),
        .O(p_1_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [3]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [3]),
        .I4(\i_/badr[3]_INST_0_i_15_n_0 ),
        .O(\i_/badr[3]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[4]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [4]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [4]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[4]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_3 
       (.I0(out[4]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [4]),
        .I3(gr5_bus1),
        .I4(\i_/badr[4]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[4]_INST_0_i_8_n_0 ),
        .O(p_1_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [4]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [4]),
        .I4(\i_/badr[4]_INST_0_i_16_n_0 ),
        .O(\i_/badr[4]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[5]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [5]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [5]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[5]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_3 
       (.I0(out[5]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [5]),
        .I3(gr5_bus1),
        .I4(\i_/badr[5]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[5]_INST_0_i_8_n_0 ),
        .O(p_1_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [5]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [5]),
        .I4(\i_/badr[5]_INST_0_i_15_n_0 ),
        .O(\i_/badr[5]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[6]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [6]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [6]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[6]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_3 
       (.I0(out[6]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [6]),
        .I3(gr5_bus1),
        .I4(\i_/badr[6]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[6]_INST_0_i_8_n_0 ),
        .O(p_1_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [6]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [6]),
        .I4(\i_/badr[6]_INST_0_i_15_n_0 ),
        .O(\i_/badr[6]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[7]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [7]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [7]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[7]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_3 
       (.I0(out[7]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [7]),
        .I3(gr5_bus1),
        .I4(\i_/badr[7]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[7]_INST_0_i_8_n_0 ),
        .O(p_1_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [7]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [7]),
        .I4(\i_/badr[7]_INST_0_i_15_n_0 ),
        .O(\i_/badr[7]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[8]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [8]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [8]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[8]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_3 
       (.I0(out[8]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [8]),
        .I3(gr5_bus1),
        .I4(\i_/badr[8]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[8]_INST_0_i_8_n_0 ),
        .O(p_1_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [8]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [8]),
        .I4(\i_/badr[8]_INST_0_i_16_n_0 ),
        .O(\i_/badr[8]_INST_0_i_8_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[9]_INST_0_i_15 
       (.I0(\i_/badr[15]_INST_0_i_11_0 [9]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_11_1 [9]),
        .I3(bank_sel),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[9]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_3 
       (.I0(out[9]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15] [9]),
        .I3(gr5_bus1),
        .I4(\i_/badr[9]_INST_0_i_7_n_0 ),
        .I5(\i_/badr[9]_INST_0_i_8_n_0 ),
        .O(p_1_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_7 
       (.I0(\i_/badr[15]_INST_0_i_3_0 [9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_3_1 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_7_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_3_2 [9]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_3_3 [9]),
        .I4(\i_/badr[9]_INST_0_i_15_n_0 ),
        .O(\i_/badr[9]_INST_0_i_8_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_23
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[31]_INST_0_i_1 ,
    \badr[31]_INST_0_i_1_0 ,
    \badr[30]_INST_0_i_1 ,
    \badr[29]_INST_0_i_1 ,
    \badr[28]_INST_0_i_1 ,
    \badr[27]_INST_0_i_1 ,
    \badr[26]_INST_0_i_1 ,
    \badr[25]_INST_0_i_1 ,
    \badr[24]_INST_0_i_1 ,
    \badr[23]_INST_0_i_1 ,
    \badr[22]_INST_0_i_1 ,
    \badr[21]_INST_0_i_1 ,
    \badr[20]_INST_0_i_1 ,
    \badr[19]_INST_0_i_1 ,
    \badr[18]_INST_0_i_1 ,
    \badr[17]_INST_0_i_1 ,
    \badr[16]_INST_0_i_1 ,
    \badr[31]_INST_0_i_1_1 ,
    \badr[31]_INST_0_i_1_2 ,
    \badr[31]_INST_0_i_1_3 ,
    \badr[30]_INST_0_i_1_0 ,
    \badr[29]_INST_0_i_1_0 ,
    \badr[28]_INST_0_i_1_0 ,
    \badr[27]_INST_0_i_1_0 ,
    \badr[26]_INST_0_i_1_0 ,
    \badr[25]_INST_0_i_1_0 ,
    \badr[24]_INST_0_i_1_0 ,
    \badr[23]_INST_0_i_1_0 ,
    \badr[22]_INST_0_i_1_0 ,
    \badr[21]_INST_0_i_1_0 ,
    \badr[20]_INST_0_i_1_0 ,
    \badr[19]_INST_0_i_1_0 ,
    \badr[18]_INST_0_i_1_0 ,
    \badr[17]_INST_0_i_1_0 ,
    \badr[16]_INST_0_i_1_0 ,
    \i_/badr[31]_INST_0_i_5_0 ,
    abus_sel_0);
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[31]_INST_0_i_1 ;
  input \badr[31]_INST_0_i_1_0 ;
  input \badr[30]_INST_0_i_1 ;
  input \badr[29]_INST_0_i_1 ;
  input \badr[28]_INST_0_i_1 ;
  input \badr[27]_INST_0_i_1 ;
  input \badr[26]_INST_0_i_1 ;
  input \badr[25]_INST_0_i_1 ;
  input \badr[24]_INST_0_i_1 ;
  input \badr[23]_INST_0_i_1 ;
  input \badr[22]_INST_0_i_1 ;
  input \badr[21]_INST_0_i_1 ;
  input \badr[20]_INST_0_i_1 ;
  input \badr[19]_INST_0_i_1 ;
  input \badr[18]_INST_0_i_1 ;
  input \badr[17]_INST_0_i_1 ;
  input \badr[16]_INST_0_i_1 ;
  input [15:0]\badr[31]_INST_0_i_1_1 ;
  input [15:0]\badr[31]_INST_0_i_1_2 ;
  input \badr[31]_INST_0_i_1_3 ;
  input \badr[30]_INST_0_i_1_0 ;
  input \badr[29]_INST_0_i_1_0 ;
  input \badr[28]_INST_0_i_1_0 ;
  input \badr[27]_INST_0_i_1_0 ;
  input \badr[26]_INST_0_i_1_0 ;
  input \badr[25]_INST_0_i_1_0 ;
  input \badr[24]_INST_0_i_1_0 ;
  input \badr[23]_INST_0_i_1_0 ;
  input \badr[22]_INST_0_i_1_0 ;
  input \badr[21]_INST_0_i_1_0 ;
  input \badr[20]_INST_0_i_1_0 ;
  input \badr[19]_INST_0_i_1_0 ;
  input \badr[18]_INST_0_i_1_0 ;
  input \badr[17]_INST_0_i_1_0 ;
  input \badr[16]_INST_0_i_1_0 ;
  input [1:0]\i_/badr[31]_INST_0_i_5_0 ;
  input [3:0]abus_sel_0;

  wire [3:0]abus_sel_0;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[17]_INST_0_i_1_0 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1_0 ;
  wire \badr[19]_INST_0_i_1 ;
  wire \badr[19]_INST_0_i_1_0 ;
  wire \badr[20]_INST_0_i_1 ;
  wire \badr[20]_INST_0_i_1_0 ;
  wire \badr[21]_INST_0_i_1 ;
  wire \badr[21]_INST_0_i_1_0 ;
  wire \badr[22]_INST_0_i_1 ;
  wire \badr[22]_INST_0_i_1_0 ;
  wire \badr[23]_INST_0_i_1 ;
  wire \badr[23]_INST_0_i_1_0 ;
  wire \badr[24]_INST_0_i_1 ;
  wire \badr[24]_INST_0_i_1_0 ;
  wire \badr[25]_INST_0_i_1 ;
  wire \badr[25]_INST_0_i_1_0 ;
  wire \badr[26]_INST_0_i_1 ;
  wire \badr[26]_INST_0_i_1_0 ;
  wire \badr[27]_INST_0_i_1 ;
  wire \badr[27]_INST_0_i_1_0 ;
  wire \badr[28]_INST_0_i_1 ;
  wire \badr[28]_INST_0_i_1_0 ;
  wire \badr[29]_INST_0_i_1 ;
  wire \badr[29]_INST_0_i_1_0 ;
  wire \badr[30]_INST_0_i_1 ;
  wire \badr[30]_INST_0_i_1_0 ;
  wire [15:0]\badr[31]_INST_0_i_1 ;
  wire \badr[31]_INST_0_i_1_0 ;
  wire [15:0]\badr[31]_INST_0_i_1_1 ;
  wire [15:0]\badr[31]_INST_0_i_1_2 ;
  wire \badr[31]_INST_0_i_1_3 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire [1:0]\i_/badr[31]_INST_0_i_5_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[16]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [0]),
        .I4(\badr[16]_INST_0_i_1 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[16]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [0]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [0]),
        .I4(\badr[16]_INST_0_i_1_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[17]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [1]),
        .I4(\badr[17]_INST_0_i_1 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[17]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [1]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [1]),
        .I4(\badr[17]_INST_0_i_1_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[18]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [2]),
        .I4(\badr[18]_INST_0_i_1 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[18]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [2]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [2]),
        .I4(\badr[18]_INST_0_i_1_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[19]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [3]),
        .I4(\badr[19]_INST_0_i_1 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[19]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [3]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [3]),
        .I4(\badr[19]_INST_0_i_1_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[20]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [4]),
        .I4(\badr[20]_INST_0_i_1 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[20]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [4]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [4]),
        .I4(\badr[20]_INST_0_i_1_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[21]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [5]),
        .I4(\badr[21]_INST_0_i_1 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[21]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [5]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [5]),
        .I4(\badr[21]_INST_0_i_1_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[22]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [6]),
        .I4(\badr[22]_INST_0_i_1 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[22]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [6]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [6]),
        .I4(\badr[22]_INST_0_i_1_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[23]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [7]),
        .I4(\badr[23]_INST_0_i_1 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[23]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [7]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [7]),
        .I4(\badr[23]_INST_0_i_1_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[24]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [8]),
        .I4(\badr[24]_INST_0_i_1 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[24]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [8]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [8]),
        .I4(\badr[24]_INST_0_i_1_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[25]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [9]),
        .I4(\badr[25]_INST_0_i_1 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[25]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [9]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [9]),
        .I4(\badr[25]_INST_0_i_1_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[26]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [10]),
        .I4(\badr[26]_INST_0_i_1 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[26]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [10]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [10]),
        .I4(\badr[26]_INST_0_i_1_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[27]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [11]),
        .I4(\badr[27]_INST_0_i_1 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[27]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [11]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [11]),
        .I4(\badr[27]_INST_0_i_1_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[28]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [12]),
        .I4(\badr[28]_INST_0_i_1 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[28]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [12]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [12]),
        .I4(\badr[28]_INST_0_i_1_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[29]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [13]),
        .I4(\badr[29]_INST_0_i_1 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[29]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [13]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [13]),
        .I4(\badr[29]_INST_0_i_1_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[30]_INST_0_i_3 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [14]),
        .I4(\badr[30]_INST_0_i_1 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[30]_INST_0_i_4 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [14]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [14]),
        .I4(\badr[30]_INST_0_i_1_0 ),
        .O(\grn_reg[14]_0 ));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[31]_INST_0_i_14 
       (.I0(\i_/badr[31]_INST_0_i_5_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_5_0 [1]),
        .I2(abus_sel_0[3]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[31]_INST_0_i_15 
       (.I0(\i_/badr[31]_INST_0_i_5_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_5_0 [1]),
        .I2(abus_sel_0[0]),
        .O(gr0_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[31]_INST_0_i_17 
       (.I0(\i_/badr[31]_INST_0_i_5_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_5_0 [1]),
        .I2(abus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h40)) 
    \i_/badr[31]_INST_0_i_18 
       (.I0(\i_/badr[31]_INST_0_i_5_0 [0]),
        .I1(\i_/badr[31]_INST_0_i_5_0 [1]),
        .I2(abus_sel_0[2]),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[31]_INST_0_i_4 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\badr[31]_INST_0_i_1 [15]),
        .I4(\badr[31]_INST_0_i_1_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[31]_INST_0_i_5 
       (.I0(gr3_bus1),
        .I1(\badr[31]_INST_0_i_1_1 [15]),
        .I2(gr4_bus1),
        .I3(\badr[31]_INST_0_i_1_2 [15]),
        .I4(\badr[31]_INST_0_i_1_3 ),
        .O(\grn_reg[15]_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_24
   (p_0_in,
    \mul_a_reg[15] ,
    \mul_a_reg[15]_0 ,
    out,
    \i_/badr[15]_INST_0_i_4_0 ,
    \i_/badr[15]_INST_0_i_14_0 ,
    abus_sel_0,
    \i_/badr[15]_INST_0_i_4_1 ,
    \i_/badr[15]_INST_0_i_4_2 ,
    \i_/badr[15]_INST_0_i_15_0 ,
    \i_/badr[15]_INST_0_i_15_1 ,
    \i_/badr[15]_INST_0_i_15_2 );
  output [15:0]p_0_in;
  input [15:0]\mul_a_reg[15] ;
  input [15:0]\mul_a_reg[15]_0 ;
  input [15:0]out;
  input [15:0]\i_/badr[15]_INST_0_i_4_0 ;
  input [2:0]\i_/badr[15]_INST_0_i_14_0 ;
  input [7:0]abus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_4_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_4_2 ;
  input [15:0]\i_/badr[15]_INST_0_i_15_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_15_1 ;
  input \i_/badr[15]_INST_0_i_15_2 ;

  wire [7:0]abus_sel_0;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \i_/badr[0]_INST_0_i_10_n_0 ;
  wire \i_/badr[0]_INST_0_i_16_n_0 ;
  wire \i_/badr[0]_INST_0_i_9_n_0 ;
  wire \i_/badr[10]_INST_0_i_10_n_0 ;
  wire \i_/badr[10]_INST_0_i_16_n_0 ;
  wire \i_/badr[10]_INST_0_i_9_n_0 ;
  wire \i_/badr[11]_INST_0_i_10_n_0 ;
  wire \i_/badr[11]_INST_0_i_16_n_0 ;
  wire \i_/badr[11]_INST_0_i_9_n_0 ;
  wire \i_/badr[12]_INST_0_i_10_n_0 ;
  wire \i_/badr[12]_INST_0_i_17_n_0 ;
  wire \i_/badr[12]_INST_0_i_9_n_0 ;
  wire \i_/badr[13]_INST_0_i_10_n_0 ;
  wire \i_/badr[13]_INST_0_i_16_n_0 ;
  wire \i_/badr[13]_INST_0_i_9_n_0 ;
  wire \i_/badr[14]_INST_0_i_10_n_0 ;
  wire \i_/badr[14]_INST_0_i_16_n_0 ;
  wire \i_/badr[14]_INST_0_i_9_n_0 ;
  wire [2:0]\i_/badr[15]_INST_0_i_14_0 ;
  wire \i_/badr[15]_INST_0_i_14_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_15_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_15_1 ;
  wire \i_/badr[15]_INST_0_i_15_2 ;
  wire \i_/badr[15]_INST_0_i_15_n_0 ;
  wire \i_/badr[15]_INST_0_i_31_n_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_4_2 ;
  wire \i_/badr[1]_INST_0_i_10_n_0 ;
  wire \i_/badr[1]_INST_0_i_16_n_0 ;
  wire \i_/badr[1]_INST_0_i_9_n_0 ;
  wire \i_/badr[2]_INST_0_i_10_n_0 ;
  wire \i_/badr[2]_INST_0_i_16_n_0 ;
  wire \i_/badr[2]_INST_0_i_9_n_0 ;
  wire \i_/badr[3]_INST_0_i_10_n_0 ;
  wire \i_/badr[3]_INST_0_i_16_n_0 ;
  wire \i_/badr[3]_INST_0_i_9_n_0 ;
  wire \i_/badr[4]_INST_0_i_10_n_0 ;
  wire \i_/badr[4]_INST_0_i_17_n_0 ;
  wire \i_/badr[4]_INST_0_i_9_n_0 ;
  wire \i_/badr[5]_INST_0_i_10_n_0 ;
  wire \i_/badr[5]_INST_0_i_16_n_0 ;
  wire \i_/badr[5]_INST_0_i_9_n_0 ;
  wire \i_/badr[6]_INST_0_i_10_n_0 ;
  wire \i_/badr[6]_INST_0_i_16_n_0 ;
  wire \i_/badr[6]_INST_0_i_9_n_0 ;
  wire \i_/badr[7]_INST_0_i_10_n_0 ;
  wire \i_/badr[7]_INST_0_i_16_n_0 ;
  wire \i_/badr[7]_INST_0_i_9_n_0 ;
  wire \i_/badr[8]_INST_0_i_10_n_0 ;
  wire \i_/badr[8]_INST_0_i_17_n_0 ;
  wire \i_/badr[8]_INST_0_i_9_n_0 ;
  wire \i_/badr[9]_INST_0_i_10_n_0 ;
  wire \i_/badr[9]_INST_0_i_16_n_0 ;
  wire \i_/badr[9]_INST_0_i_9_n_0 ;
  wire [15:0]\mul_a_reg[15] ;
  wire [15:0]\mul_a_reg[15]_0 ;
  wire [15:0]out;
  wire [15:0]p_0_in;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [0]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [0]),
        .I4(\i_/badr[0]_INST_0_i_16_n_0 ),
        .O(\i_/badr[0]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[0]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [0]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [0]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[0]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[0]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [0]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [0]),
        .I3(gr5_bus1),
        .I4(\i_/badr[0]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[0]_INST_0_i_10_n_0 ),
        .O(p_0_in[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[0]_INST_0_i_9 
       (.I0(out[0]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [0]),
        .I3(gr7_bus1),
        .O(\i_/badr[0]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [10]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [10]),
        .I4(\i_/badr[10]_INST_0_i_16_n_0 ),
        .O(\i_/badr[10]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[10]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [10]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [10]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[10]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[10]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [10]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [10]),
        .I3(gr5_bus1),
        .I4(\i_/badr[10]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[10]_INST_0_i_10_n_0 ),
        .O(p_0_in[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[10]_INST_0_i_9 
       (.I0(out[10]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [10]),
        .I3(gr7_bus1),
        .O(\i_/badr[10]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [11]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [11]),
        .I4(\i_/badr[11]_INST_0_i_16_n_0 ),
        .O(\i_/badr[11]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[11]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [11]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [11]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[11]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[11]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [11]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [11]),
        .I3(gr5_bus1),
        .I4(\i_/badr[11]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[11]_INST_0_i_10_n_0 ),
        .O(p_0_in[11]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[11]_INST_0_i_9 
       (.I0(out[11]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [11]),
        .I3(gr7_bus1),
        .O(\i_/badr[11]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [12]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [12]),
        .I4(\i_/badr[12]_INST_0_i_17_n_0 ),
        .O(\i_/badr[12]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[12]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [12]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [12]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[12]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[12]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [12]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [12]),
        .I3(gr5_bus1),
        .I4(\i_/badr[12]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[12]_INST_0_i_10_n_0 ),
        .O(p_0_in[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[12]_INST_0_i_9 
       (.I0(out[12]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [12]),
        .I3(gr7_bus1),
        .O(\i_/badr[12]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [13]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [13]),
        .I4(\i_/badr[13]_INST_0_i_16_n_0 ),
        .O(\i_/badr[13]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[13]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [13]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [13]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[13]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[13]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [13]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [13]),
        .I3(gr5_bus1),
        .I4(\i_/badr[13]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[13]_INST_0_i_10_n_0 ),
        .O(p_0_in[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[13]_INST_0_i_9 
       (.I0(out[13]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [13]),
        .I3(gr7_bus1),
        .O(\i_/badr[13]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [14]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [14]),
        .I4(\i_/badr[14]_INST_0_i_16_n_0 ),
        .O(\i_/badr[14]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[14]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [14]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [14]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[14]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[14]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [14]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [14]),
        .I3(gr5_bus1),
        .I4(\i_/badr[14]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[14]_INST_0_i_10_n_0 ),
        .O(p_0_in[14]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[14]_INST_0_i_9 
       (.I0(out[14]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [14]),
        .I3(gr7_bus1),
        .O(\i_/badr[14]_INST_0_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/badr[15]_INST_0_i_12 
       (.I0(\i_/badr[15]_INST_0_i_14_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_14_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_14_0 [1]),
        .I3(abus_sel_0[6]),
        .O(gr6_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/badr[15]_INST_0_i_13 
       (.I0(\i_/badr[15]_INST_0_i_14_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_14_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_14_0 [1]),
        .I3(abus_sel_0[5]),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[15]_INST_0_i_14 
       (.I0(out[15]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [15]),
        .I3(gr7_bus1),
        .O(\i_/badr[15]_INST_0_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [15]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [15]),
        .I4(\i_/badr[15]_INST_0_i_31_n_0 ),
        .O(\i_/badr[15]_INST_0_i_15_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/badr[15]_INST_0_i_27 
       (.I0(\i_/badr[15]_INST_0_i_14_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_14_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_14_0 [1]),
        .I3(abus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/badr[15]_INST_0_i_28 
       (.I0(\i_/badr[15]_INST_0_i_14_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_14_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_14_0 [1]),
        .I3(abus_sel_0[7]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/badr[15]_INST_0_i_29 
       (.I0(\i_/badr[15]_INST_0_i_14_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_14_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_14_0 [1]),
        .I3(abus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/badr[15]_INST_0_i_30 
       (.I0(\i_/badr[15]_INST_0_i_14_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_14_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_14_0 [1]),
        .I3(abus_sel_0[4]),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[15]_INST_0_i_31 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [15]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [15]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[15]_INST_0_i_31_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[15]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [15]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [15]),
        .I3(gr5_bus1),
        .I4(\i_/badr[15]_INST_0_i_14_n_0 ),
        .I5(\i_/badr[15]_INST_0_i_15_n_0 ),
        .O(p_0_in[15]));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [1]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [1]),
        .I4(\i_/badr[1]_INST_0_i_16_n_0 ),
        .O(\i_/badr[1]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[1]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [1]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [1]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[1]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[1]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [1]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [1]),
        .I3(gr5_bus1),
        .I4(\i_/badr[1]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[1]_INST_0_i_10_n_0 ),
        .O(p_0_in[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[1]_INST_0_i_9 
       (.I0(out[1]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [1]),
        .I3(gr7_bus1),
        .O(\i_/badr[1]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [2]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [2]),
        .I4(\i_/badr[2]_INST_0_i_16_n_0 ),
        .O(\i_/badr[2]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[2]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [2]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [2]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[2]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[2]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [2]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [2]),
        .I3(gr5_bus1),
        .I4(\i_/badr[2]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[2]_INST_0_i_10_n_0 ),
        .O(p_0_in[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[2]_INST_0_i_9 
       (.I0(out[2]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [2]),
        .I3(gr7_bus1),
        .O(\i_/badr[2]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [3]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [3]),
        .I4(\i_/badr[3]_INST_0_i_16_n_0 ),
        .O(\i_/badr[3]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[3]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [3]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [3]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[3]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[3]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [3]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [3]),
        .I3(gr5_bus1),
        .I4(\i_/badr[3]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[3]_INST_0_i_10_n_0 ),
        .O(p_0_in[3]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[3]_INST_0_i_9 
       (.I0(out[3]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [3]),
        .I3(gr7_bus1),
        .O(\i_/badr[3]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [4]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [4]),
        .I4(\i_/badr[4]_INST_0_i_17_n_0 ),
        .O(\i_/badr[4]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[4]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [4]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [4]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[4]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[4]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [4]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [4]),
        .I3(gr5_bus1),
        .I4(\i_/badr[4]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[4]_INST_0_i_10_n_0 ),
        .O(p_0_in[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[4]_INST_0_i_9 
       (.I0(out[4]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [4]),
        .I3(gr7_bus1),
        .O(\i_/badr[4]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [5]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [5]),
        .I4(\i_/badr[5]_INST_0_i_16_n_0 ),
        .O(\i_/badr[5]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[5]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [5]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [5]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[5]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[5]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [5]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [5]),
        .I3(gr5_bus1),
        .I4(\i_/badr[5]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[5]_INST_0_i_10_n_0 ),
        .O(p_0_in[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[5]_INST_0_i_9 
       (.I0(out[5]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [5]),
        .I3(gr7_bus1),
        .O(\i_/badr[5]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [6]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [6]),
        .I4(\i_/badr[6]_INST_0_i_16_n_0 ),
        .O(\i_/badr[6]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[6]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [6]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [6]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[6]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[6]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [6]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [6]),
        .I3(gr5_bus1),
        .I4(\i_/badr[6]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[6]_INST_0_i_10_n_0 ),
        .O(p_0_in[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[6]_INST_0_i_9 
       (.I0(out[6]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [6]),
        .I3(gr7_bus1),
        .O(\i_/badr[6]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [7]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [7]),
        .I4(\i_/badr[7]_INST_0_i_16_n_0 ),
        .O(\i_/badr[7]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[7]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [7]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [7]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[7]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[7]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [7]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [7]),
        .I3(gr5_bus1),
        .I4(\i_/badr[7]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[7]_INST_0_i_10_n_0 ),
        .O(p_0_in[7]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[7]_INST_0_i_9 
       (.I0(out[7]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [7]),
        .I3(gr7_bus1),
        .O(\i_/badr[7]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [8]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [8]),
        .I4(\i_/badr[8]_INST_0_i_17_n_0 ),
        .O(\i_/badr[8]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[8]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [8]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [8]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[8]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[8]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [8]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [8]),
        .I3(gr5_bus1),
        .I4(\i_/badr[8]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[8]_INST_0_i_10_n_0 ),
        .O(p_0_in[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[8]_INST_0_i_9 
       (.I0(out[8]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [8]),
        .I3(gr7_bus1),
        .O(\i_/badr[8]_INST_0_i_9_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_10 
       (.I0(gr3_bus1),
        .I1(\i_/badr[15]_INST_0_i_4_1 [9]),
        .I2(gr4_bus1),
        .I3(\i_/badr[15]_INST_0_i_4_2 [9]),
        .I4(\i_/badr[9]_INST_0_i_16_n_0 ),
        .O(\i_/badr[9]_INST_0_i_10_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[9]_INST_0_i_16 
       (.I0(\i_/badr[15]_INST_0_i_15_0 [9]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_15_1 [9]),
        .I3(\i_/badr[15]_INST_0_i_15_2 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[9]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \i_/badr[9]_INST_0_i_4 
       (.I0(\mul_a_reg[15] [9]),
        .I1(gr6_bus1),
        .I2(\mul_a_reg[15]_0 [9]),
        .I3(gr5_bus1),
        .I4(\i_/badr[9]_INST_0_i_9_n_0 ),
        .I5(\i_/badr[9]_INST_0_i_10_n_0 ),
        .O(p_0_in[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/badr[9]_INST_0_i_9 
       (.I0(out[9]),
        .I1(gr0_bus1),
        .I2(\i_/badr[15]_INST_0_i_4_0 [9]),
        .I3(gr7_bus1),
        .O(\i_/badr[9]_INST_0_i_9_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_25
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_8 ,
    \i_/bdatw[15]_INST_0_i_24_0 ,
    \i_/bdatw[15]_INST_0_i_24_1 ,
    \i_/bdatw[15]_INST_0_i_24_2 ,
    \i_/bdatw[15]_INST_0_i_24_3 ,
    \i_/bdatw[15]_INST_0_i_48_0 ,
    bbus_sel_0,
    \i_/bdatw[15]_INST_0_i_48_1 ,
    \i_/bdatw[15]_INST_0_i_48_2 ,
    bank_sel,
    \i_/bdatw[15]_INST_0_i_65_0 ,
    ctl_selb_rn,
    \i_/bdatw[15]_INST_0_i_65_1 ,
    \i_/bdatw[15]_INST_0_i_65_2 ,
    ctl_selb_0,
    \i_/bdatw[15]_INST_0_i_65_3 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_8 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_24_3 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_48_0 ;
  input [5:0]bbus_sel_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_48_2 ;
  input [0:0]bank_sel;
  input \i_/bdatw[15]_INST_0_i_65_0 ;
  input [1:0]ctl_selb_rn;
  input \i_/bdatw[15]_INST_0_i_65_1 ;
  input \i_/bdatw[15]_INST_0_i_65_2 ;
  input [0:0]ctl_selb_0;
  input \i_/bdatw[15]_INST_0_i_65_3 ;

  wire [0:0]bank_sel;
  wire [5:0]bbus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_8 ;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_16_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_64_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_22_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_23_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_41_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_24_3 ;
  wire \i_/bdatw[15]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_35_n_0 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_48_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_48_2 ;
  wire \i_/bdatw[15]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_49_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_55_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_65_0 ;
  wire \i_/bdatw[15]_INST_0_i_65_1 ;
  wire \i_/bdatw[15]_INST_0_i_65_2 ;
  wire \i_/bdatw[15]_INST_0_i_65_3 ;
  wire \i_/bdatw[15]_INST_0_i_65_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_13_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_43_n_0 ;
  wire \i_/iv[15]_i_172_n_0 ;
  wire \i_/sr[7]_i_58_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [2]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [2]),
        .I4(\i_/bdatw[10]_INST_0_i_27_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [2]),
        .I2(gr4_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[10]_INST_0_i_28_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[10]_INST_0_i_21 
       (.I0(\i_/bdatw[10]_INST_0_i_35_n_0 ),
        .I1(\i_/bdatw[10]_INST_0_i_36_n_0 ),
        .I2(out[10]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [10]),
        .I5(gr3_bus1),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[10]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [2]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [2]),
        .I3(bank_sel),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[10]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [10]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [3]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [3]),
        .I4(\i_/bdatw[11]_INST_0_i_27_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [3]),
        .I2(gr4_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[11]_INST_0_i_28_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[11]_INST_0_i_21 
       (.I0(\i_/bdatw[11]_INST_0_i_35_n_0 ),
        .I1(\i_/bdatw[11]_INST_0_i_36_n_0 ),
        .I2(out[11]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [11]),
        .I5(gr3_bus1),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[11]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [3]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [3]),
        .I3(bank_sel),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[11]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [11]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [4]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [4]),
        .I4(\i_/bdatw[12]_INST_0_i_31_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_15 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [4]),
        .I2(gr4_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[12]_INST_0_i_32_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[12]_INST_0_i_25 
       (.I0(\i_/bdatw[12]_INST_0_i_39_n_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_40_n_0 ),
        .I2(out[12]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [12]),
        .I5(gr3_bus1),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[12]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [4]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [4]),
        .I3(bank_sel),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[12]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_39 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [12]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_46_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_46_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [5]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_35_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[13]_INST_0_i_14 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I3(bbus_sel_0[2]),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[13]_INST_0_i_15 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I3(bbus_sel_0[1]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_16 
       (.I0(out[5]),
        .I1(gr4_bus1),
        .I2(\bdatw[15]_INST_0_i_8 [5]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[13]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[13]_INST_0_i_29 
       (.I0(\i_/bdatw[13]_INST_0_i_49_n_0 ),
        .I1(\i_/bdatw[13]_INST_0_i_50_n_0 ),
        .I2(out[13]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [13]),
        .I5(gr3_bus1),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[13]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I3(bbus_sel_0[5]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[13]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I3(bbus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_49 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [13]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_64_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_50 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_55 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_65_0 ),
        .I2(ctl_selb_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_65_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_65_2 ),
        .I5(ctl_selb_0),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_56 
       (.I0(bank_sel),
        .I1(\i_/bdatw[15]_INST_0_i_65_3 ),
        .I2(ctl_selb_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_65_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_65_2 ),
        .I5(ctl_selb_0),
        .O(gr5_bus1));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_6 
       (.I0(\grn_reg[5]_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [5]),
        .I2(gr2_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_3 [5]),
        .I4(gr1_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_16_n_0 ),
        .O(\grn_reg[5] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_64_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[14]_INST_0_i_11 
       (.I0(\i_/bdatw[14]_INST_0_i_22_n_0 ),
        .I1(\i_/bdatw[14]_INST_0_i_23_n_0 ),
        .I2(out[6]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [6]),
        .I5(gr3_bus1),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[14]_INST_0_i_16 
       (.I0(\i_/bdatw[14]_INST_0_i_30_n_0 ),
        .I1(\i_/bdatw[14]_INST_0_i_31_n_0 ),
        .I2(out[14]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [14]),
        .I5(gr3_bus1),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_22 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [6]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_37_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_22_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [14]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[15]_INST_0_i_17 
       (.I0(\i_/bdatw[15]_INST_0_i_34_n_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_35_n_0 ),
        .I2(out[7]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [7]),
        .I5(gr3_bus1),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[15]_INST_0_i_24 
       (.I0(\i_/bdatw[15]_INST_0_i_48_n_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_49_n_0 ),
        .I2(out[15]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [15]),
        .I5(gr3_bus1),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [7]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_55_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I3(bbus_sel_0[4]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'h0D00)) 
    \i_/bdatw[15]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_48_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_48_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_48_0 [0]),
        .I3(bbus_sel_0[3]),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_48 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [15]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_65_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_49 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_49_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_55 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_55_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_65 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_65_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [0]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [0]),
        .I4(\i_/bdatw[8]_INST_0_i_27_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_13 
       (.I0(out[0]),
        .I1(gr4_bus1),
        .I2(\bdatw[15]_INST_0_i_8 [0]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_13_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[8]_INST_0_i_23 
       (.I0(\i_/bdatw[8]_INST_0_i_35_n_0 ),
        .I1(\i_/bdatw[8]_INST_0_i_36_n_0 ),
        .I2(out[8]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [8]),
        .I5(gr3_bus1),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_35 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [8]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_6 
       (.I0(\grn_reg[0]_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I2(gr2_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_3 [0]),
        .I4(gr1_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_13_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_13 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [1]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [1]),
        .I4(\i_/bdatw[9]_INST_0_i_28_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_14 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [1]),
        .I2(gr4_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[9]_INST_0_i_29_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[9]_INST_0_i_22 
       (.I0(\i_/bdatw[9]_INST_0_i_36_n_0 ),
        .I1(\i_/bdatw[9]_INST_0_i_37_n_0 ),
        .I2(out[9]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [9]),
        .I5(gr3_bus1),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[9]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [1]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [1]),
        .I3(bank_sel),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[9]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_36 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_24_0 [9]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_24_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_48_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_48_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/iv[15]_i_140 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [5]),
        .I2(gr4_bus1),
        .I3(out[5]),
        .I4(\i_/iv[15]_i_172_n_0 ),
        .O(\grn_reg[5]_1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/iv[15]_i_172 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [5]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [5]),
        .I3(bank_sel),
        .I4(bbus_sel_0[1]),
        .O(\i_/iv[15]_i_172_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/sr[7]_i_56 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [0]),
        .I2(gr4_bus1),
        .I3(out[0]),
        .I4(\i_/sr[7]_i_58_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/sr[7]_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_24_2 [0]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_24_3 [0]),
        .I3(bank_sel),
        .I4(bbus_sel_0[1]),
        .O(\i_/sr[7]_i_58_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_26
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[5]_0 ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    \grn_reg[5]_1 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_1 ,
    out,
    \bdatw[15]_INST_0_i_8 ,
    \i_/bdatw[15]_INST_0_i_23_0 ,
    \i_/bdatw[15]_INST_0_i_23_1 ,
    \i_/bdatw[15]_INST_0_i_23_2 ,
    \i_/bdatw[15]_INST_0_i_23_3 ,
    \i_/bdatw[15]_INST_0_i_46_0 ,
    bbus_sel_0,
    \i_/bdatw[15]_INST_0_i_46_1 ,
    \i_/bdatw[15]_INST_0_i_46_2 ,
    \i_/bdatw[15]_INST_0_i_64_0 ,
    \i_/bdatw[15]_INST_0_i_64_1 ,
    ctl_selb_rn,
    \i_/bdatw[15]_INST_0_i_64_2 ,
    \i_/bdatw[15]_INST_0_i_64_3 ,
    ctl_selb_0,
    \i_/bdatw[15]_INST_0_i_64_4 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[0]_0 ;
  output \grn_reg[5]_1 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_1 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_8 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_23_3 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_46_0 ;
  input [5:0]bbus_sel_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_46_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_46_2 ;
  input \i_/bdatw[15]_INST_0_i_64_0 ;
  input \i_/bdatw[15]_INST_0_i_64_1 ;
  input [1:0]ctl_selb_rn;
  input \i_/bdatw[15]_INST_0_i_64_2 ;
  input \i_/bdatw[15]_INST_0_i_64_3 ;
  input [0:0]ctl_selb_0;
  input \i_/bdatw[15]_INST_0_i_64_4 ;

  wire [5:0]bbus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_8 ;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[0]_1 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[5]_1 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_20_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_21_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_40_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_23_3 ;
  wire \i_/bdatw[15]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_31_n_0 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_46_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_46_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_46_2 ;
  wire \i_/bdatw[15]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_64_0 ;
  wire \i_/bdatw[15]_INST_0_i_64_1 ;
  wire \i_/bdatw[15]_INST_0_i_64_2 ;
  wire \i_/bdatw[15]_INST_0_i_64_3 ;
  wire \i_/bdatw[15]_INST_0_i_64_4 ;
  wire \i_/bdatw[15]_INST_0_i_64_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_15_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_28_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_42_n_0 ;
  wire \i_/iv[15]_i_171_n_0 ;
  wire \i_/sr[7]_i_57_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [2]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [2]),
        .I4(\i_/bdatw[10]_INST_0_i_25_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [2]),
        .I2(gr4_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[10]_INST_0_i_26_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[10]_INST_0_i_20 
       (.I0(\i_/bdatw[10]_INST_0_i_33_n_0 ),
        .I1(\i_/bdatw[10]_INST_0_i_34_n_0 ),
        .I2(out[10]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [10]),
        .I5(gr3_bus1),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [2]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[10]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [2]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[10]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [10]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_10 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [3]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [3]),
        .I4(\i_/bdatw[11]_INST_0_i_25_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_11 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [3]),
        .I2(gr4_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[11]_INST_0_i_26_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[11]_INST_0_i_20 
       (.I0(\i_/bdatw[11]_INST_0_i_33_n_0 ),
        .I1(\i_/bdatw[11]_INST_0_i_34_n_0 ),
        .I2(out[11]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [11]),
        .I5(gr3_bus1),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[11]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [3]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[11]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [11]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_12 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [4]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [4]),
        .I4(\i_/bdatw[12]_INST_0_i_29_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_13 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [4]),
        .I2(gr4_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[12]_INST_0_i_30_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[12]_INST_0_i_24 
       (.I0(\i_/bdatw[12]_INST_0_i_37_n_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_38_n_0 ),
        .I2(out[12]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [12]),
        .I5(gr3_bus1),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_29_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[12]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [4]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[12]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [12]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_45_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_45_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [5]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_38_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[13]_INST_0_i_18 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_46_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_46_0 [1]),
        .I3(bbus_sel_0[2]),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[13]_INST_0_i_19 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_46_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_46_0 [1]),
        .I3(bbus_sel_0[1]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_20 
       (.I0(out[5]),
        .I1(gr4_bus1),
        .I2(\bdatw[15]_INST_0_i_8 [5]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[13]_INST_0_i_20_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[13]_INST_0_i_28 
       (.I0(\i_/bdatw[13]_INST_0_i_47_n_0 ),
        .I1(\i_/bdatw[13]_INST_0_i_48_n_0 ),
        .I2(out[13]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [13]),
        .I5(gr3_bus1),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[13]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_46_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_46_0 [1]),
        .I3(bbus_sel_0[5]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[13]_INST_0_i_37 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_46_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_46_0 [1]),
        .I3(bbus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_47 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [13]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_63_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_64_4 ),
        .I2(ctl_selb_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_64_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_64_3 ),
        .I5(ctl_selb_0),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_64_1 ),
        .I2(ctl_selb_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_64_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_64_3 ),
        .I5(ctl_selb_0),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_63_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_7 
       (.I0(\grn_reg[5]_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [5]),
        .I2(gr2_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_3 [5]),
        .I4(gr1_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_20_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[14]_INST_0_i_10 
       (.I0(\i_/bdatw[14]_INST_0_i_20_n_0 ),
        .I1(\i_/bdatw[14]_INST_0_i_21_n_0 ),
        .I2(out[6]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [6]),
        .I5(gr3_bus1),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[14]_INST_0_i_15 
       (.I0(\i_/bdatw[14]_INST_0_i_28_n_0 ),
        .I1(\i_/bdatw[14]_INST_0_i_29_n_0 ),
        .I2(out[14]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [14]),
        .I5(gr3_bus1),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [6]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_36_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_20_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_21_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_28 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [14]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_40_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_28_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_36_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[15]_INST_0_i_16 
       (.I0(\i_/bdatw[15]_INST_0_i_30_n_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_31_n_0 ),
        .I2(out[7]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [7]),
        .I5(gr3_bus1),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[15]_INST_0_i_23 
       (.I0(\i_/bdatw[15]_INST_0_i_46_n_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_47_n_0 ),
        .I2(out[15]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [15]),
        .I5(gr3_bus1),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_30 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [7]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_54_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[15]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_46_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_46_0 [1]),
        .I3(bbus_sel_0[4]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'h1000)) 
    \i_/bdatw[15]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_46_0 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_46_0 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_46_0 [1]),
        .I3(bbus_sel_0[3]),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_46 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [15]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_64_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_54 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_54_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_64 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_64_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_14 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [0]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [0]),
        .I4(\i_/bdatw[8]_INST_0_i_28_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_15 
       (.I0(out[0]),
        .I1(gr4_bus1),
        .I2(\bdatw[15]_INST_0_i_8 [0]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[8]_INST_0_i_22 
       (.I0(\i_/bdatw[8]_INST_0_i_33_n_0 ),
        .I1(\i_/bdatw[8]_INST_0_i_34_n_0 ),
        .I2(out[8]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [8]),
        .I5(gr3_bus1),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_28 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [0]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_33 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [8]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_41_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_7 
       (.I0(\grn_reg[0]_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I2(gr2_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_3 [0]),
        .I4(gr1_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_15_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [1]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [1]),
        .I4(\i_/bdatw[9]_INST_0_i_26_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [1]),
        .I2(gr4_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[9]_INST_0_i_27_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[9]_INST_0_i_21 
       (.I0(\i_/bdatw[9]_INST_0_i_34_n_0 ),
        .I1(\i_/bdatw[9]_INST_0_i_35_n_0 ),
        .I2(out[9]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_8 [9]),
        .I5(gr3_bus1),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [1]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[9]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [1]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[9]_INST_0_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_34 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_23_0 [9]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_23_1 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_46_1 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_46_2 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/iv[15]_i_139 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [5]),
        .I2(gr4_bus1),
        .I3(out[5]),
        .I4(\i_/iv[15]_i_171_n_0 ),
        .O(\grn_reg[5]_1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/iv[15]_i_171 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [5]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [5]),
        .I3(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/iv[15]_i_171_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/sr[7]_i_55 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_8 [0]),
        .I2(gr4_bus1),
        .I3(out[0]),
        .I4(\i_/sr[7]_i_57_n_0 ),
        .O(\grn_reg[0]_1 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/sr[7]_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_23_2 [0]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_23_3 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_64_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/sr[7]_i_57_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_3
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \badr[15]_INST_0_i_5 ,
    \i_/badr[15]_INST_0_i_17_0 ,
    abus_sel_0,
    \i_/badr[15]_INST_0_i_17_1 ,
    \i_/badr[15]_INST_0_i_17_2 ,
    \i_/badr[15]_INST_0_i_17_3 ,
    \badr[15]_INST_0_i_5_0 ,
    \badr[15]_INST_0_i_5_1 ,
    \i_/badr[15]_INST_0_i_18_0 ,
    \i_/badr[15]_INST_0_i_18_1 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\badr[15]_INST_0_i_5 ;
  input [2:0]\i_/badr[15]_INST_0_i_17_0 ;
  input [7:0]abus_sel_0;
  input [15:0]\i_/badr[15]_INST_0_i_17_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_17_2 ;
  input \i_/badr[15]_INST_0_i_17_3 ;
  input [15:0]\badr[15]_INST_0_i_5_0 ;
  input [15:0]\badr[15]_INST_0_i_5_1 ;
  input [15:0]\i_/badr[15]_INST_0_i_18_0 ;
  input [15:0]\i_/badr[15]_INST_0_i_18_1 ;

  wire [7:0]abus_sel_0;
  wire [15:0]\badr[15]_INST_0_i_5 ;
  wire [15:0]\badr[15]_INST_0_i_5_0 ;
  wire [15:0]\badr[15]_INST_0_i_5_1 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire \i_/badr[0]_INST_0_i_17_n_0 ;
  wire \i_/badr[0]_INST_0_i_18_n_0 ;
  wire \i_/badr[10]_INST_0_i_17_n_0 ;
  wire \i_/badr[10]_INST_0_i_18_n_0 ;
  wire \i_/badr[11]_INST_0_i_17_n_0 ;
  wire \i_/badr[11]_INST_0_i_18_n_0 ;
  wire \i_/badr[12]_INST_0_i_18_n_0 ;
  wire \i_/badr[12]_INST_0_i_19_n_0 ;
  wire \i_/badr[13]_INST_0_i_17_n_0 ;
  wire \i_/badr[13]_INST_0_i_18_n_0 ;
  wire \i_/badr[14]_INST_0_i_17_n_0 ;
  wire \i_/badr[14]_INST_0_i_18_n_0 ;
  wire [2:0]\i_/badr[15]_INST_0_i_17_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_17_1 ;
  wire [15:0]\i_/badr[15]_INST_0_i_17_2 ;
  wire \i_/badr[15]_INST_0_i_17_3 ;
  wire [15:0]\i_/badr[15]_INST_0_i_18_0 ;
  wire [15:0]\i_/badr[15]_INST_0_i_18_1 ;
  wire \i_/badr[15]_INST_0_i_34_n_0 ;
  wire \i_/badr[15]_INST_0_i_37_n_0 ;
  wire \i_/badr[1]_INST_0_i_17_n_0 ;
  wire \i_/badr[1]_INST_0_i_18_n_0 ;
  wire \i_/badr[2]_INST_0_i_17_n_0 ;
  wire \i_/badr[2]_INST_0_i_18_n_0 ;
  wire \i_/badr[3]_INST_0_i_17_n_0 ;
  wire \i_/badr[3]_INST_0_i_18_n_0 ;
  wire \i_/badr[4]_INST_0_i_18_n_0 ;
  wire \i_/badr[4]_INST_0_i_19_n_0 ;
  wire \i_/badr[5]_INST_0_i_17_n_0 ;
  wire \i_/badr[5]_INST_0_i_18_n_0 ;
  wire \i_/badr[6]_INST_0_i_17_n_0 ;
  wire \i_/badr[6]_INST_0_i_18_n_0 ;
  wire \i_/badr[7]_INST_0_i_17_n_0 ;
  wire \i_/badr[7]_INST_0_i_18_n_0 ;
  wire \i_/badr[8]_INST_0_i_18_n_0 ;
  wire \i_/badr[8]_INST_0_i_19_n_0 ;
  wire \i_/badr[9]_INST_0_i_17_n_0 ;
  wire \i_/badr[9]_INST_0_i_18_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [0]),
        .I4(\i_/badr[0]_INST_0_i_17_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[0]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [0]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [0]),
        .I4(\i_/badr[0]_INST_0_i_18_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[0]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [0]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [0]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[0]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[0]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [0]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [0]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[0]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [10]),
        .I4(\i_/badr[10]_INST_0_i_17_n_0 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[10]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [10]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [10]),
        .I4(\i_/badr[10]_INST_0_i_18_n_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[10]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [10]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [10]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[10]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[10]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [10]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [10]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[10]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [11]),
        .I4(\i_/badr[11]_INST_0_i_17_n_0 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[11]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [11]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [11]),
        .I4(\i_/badr[11]_INST_0_i_18_n_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[11]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [11]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [11]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[11]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[11]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [11]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [11]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[11]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [12]),
        .I4(\i_/badr[12]_INST_0_i_18_n_0 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[12]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [12]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [12]),
        .I4(\i_/badr[12]_INST_0_i_19_n_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[12]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [12]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [12]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[12]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[12]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [12]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [12]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[12]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [13]),
        .I4(\i_/badr[13]_INST_0_i_17_n_0 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[13]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [13]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [13]),
        .I4(\i_/badr[13]_INST_0_i_18_n_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[13]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [13]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [13]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[13]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[13]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [13]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [13]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[13]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [14]),
        .I4(\i_/badr[14]_INST_0_i_17_n_0 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[14]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [14]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [14]),
        .I4(\i_/badr[14]_INST_0_i_18_n_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[14]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [14]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [14]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[14]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[14]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [14]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [14]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[14]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [15]),
        .I4(\i_/badr[15]_INST_0_i_34_n_0 ),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[15]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [15]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [15]),
        .I4(\i_/badr[15]_INST_0_i_37_n_0 ),
        .O(\grn_reg[15]_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/badr[15]_INST_0_i_32 
       (.I0(\i_/badr[15]_INST_0_i_17_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_17_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_17_0 [1]),
        .I3(abus_sel_0[7]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/badr[15]_INST_0_i_33 
       (.I0(\i_/badr[15]_INST_0_i_17_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_17_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_17_0 [1]),
        .I3(abus_sel_0[0]),
        .O(gr0_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[15]_INST_0_i_34 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [15]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [15]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[15]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/badr[15]_INST_0_i_35 
       (.I0(\i_/badr[15]_INST_0_i_17_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_17_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_17_0 [1]),
        .I3(abus_sel_0[3]),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/badr[15]_INST_0_i_36 
       (.I0(\i_/badr[15]_INST_0_i_17_0 [2]),
        .I1(\i_/badr[15]_INST_0_i_17_0 [0]),
        .I2(\i_/badr[15]_INST_0_i_17_0 [1]),
        .I3(abus_sel_0[4]),
        .O(gr4_bus1));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[15]_INST_0_i_37 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [15]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [15]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[15]_INST_0_i_37_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [1]),
        .I4(\i_/badr[1]_INST_0_i_17_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[1]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [1]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [1]),
        .I4(\i_/badr[1]_INST_0_i_18_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[1]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [1]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [1]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[1]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[1]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [1]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [1]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[1]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [2]),
        .I4(\i_/badr[2]_INST_0_i_17_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[2]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [2]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [2]),
        .I4(\i_/badr[2]_INST_0_i_18_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[2]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [2]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [2]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[2]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[2]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [2]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [2]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[2]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [3]),
        .I4(\i_/badr[3]_INST_0_i_17_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[3]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [3]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [3]),
        .I4(\i_/badr[3]_INST_0_i_18_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[3]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [3]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [3]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[3]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[3]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [3]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [3]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[3]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [4]),
        .I4(\i_/badr[4]_INST_0_i_18_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[4]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [4]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [4]),
        .I4(\i_/badr[4]_INST_0_i_19_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[4]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [4]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [4]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[4]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[4]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [4]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [4]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[4]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [5]),
        .I4(\i_/badr[5]_INST_0_i_17_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[5]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [5]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [5]),
        .I4(\i_/badr[5]_INST_0_i_18_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[5]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [5]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [5]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[5]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[5]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [5]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [5]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[5]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [6]),
        .I4(\i_/badr[6]_INST_0_i_17_n_0 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[6]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [6]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [6]),
        .I4(\i_/badr[6]_INST_0_i_18_n_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[6]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [6]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [6]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[6]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[6]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [6]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [6]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[6]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [7]),
        .I4(\i_/badr[7]_INST_0_i_17_n_0 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[7]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [7]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [7]),
        .I4(\i_/badr[7]_INST_0_i_18_n_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[7]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [7]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [7]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[7]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[7]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [7]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [7]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[7]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [8]),
        .I4(\i_/badr[8]_INST_0_i_18_n_0 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[8]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [8]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [8]),
        .I4(\i_/badr[8]_INST_0_i_19_n_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[8]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [8]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [8]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[8]_INST_0_i_18_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[8]_INST_0_i_19 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [8]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [8]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[8]_INST_0_i_19_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_11 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\badr[15]_INST_0_i_5 [9]),
        .I4(\i_/badr[9]_INST_0_i_17_n_0 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/badr[9]_INST_0_i_12 
       (.I0(gr3_bus1),
        .I1(\badr[15]_INST_0_i_5_0 [9]),
        .I2(gr4_bus1),
        .I3(\badr[15]_INST_0_i_5_1 [9]),
        .I4(\i_/badr[9]_INST_0_i_18_n_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[9]_INST_0_i_17 
       (.I0(\i_/badr[15]_INST_0_i_17_1 [9]),
        .I1(abus_sel_0[6]),
        .I2(\i_/badr[15]_INST_0_i_17_2 [9]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[5]),
        .O(\i_/badr[9]_INST_0_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/badr[9]_INST_0_i_18 
       (.I0(\i_/badr[15]_INST_0_i_18_0 [9]),
        .I1(abus_sel_0[2]),
        .I2(\i_/badr[15]_INST_0_i_18_1 [9]),
        .I3(\i_/badr[15]_INST_0_i_17_3 ),
        .I4(abus_sel_0[1]),
        .O(\i_/badr[9]_INST_0_i_18_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_4
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_9 ,
    \i_/bdatw[15]_INST_0_i_26_0 ,
    bbus_sel_0,
    \i_/bdatw[15]_INST_0_i_26_1 ,
    \i_/bdatw[15]_INST_0_i_26_2 ,
    \i_/bdatw[15]_INST_0_i_50_0 ,
    \i_/bdatw[15]_INST_0_i_50_1 ,
    \i_/bdatw[15]_INST_0_i_66_0 ,
    \i_/bdatw[15]_INST_0_i_66_1 ,
    ctl_selb_rn,
    \i_/bdatw[15]_INST_0_i_66_2 ,
    \i_/bdatw[15]_INST_0_i_66_3 ,
    ctl_selb_0,
    \i_/bdatw[15]_INST_0_i_26_3 ,
    \i_/bdatw[15]_INST_0_i_26_4 ,
    \i_/bdatw[15]_INST_0_i_66_4 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_9 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_26_0 ;
  input [5:0]bbus_sel_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_26_1 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_26_2 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_50_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_50_1 ;
  input \i_/bdatw[15]_INST_0_i_66_0 ;
  input \i_/bdatw[15]_INST_0_i_66_1 ;
  input [1:0]ctl_selb_rn;
  input \i_/bdatw[15]_INST_0_i_66_2 ;
  input \i_/bdatw[15]_INST_0_i_66_3 ;
  input [0:0]ctl_selb_0;
  input [15:0]\i_/bdatw[15]_INST_0_i_26_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_26_4 ;
  input \i_/bdatw[15]_INST_0_i_66_4 ;

  wire [5:0]bbus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_9 ;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_36_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_47_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_52_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_65_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_24_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_25_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_42_n_0 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_26_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_26_1 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_26_2 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_26_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_26_4 ;
  wire \i_/bdatw[15]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_39_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_50_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_50_1 ;
  wire \i_/bdatw[15]_INST_0_i_50_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_51_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_56_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_66_0 ;
  wire \i_/bdatw[15]_INST_0_i_66_1 ;
  wire \i_/bdatw[15]_INST_0_i_66_2 ;
  wire \i_/bdatw[15]_INST_0_i_66_3 ;
  wire \i_/bdatw[15]_INST_0_i_66_4 ;
  wire \i_/bdatw[15]_INST_0_i_66_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_37_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_38_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_44_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [2]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [2]),
        .I4(\i_/bdatw[10]_INST_0_i_31_n_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [2]),
        .I2(gr4_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[10]_INST_0_i_32_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[10]_INST_0_i_23 
       (.I0(\i_/bdatw[10]_INST_0_i_37_n_0 ),
        .I1(\i_/bdatw[10]_INST_0_i_38_n_0 ),
        .I2(out[10]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [10]),
        .I5(gr3_bus1),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [2]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[10]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [2]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [2]),
        .I3(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[10]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [10]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [10]),
        .I4(\i_/bdatw[10]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[10]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [10]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [10]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[10]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [3]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [3]),
        .I4(\i_/bdatw[11]_INST_0_i_31_n_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_18 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [3]),
        .I2(gr4_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[11]_INST_0_i_32_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[11]_INST_0_i_23 
       (.I0(\i_/bdatw[11]_INST_0_i_37_n_0 ),
        .I1(\i_/bdatw[11]_INST_0_i_38_n_0 ),
        .I2(out[11]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [11]),
        .I5(gr3_bus1),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_31_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[11]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [3]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [3]),
        .I3(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[11]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [11]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [11]),
        .I4(\i_/bdatw[11]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[11]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [11]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [11]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[11]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_19 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [4]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [4]),
        .I4(\i_/bdatw[12]_INST_0_i_35_n_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_20 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [4]),
        .I2(gr4_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[12]_INST_0_i_36_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[12]_INST_0_i_27 
       (.I0(\i_/bdatw[12]_INST_0_i_41_n_0 ),
        .I1(\i_/bdatw[12]_INST_0_i_42_n_0 ),
        .I2(out[12]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [12]),
        .I5(gr3_bus1),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_35 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[12]_INST_0_i_36 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [4]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [4]),
        .I3(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[12]_INST_0_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_41 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [12]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [12]),
        .I4(\i_/bdatw[12]_INST_0_i_47_n_0 ),
        .O(\i_/bdatw[12]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [12]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [12]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[12]_INST_0_i_42_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_47 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_47_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_22 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [5]),
        .I2(gr4_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[13]_INST_0_i_39_n_0 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_23 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [5]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [5]),
        .I4(\i_/bdatw[13]_INST_0_i_42_n_0 ),
        .O(\grn_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[13]_INST_0_i_31 
       (.I0(\i_/bdatw[13]_INST_0_i_51_n_0 ),
        .I1(\i_/bdatw[13]_INST_0_i_52_n_0 ),
        .I2(out[13]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [13]),
        .I5(gr3_bus1),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[13]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [5]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [5]),
        .I3(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[13]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[13]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_26_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_26_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_0 [0]),
        .I3(bbus_sel_0[5]),
        .O(gr7_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[13]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_26_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_26_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_0 [0]),
        .I3(bbus_sel_0[0]),
        .O(gr0_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_51 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [13]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [13]),
        .I4(\i_/bdatw[13]_INST_0_i_65_n_0 ),
        .O(\i_/bdatw[13]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [13]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [13]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[13]_INST_0_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_66_4 ),
        .I2(ctl_selb_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_66_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_66_3 ),
        .I5(ctl_selb_0),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_66_1 ),
        .I2(ctl_selb_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_66_2 ),
        .I4(\i_/bdatw[15]_INST_0_i_66_3 ),
        .I5(ctl_selb_0),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_65 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_65_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[14]_INST_0_i_13 
       (.I0(\i_/bdatw[14]_INST_0_i_24_n_0 ),
        .I1(\i_/bdatw[14]_INST_0_i_25_n_0 ),
        .I2(out[6]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [6]),
        .I5(gr3_bus1),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[14]_INST_0_i_18 
       (.I0(\i_/bdatw[14]_INST_0_i_32_n_0 ),
        .I1(\i_/bdatw[14]_INST_0_i_33_n_0 ),
        .I2(out[14]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [14]),
        .I5(gr3_bus1),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_24 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [6]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [6]),
        .I4(\i_/bdatw[14]_INST_0_i_38_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_25 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [6]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [6]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[14]_INST_0_i_32 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [14]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [14]),
        .I4(\i_/bdatw[14]_INST_0_i_42_n_0 ),
        .O(\i_/bdatw[14]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [14]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [14]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[14]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[15]_INST_0_i_20 
       (.I0(\i_/bdatw[15]_INST_0_i_38_n_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_39_n_0 ),
        .I2(out[7]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [7]),
        .I5(gr3_bus1),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[15]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_50_n_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_51_n_0 ),
        .I2(out[15]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [15]),
        .I5(gr3_bus1),
        .O(\grn_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [7]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [7]),
        .I4(\i_/bdatw[15]_INST_0_i_56_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [7]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [7]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_26_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_26_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_0 [0]),
        .I3(bbus_sel_0[4]),
        .O(gr4_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_41 
       (.I0(\i_/bdatw[15]_INST_0_i_26_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_26_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_0 [0]),
        .I3(bbus_sel_0[3]),
        .O(gr3_bus1));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[15]_INST_0_i_50 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [15]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [15]),
        .I4(\i_/bdatw[15]_INST_0_i_66_n_0 ),
        .O(\i_/bdatw[15]_INST_0_i_50_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_51 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [15]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [15]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[15]_INST_0_i_51_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_56 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_56_n_0 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_57 
       (.I0(\i_/bdatw[15]_INST_0_i_26_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_26_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_0 [0]),
        .I3(bbus_sel_0[2]),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'hD000)) 
    \i_/bdatw[15]_INST_0_i_58 
       (.I0(\i_/bdatw[15]_INST_0_i_26_0 [1]),
        .I1(\i_/bdatw[15]_INST_0_i_26_0 [2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_0 [0]),
        .I3(bbus_sel_0[1]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_66_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_17 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [0]),
        .I2(gr4_bus1),
        .I3(out[0]),
        .I4(\i_/bdatw[8]_INST_0_i_29_n_0 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [0]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [0]),
        .I4(\i_/bdatw[8]_INST_0_i_30_n_0 ),
        .O(\grn_reg[0]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[8]_INST_0_i_25 
       (.I0(\i_/bdatw[8]_INST_0_i_37_n_0 ),
        .I1(\i_/bdatw[8]_INST_0_i_38_n_0 ),
        .I2(out[8]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [8]),
        .I5(gr3_bus1),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[8]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [0]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [0]),
        .I3(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[8]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [0]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_30_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_37 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [8]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [8]),
        .I4(\i_/bdatw[8]_INST_0_i_43_n_0 ),
        .O(\i_/bdatw[8]_INST_0_i_37_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_38 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [8]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [8]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[8]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_18 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [1]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [1]),
        .I4(\i_/bdatw[9]_INST_0_i_32_n_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_19 
       (.I0(gr3_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [1]),
        .I2(gr4_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[9]_INST_0_i_33_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \i_/bdatw[9]_INST_0_i_24 
       (.I0(\i_/bdatw[9]_INST_0_i_38_n_0 ),
        .I1(\i_/bdatw[9]_INST_0_i_39_n_0 ),
        .I2(out[9]),
        .I3(gr4_bus1),
        .I4(\bdatw[15]_INST_0_i_9 [9]),
        .I5(gr3_bus1),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [1]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_32_n_0 ));
  LUT5 #(
    .INIT(32'hF8008800)) 
    \i_/bdatw[9]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [1]),
        .I1(bbus_sel_0[2]),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [1]),
        .I3(\i_/bdatw[15]_INST_0_i_66_0 ),
        .I4(bbus_sel_0[1]),
        .O(\i_/bdatw[9]_INST_0_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_38 
       (.I0(gr7_bus1),
        .I1(\i_/bdatw[15]_INST_0_i_26_1 [9]),
        .I2(gr0_bus1),
        .I3(\i_/bdatw[15]_INST_0_i_26_2 [9]),
        .I4(\i_/bdatw[9]_INST_0_i_44_n_0 ),
        .O(\i_/bdatw[9]_INST_0_i_38_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_26_3 [9]),
        .I1(gr2_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_26_4 [9]),
        .I3(gr1_bus1),
        .O(\i_/bdatw[9]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_50_0 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_50_1 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_44_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_5
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[15]_0 ,
    \grn_reg[14]_0 ,
    \grn_reg[13]_0 ,
    \grn_reg[12]_0 ,
    \grn_reg[11]_0 ,
    \grn_reg[10]_0 ,
    \grn_reg[9]_0 ,
    \grn_reg[8]_0 ,
    \grn_reg[7]_0 ,
    \grn_reg[6]_0 ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[31]_INST_0_i_5 ,
    \bdatw[31]_INST_0_i_5_0 ,
    \bdatw[30]_INST_0_i_3 ,
    \bdatw[29]_INST_0_i_3 ,
    \bdatw[28]_INST_0_i_3 ,
    \bdatw[27]_INST_0_i_3 ,
    \bdatw[26]_INST_0_i_3 ,
    \bdatw[25]_INST_0_i_3 ,
    \bdatw[24]_INST_0_i_3 ,
    \bdatw[23]_INST_0_i_3 ,
    \bdatw[22]_INST_0_i_3 ,
    \bdatw[21]_INST_0_i_3 ,
    \bdatw[20]_INST_0_i_3 ,
    \bdatw[19]_INST_0_i_3 ,
    \bdatw[18]_INST_0_i_3 ,
    \bdatw[17]_INST_0_i_3 ,
    \bdatw[16]_INST_0_i_3 ,
    \bdatw[31]_INST_0_i_5_1 ,
    \bdatw[31]_INST_0_i_5_2 ,
    \bdatw[31]_INST_0_i_5_3 ,
    \bdatw[30]_INST_0_i_3_0 ,
    \bdatw[29]_INST_0_i_3_0 ,
    \bdatw[28]_INST_0_i_3_0 ,
    \bdatw[27]_INST_0_i_3_0 ,
    \bdatw[26]_INST_0_i_3_0 ,
    \bdatw[25]_INST_0_i_3_0 ,
    \bdatw[24]_INST_0_i_3_0 ,
    \bdatw[23]_INST_0_i_3_0 ,
    \bdatw[22]_INST_0_i_3_0 ,
    \bdatw[21]_INST_0_i_3_0 ,
    \bdatw[20]_INST_0_i_3_0 ,
    \bdatw[19]_INST_0_i_3_0 ,
    \bdatw[18]_INST_0_i_3_0 ,
    \bdatw[17]_INST_0_i_3_0 ,
    \bdatw[16]_INST_0_i_3_0 ,
    \i_/bdatw[31]_INST_0_i_17_0 ,
    bbus_sel_0);
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[15]_0 ;
  output \grn_reg[14]_0 ;
  output \grn_reg[13]_0 ;
  output \grn_reg[12]_0 ;
  output \grn_reg[11]_0 ;
  output \grn_reg[10]_0 ;
  output \grn_reg[9]_0 ;
  output \grn_reg[8]_0 ;
  output \grn_reg[7]_0 ;
  output \grn_reg[6]_0 ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[31]_INST_0_i_5 ;
  input \bdatw[31]_INST_0_i_5_0 ;
  input \bdatw[30]_INST_0_i_3 ;
  input \bdatw[29]_INST_0_i_3 ;
  input \bdatw[28]_INST_0_i_3 ;
  input \bdatw[27]_INST_0_i_3 ;
  input \bdatw[26]_INST_0_i_3 ;
  input \bdatw[25]_INST_0_i_3 ;
  input \bdatw[24]_INST_0_i_3 ;
  input \bdatw[23]_INST_0_i_3 ;
  input \bdatw[22]_INST_0_i_3 ;
  input \bdatw[21]_INST_0_i_3 ;
  input \bdatw[20]_INST_0_i_3 ;
  input \bdatw[19]_INST_0_i_3 ;
  input \bdatw[18]_INST_0_i_3 ;
  input \bdatw[17]_INST_0_i_3 ;
  input \bdatw[16]_INST_0_i_3 ;
  input [15:0]\bdatw[31]_INST_0_i_5_1 ;
  input [15:0]\bdatw[31]_INST_0_i_5_2 ;
  input \bdatw[31]_INST_0_i_5_3 ;
  input \bdatw[30]_INST_0_i_3_0 ;
  input \bdatw[29]_INST_0_i_3_0 ;
  input \bdatw[28]_INST_0_i_3_0 ;
  input \bdatw[27]_INST_0_i_3_0 ;
  input \bdatw[26]_INST_0_i_3_0 ;
  input \bdatw[25]_INST_0_i_3_0 ;
  input \bdatw[24]_INST_0_i_3_0 ;
  input \bdatw[23]_INST_0_i_3_0 ;
  input \bdatw[22]_INST_0_i_3_0 ;
  input \bdatw[21]_INST_0_i_3_0 ;
  input \bdatw[20]_INST_0_i_3_0 ;
  input \bdatw[19]_INST_0_i_3_0 ;
  input \bdatw[18]_INST_0_i_3_0 ;
  input \bdatw[17]_INST_0_i_3_0 ;
  input \bdatw[16]_INST_0_i_3_0 ;
  input [1:0]\i_/bdatw[31]_INST_0_i_17_0 ;
  input [3:0]bbus_sel_0;

  wire [3:0]bbus_sel_0;
  wire \bdatw[16]_INST_0_i_3 ;
  wire \bdatw[16]_INST_0_i_3_0 ;
  wire \bdatw[17]_INST_0_i_3 ;
  wire \bdatw[17]_INST_0_i_3_0 ;
  wire \bdatw[18]_INST_0_i_3 ;
  wire \bdatw[18]_INST_0_i_3_0 ;
  wire \bdatw[19]_INST_0_i_3 ;
  wire \bdatw[19]_INST_0_i_3_0 ;
  wire \bdatw[20]_INST_0_i_3 ;
  wire \bdatw[20]_INST_0_i_3_0 ;
  wire \bdatw[21]_INST_0_i_3 ;
  wire \bdatw[21]_INST_0_i_3_0 ;
  wire \bdatw[22]_INST_0_i_3 ;
  wire \bdatw[22]_INST_0_i_3_0 ;
  wire \bdatw[23]_INST_0_i_3 ;
  wire \bdatw[23]_INST_0_i_3_0 ;
  wire \bdatw[24]_INST_0_i_3 ;
  wire \bdatw[24]_INST_0_i_3_0 ;
  wire \bdatw[25]_INST_0_i_3 ;
  wire \bdatw[25]_INST_0_i_3_0 ;
  wire \bdatw[26]_INST_0_i_3 ;
  wire \bdatw[26]_INST_0_i_3_0 ;
  wire \bdatw[27]_INST_0_i_3 ;
  wire \bdatw[27]_INST_0_i_3_0 ;
  wire \bdatw[28]_INST_0_i_3 ;
  wire \bdatw[28]_INST_0_i_3_0 ;
  wire \bdatw[29]_INST_0_i_3 ;
  wire \bdatw[29]_INST_0_i_3_0 ;
  wire \bdatw[30]_INST_0_i_3 ;
  wire \bdatw[30]_INST_0_i_3_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_5 ;
  wire \bdatw[31]_INST_0_i_5_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_5_1 ;
  wire [15:0]\bdatw[31]_INST_0_i_5_2 ;
  wire \bdatw[31]_INST_0_i_5_3 ;
  wire gr0_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[10]_0 ;
  wire \grn_reg[11] ;
  wire \grn_reg[11]_0 ;
  wire \grn_reg[12] ;
  wire \grn_reg[12]_0 ;
  wire \grn_reg[13] ;
  wire \grn_reg[13]_0 ;
  wire \grn_reg[14] ;
  wire \grn_reg[14]_0 ;
  wire \grn_reg[15] ;
  wire \grn_reg[15]_0 ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[6]_0 ;
  wire \grn_reg[7] ;
  wire \grn_reg[7]_0 ;
  wire \grn_reg[8] ;
  wire \grn_reg[8]_0 ;
  wire \grn_reg[9] ;
  wire \grn_reg[9]_0 ;
  wire [1:0]\i_/bdatw[31]_INST_0_i_17_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[16]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [0]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [0]),
        .I4(\bdatw[16]_INST_0_i_3_0 ),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[16]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[0]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [0]),
        .I4(\bdatw[16]_INST_0_i_3 ),
        .O(\grn_reg[0] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[17]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [1]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [1]),
        .I4(\bdatw[17]_INST_0_i_3_0 ),
        .O(\grn_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[17]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[1]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [1]),
        .I4(\bdatw[17]_INST_0_i_3 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[18]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [2]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [2]),
        .I4(\bdatw[18]_INST_0_i_3_0 ),
        .O(\grn_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[18]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[2]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [2]),
        .I4(\bdatw[18]_INST_0_i_3 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[19]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [3]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [3]),
        .I4(\bdatw[19]_INST_0_i_3_0 ),
        .O(\grn_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[19]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[3]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [3]),
        .I4(\bdatw[19]_INST_0_i_3 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[20]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [4]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [4]),
        .I4(\bdatw[20]_INST_0_i_3_0 ),
        .O(\grn_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[20]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[4]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [4]),
        .I4(\bdatw[20]_INST_0_i_3 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[21]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [5]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [5]),
        .I4(\bdatw[21]_INST_0_i_3_0 ),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[21]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[5]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [5]),
        .I4(\bdatw[21]_INST_0_i_3 ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[22]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [6]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [6]),
        .I4(\bdatw[22]_INST_0_i_3_0 ),
        .O(\grn_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[22]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [6]),
        .I4(\bdatw[22]_INST_0_i_3 ),
        .O(\grn_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[23]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [7]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [7]),
        .I4(\bdatw[23]_INST_0_i_3_0 ),
        .O(\grn_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[23]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [7]),
        .I4(\bdatw[23]_INST_0_i_3 ),
        .O(\grn_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[24]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [8]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [8]),
        .I4(\bdatw[24]_INST_0_i_3_0 ),
        .O(\grn_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[24]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [8]),
        .I4(\bdatw[24]_INST_0_i_3 ),
        .O(\grn_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[25]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [9]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [9]),
        .I4(\bdatw[25]_INST_0_i_3_0 ),
        .O(\grn_reg[9]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[25]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [9]),
        .I4(\bdatw[25]_INST_0_i_3 ),
        .O(\grn_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[26]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [10]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [10]),
        .I4(\bdatw[26]_INST_0_i_3_0 ),
        .O(\grn_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[26]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [10]),
        .I4(\bdatw[26]_INST_0_i_3 ),
        .O(\grn_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[27]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [11]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [11]),
        .I4(\bdatw[27]_INST_0_i_3_0 ),
        .O(\grn_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[27]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [11]),
        .I4(\bdatw[27]_INST_0_i_3 ),
        .O(\grn_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[28]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [12]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [12]),
        .I4(\bdatw[28]_INST_0_i_3_0 ),
        .O(\grn_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[28]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [12]),
        .I4(\bdatw[28]_INST_0_i_3 ),
        .O(\grn_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[29]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [13]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [13]),
        .I4(\bdatw[29]_INST_0_i_3_0 ),
        .O(\grn_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[29]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [13]),
        .I4(\bdatw[29]_INST_0_i_3 ),
        .O(\grn_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[30]_INST_0_i_8 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [14]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [14]),
        .I4(\bdatw[30]_INST_0_i_3_0 ),
        .O(\grn_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[30]_INST_0_i_9 
       (.I0(gr7_bus1),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [14]),
        .I4(\bdatw[30]_INST_0_i_3 ),
        .O(\grn_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[31]_INST_0_i_16 
       (.I0(gr3_bus1),
        .I1(\bdatw[31]_INST_0_i_5_1 [15]),
        .I2(gr4_bus1),
        .I3(\bdatw[31]_INST_0_i_5_2 [15]),
        .I4(\bdatw[31]_INST_0_i_5_3 ),
        .O(\grn_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[31]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[31]_INST_0_i_5 [15]),
        .I4(\bdatw[31]_INST_0_i_5_0 ),
        .O(\grn_reg[15] ));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_40 
       (.I0(\i_/bdatw[31]_INST_0_i_17_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_17_0 [1]),
        .I2(bbus_sel_0[1]),
        .O(gr3_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_41 
       (.I0(\i_/bdatw[31]_INST_0_i_17_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_17_0 [1]),
        .I2(bbus_sel_0[2]),
        .O(gr4_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_43 
       (.I0(\i_/bdatw[31]_INST_0_i_17_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_17_0 [1]),
        .I2(bbus_sel_0[3]),
        .O(gr7_bus1));
  LUT3 #(
    .INIT(8'h80)) 
    \i_/bdatw[31]_INST_0_i_44 
       (.I0(\i_/bdatw[31]_INST_0_i_17_0 [0]),
        .I1(\i_/bdatw[31]_INST_0_i_17_0 [1]),
        .I2(bbus_sel_0[0]),
        .O(gr0_bus1));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bank_bus" *) 
module niho_rgf_bank_bus_6
   (\grn_reg[15] ,
    \grn_reg[14] ,
    \grn_reg[13] ,
    \grn_reg[12] ,
    \grn_reg[11] ,
    \grn_reg[10] ,
    \grn_reg[9] ,
    \grn_reg[8] ,
    \grn_reg[7] ,
    \grn_reg[6] ,
    \grn_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \grn_reg[5]_0 ,
    \grn_reg[4]_0 ,
    \grn_reg[3]_0 ,
    \grn_reg[2]_0 ,
    \grn_reg[1]_0 ,
    \grn_reg[0]_0 ,
    out,
    \bdatw[15]_INST_0_i_9 ,
    \i_/bdatw[15]_INST_0_i_27_0 ,
    \i_/bdatw[15]_INST_0_i_67_0 ,
    \i_/bdatw[15]_INST_0_i_27_1 ,
    \i_/bdatw[15]_INST_0_i_27_2 ,
    ctl_selb_0,
    \i_/bdatw[15]_INST_0_i_27_3 ,
    \i_/bdatw[15]_INST_0_i_27_4 ,
    \i_/bdatw[15]_INST_0_i_27_5 ,
    \i_/bdatw[15]_INST_0_i_52_0 ,
    ctl_selb_rn,
    \i_/bdatw[15]_INST_0_i_27_6 ,
    \i_/bdatw[15]_INST_0_i_27_7 ,
    \i_/bdatw[15]_INST_0_i_53_0 ,
    \i_/bdatw[15]_INST_0_i_53_1 ,
    \i_/bdatw[15]_INST_0_i_53_2 ,
    bbus_sel_0,
    \i_/bdatw[15]_INST_0_i_67_1 ,
    \i_/bdatw[15]_INST_0_i_52_1 ,
    \i_/bdatw[15]_INST_0_i_27_8 );
  output \grn_reg[15] ;
  output \grn_reg[14] ;
  output \grn_reg[13] ;
  output \grn_reg[12] ;
  output \grn_reg[11] ;
  output \grn_reg[10] ;
  output \grn_reg[9] ;
  output \grn_reg[8] ;
  output \grn_reg[7] ;
  output \grn_reg[6] ;
  output \grn_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \grn_reg[5]_0 ;
  output \grn_reg[4]_0 ;
  output \grn_reg[3]_0 ;
  output \grn_reg[2]_0 ;
  output \grn_reg[1]_0 ;
  output \grn_reg[0]_0 ;
  input [15:0]out;
  input [15:0]\bdatw[15]_INST_0_i_9 ;
  input \i_/bdatw[15]_INST_0_i_27_0 ;
  input \i_/bdatw[15]_INST_0_i_67_0 ;
  input \i_/bdatw[15]_INST_0_i_27_1 ;
  input \i_/bdatw[15]_INST_0_i_27_2 ;
  input [0:0]ctl_selb_0;
  input \i_/bdatw[15]_INST_0_i_27_3 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_4 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_5 ;
  input \i_/bdatw[15]_INST_0_i_52_0 ;
  input [1:0]ctl_selb_rn;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_6 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_27_7 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_53_0 ;
  input [15:0]\i_/bdatw[15]_INST_0_i_53_1 ;
  input [2:0]\i_/bdatw[15]_INST_0_i_53_2 ;
  input [1:0]bbus_sel_0;
  input \i_/bdatw[15]_INST_0_i_67_1 ;
  input \i_/bdatw[15]_INST_0_i_52_1 ;
  input \i_/bdatw[15]_INST_0_i_27_8 ;

  wire [1:0]bbus_sel_0;
  wire [15:0]\bdatw[15]_INST_0_i_9 ;
  wire [0:0]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire gr0_bus1;
  wire gr1_bus1;
  wire gr2_bus1;
  wire gr3_bus1;
  wire gr4_bus1;
  wire gr5_bus1;
  wire gr6_bus1;
  wire gr7_bus1;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire \grn_reg[10] ;
  wire \grn_reg[11] ;
  wire \grn_reg[12] ;
  wire \grn_reg[13] ;
  wire \grn_reg[14] ;
  wire \grn_reg[15] ;
  wire \grn_reg[1] ;
  wire \grn_reg[1]_0 ;
  wire \grn_reg[2] ;
  wire \grn_reg[2]_0 ;
  wire \grn_reg[3] ;
  wire \grn_reg[3]_0 ;
  wire \grn_reg[4] ;
  wire \grn_reg[4]_0 ;
  wire \grn_reg[5] ;
  wire \grn_reg[5]_0 ;
  wire \grn_reg[6] ;
  wire \grn_reg[7] ;
  wire \grn_reg[8] ;
  wire \grn_reg[9] ;
  wire \i_/bdatw[10]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[10]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_29_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[11]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_33_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[12]_INST_0_i_48_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_46_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_54_n_0 ;
  wire \i_/bdatw[13]_INST_0_i_66_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_26_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_27_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_34_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_35_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[14]_INST_0_i_43_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_27_0 ;
  wire \i_/bdatw[15]_INST_0_i_27_1 ;
  wire \i_/bdatw[15]_INST_0_i_27_2 ;
  wire \i_/bdatw[15]_INST_0_i_27_3 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_4 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_5 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_6 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_27_7 ;
  wire \i_/bdatw[15]_INST_0_i_27_8 ;
  wire \i_/bdatw[15]_INST_0_i_42_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_45_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_52_0 ;
  wire \i_/bdatw[15]_INST_0_i_52_1 ;
  wire \i_/bdatw[15]_INST_0_i_52_n_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_53_0 ;
  wire [15:0]\i_/bdatw[15]_INST_0_i_53_1 ;
  wire [2:0]\i_/bdatw[15]_INST_0_i_53_2 ;
  wire \i_/bdatw[15]_INST_0_i_53_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_63_n_0 ;
  wire \i_/bdatw[15]_INST_0_i_67_0 ;
  wire \i_/bdatw[15]_INST_0_i_67_1 ;
  wire \i_/bdatw[15]_INST_0_i_67_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_32_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_39_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[8]_INST_0_i_44_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_30_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_31_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_40_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_41_n_0 ;
  wire \i_/bdatw[9]_INST_0_i_45_n_0 ;
  wire [15:0]out;

  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[10]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [2]),
        .I2(gr0_bus1),
        .I3(out[2]),
        .I4(\i_/bdatw[10]_INST_0_i_29_n_0 ),
        .O(\grn_reg[2] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_17 
       (.I0(\i_/bdatw[10]_INST_0_i_30_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [2]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [2]),
        .O(\grn_reg[2]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_24 
       (.I0(\i_/bdatw[10]_INST_0_i_39_n_0 ),
        .I1(out[10]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [10]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[10]_INST_0_i_40_n_0 ),
        .O(\grn_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [2]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [2]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [2]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [2]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[10]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [10]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [10]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[10]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[10]_INST_0_i_40 
       (.I0(\i_/bdatw[10]_INST_0_i_44_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [10]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [10]),
        .O(\i_/bdatw[10]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[10]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [10]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [10]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[10]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[11]_INST_0_i_15 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [3]),
        .I2(gr0_bus1),
        .I3(out[3]),
        .I4(\i_/bdatw[11]_INST_0_i_29_n_0 ),
        .O(\grn_reg[3] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_16 
       (.I0(\i_/bdatw[11]_INST_0_i_30_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [3]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [3]),
        .O(\grn_reg[3]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_24 
       (.I0(\i_/bdatw[11]_INST_0_i_39_n_0 ),
        .I1(out[11]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [11]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[11]_INST_0_i_40_n_0 ),
        .O(\grn_reg[11] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_29 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [3]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [3]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_29_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [3]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [3]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[11]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [11]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [11]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[11]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[11]_INST_0_i_40 
       (.I0(\i_/bdatw[11]_INST_0_i_44_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [11]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [11]),
        .O(\i_/bdatw[11]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[11]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [11]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [11]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[11]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[12]_INST_0_i_17 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [4]),
        .I2(gr0_bus1),
        .I3(out[4]),
        .I4(\i_/bdatw[12]_INST_0_i_33_n_0 ),
        .O(\grn_reg[4] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_18 
       (.I0(\i_/bdatw[12]_INST_0_i_34_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [4]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [4]),
        .O(\grn_reg[4]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_28 
       (.I0(\i_/bdatw[12]_INST_0_i_43_n_0 ),
        .I1(out[12]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [12]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[12]_INST_0_i_44_n_0 ),
        .O(\grn_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_33 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [4]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [4]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_33_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [4]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [4]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[12]_INST_0_i_34_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [12]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [12]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[12]_INST_0_i_43_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[12]_INST_0_i_44 
       (.I0(\i_/bdatw[12]_INST_0_i_48_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [12]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [12]),
        .O(\i_/bdatw[12]_INST_0_i_44_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[12]_INST_0_i_48 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [12]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [12]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[12]_INST_0_i_48_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_24 
       (.I0(\i_/bdatw[13]_INST_0_i_43_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [5]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [5]),
        .O(\grn_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[13]_INST_0_i_25 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [5]),
        .I2(gr0_bus1),
        .I3(out[5]),
        .I4(\i_/bdatw[13]_INST_0_i_46_n_0 ),
        .O(\grn_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_32 
       (.I0(\i_/bdatw[13]_INST_0_i_53_n_0 ),
        .I1(out[13]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [13]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[13]_INST_0_i_54_n_0 ),
        .O(\grn_reg[13] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [5]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [5]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[13]_INST_0_i_43_n_0 ));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[13]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_53_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_53_2 [1]),
        .I3(bbus_sel_0[0]),
        .O(gr1_bus1));
  LUT4 #(
    .INIT(16'h4000)) 
    \i_/bdatw[13]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_53_2 [2]),
        .I1(\i_/bdatw[15]_INST_0_i_53_2 [0]),
        .I2(\i_/bdatw[15]_INST_0_i_53_2 [1]),
        .I3(bbus_sel_0[1]),
        .O(gr2_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_46 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [5]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [5]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_46_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [13]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [13]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[13]_INST_0_i_53_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[13]_INST_0_i_54 
       (.I0(\i_/bdatw[13]_INST_0_i_66_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [13]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [13]),
        .O(\i_/bdatw[13]_INST_0_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_61 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_67_1 ),
        .I2(ctl_selb_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_27_2 ),
        .I5(ctl_selb_0),
        .O(gr4_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[13]_INST_0_i_62 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_27_2 ),
        .I5(ctl_selb_0),
        .O(gr3_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[13]_INST_0_i_66 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [13]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [13]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[13]_INST_0_i_66_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_14 
       (.I0(\i_/bdatw[14]_INST_0_i_26_n_0 ),
        .I1(out[6]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [6]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_27_n_0 ),
        .O(\grn_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_19 
       (.I0(\i_/bdatw[14]_INST_0_i_34_n_0 ),
        .I1(out[14]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [14]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[14]_INST_0_i_35_n_0 ),
        .O(\grn_reg[14] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_26 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [6]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [6]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_27 
       (.I0(\i_/bdatw[14]_INST_0_i_39_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [6]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [6]),
        .O(\i_/bdatw[14]_INST_0_i_27_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_34 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [14]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [14]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[14]_INST_0_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[14]_INST_0_i_35 
       (.I0(\i_/bdatw[14]_INST_0_i_43_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [14]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [14]),
        .O(\i_/bdatw[14]_INST_0_i_35_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [6]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [6]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[14]_INST_0_i_39_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[14]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [14]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [14]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[14]_INST_0_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_21 
       (.I0(\i_/bdatw[15]_INST_0_i_42_n_0 ),
        .I1(out[7]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [7]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_45_n_0 ),
        .O(\grn_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_27 
       (.I0(\i_/bdatw[15]_INST_0_i_52_n_0 ),
        .I1(out[15]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [15]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[15]_INST_0_i_53_n_0 ),
        .O(\grn_reg[15] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_42 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [7]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [7]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_42_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_43 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_27_8 ),
        .I2(\i_/bdatw[15]_INST_0_i_27_3 ),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_27_2 ),
        .I5(ctl_selb_0),
        .O(gr0_bus1));
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \i_/bdatw[15]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_67_0 ),
        .I2(\i_/bdatw[15]_INST_0_i_27_1 ),
        .I3(\i_/bdatw[15]_INST_0_i_27_2 ),
        .I4(ctl_selb_0),
        .I5(\i_/bdatw[15]_INST_0_i_27_3 ),
        .O(gr7_bus1));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_63_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [7]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [7]),
        .O(\i_/bdatw[15]_INST_0_i_45_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_52 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [15]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [15]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[15]_INST_0_i_52_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[15]_INST_0_i_53 
       (.I0(\i_/bdatw[15]_INST_0_i_67_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [15]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [15]),
        .O(\i_/bdatw[15]_INST_0_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_59 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_52_1 ),
        .I2(ctl_selb_rn[0]),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_27_2 ),
        .I5(ctl_selb_0),
        .O(gr6_bus1));
  LUT6 #(
    .INIT(64'h0000020000000000)) 
    \i_/bdatw[15]_INST_0_i_60 
       (.I0(\i_/bdatw[15]_INST_0_i_27_0 ),
        .I1(\i_/bdatw[15]_INST_0_i_52_0 ),
        .I2(ctl_selb_rn[1]),
        .I3(\i_/bdatw[15]_INST_0_i_27_1 ),
        .I4(\i_/bdatw[15]_INST_0_i_27_2 ),
        .I5(ctl_selb_0),
        .O(gr5_bus1));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_63 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [7]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [7]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[15]_INST_0_i_63_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[15]_INST_0_i_67 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [15]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [15]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[15]_INST_0_i_67_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_19 
       (.I0(\i_/bdatw[8]_INST_0_i_31_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [0]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [0]),
        .O(\grn_reg[0]_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[8]_INST_0_i_20 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [0]),
        .I2(gr0_bus1),
        .I3(out[0]),
        .I4(\i_/bdatw[8]_INST_0_i_32_n_0 ),
        .O(\grn_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_26 
       (.I0(\i_/bdatw[8]_INST_0_i_39_n_0 ),
        .I1(out[8]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [8]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[8]_INST_0_i_40_n_0 ),
        .O(\grn_reg[8] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [0]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [0]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_32 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [0]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [0]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_32_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_39 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [8]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [8]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[8]_INST_0_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[8]_INST_0_i_40 
       (.I0(\i_/bdatw[8]_INST_0_i_44_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [8]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [8]),
        .O(\i_/bdatw[8]_INST_0_i_40_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[8]_INST_0_i_44 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [8]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [8]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[8]_INST_0_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFF888)) 
    \i_/bdatw[9]_INST_0_i_16 
       (.I0(gr7_bus1),
        .I1(\bdatw[15]_INST_0_i_9 [1]),
        .I2(gr0_bus1),
        .I3(out[1]),
        .I4(\i_/bdatw[9]_INST_0_i_30_n_0 ),
        .O(\grn_reg[1] ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_17 
       (.I0(\i_/bdatw[9]_INST_0_i_31_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [1]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [1]),
        .O(\grn_reg[1]_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_25 
       (.I0(\i_/bdatw[9]_INST_0_i_40_n_0 ),
        .I1(out[9]),
        .I2(gr0_bus1),
        .I3(\bdatw[15]_INST_0_i_9 [9]),
        .I4(gr7_bus1),
        .I5(\i_/bdatw[9]_INST_0_i_41_n_0 ),
        .O(\grn_reg[9] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_30 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [1]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [1]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_31 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [1]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [1]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[9]_INST_0_i_31_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_40 
       (.I0(\i_/bdatw[15]_INST_0_i_27_4 [9]),
        .I1(gr6_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_5 [9]),
        .I3(gr5_bus1),
        .O(\i_/bdatw[9]_INST_0_i_40_n_0 ));
  LUT5 #(
    .INIT(32'hFFEAEAEA)) 
    \i_/bdatw[9]_INST_0_i_41 
       (.I0(\i_/bdatw[9]_INST_0_i_45_n_0 ),
        .I1(gr1_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_27_6 [9]),
        .I3(gr2_bus1),
        .I4(\i_/bdatw[15]_INST_0_i_27_7 [9]),
        .O(\i_/bdatw[9]_INST_0_i_41_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \i_/bdatw[9]_INST_0_i_45 
       (.I0(\i_/bdatw[15]_INST_0_i_53_0 [9]),
        .I1(gr4_bus1),
        .I2(\i_/bdatw[15]_INST_0_i_53_1 [9]),
        .I3(gr3_bus1),
        .O(\i_/bdatw[9]_INST_0_i_45_n_0 ));
endmodule

module niho_rgf_bus
   (DI,
    \sr_reg[15] ,
    \sp_reg[15] ,
    \tr_reg[11] ,
    \tr_reg[7] ,
    \tr_reg[3] ,
    \tr_reg[31] ,
    \tr_reg[30] ,
    \tr_reg[29] ,
    \tr_reg[28] ,
    \tr_reg[27] ,
    \tr_reg[26] ,
    \tr_reg[25] ,
    \tr_reg[24] ,
    \tr_reg[23] ,
    \tr_reg[22] ,
    \tr_reg[21] ,
    \tr_reg[20] ,
    \tr_reg[19] ,
    \tr_reg[18] ,
    \tr_reg[17] ,
    \tr_reg[16] ,
    \mul_a_reg[15] ,
    p_1_in,
    p_0_in,
    \mul_a_reg[14] ,
    \mul_a_reg[13] ,
    \mul_a_reg[12] ,
    \mul_a_reg[11] ,
    \mul_a_reg[10] ,
    \mul_a_reg[9] ,
    \mul_a_reg[8] ,
    \mul_a_reg[7] ,
    \mul_a_reg[6] ,
    \mul_a_reg[5] ,
    \mul_a_reg[4] ,
    \mul_a_reg[3] ,
    \mul_a_reg[2] ,
    \mul_a_reg[1] ,
    \mul_a_reg[0] ,
    out,
    abus_sel_cr,
    \mul_a_reg[15]_0 ,
    \mul_a_reg[15]_1 ,
    \mul_a_reg[15]_2 ,
    \mul_a_reg[15]_3 ,
    \mul_a_reg[14]_0 ,
    \mul_a_reg[14]_1 ,
    \mul_a_reg[14]_2 ,
    \mul_a_reg[14]_3 ,
    \mul_a_reg[13]_0 ,
    \mul_a_reg[13]_1 ,
    \mul_a_reg[13]_2 ,
    \mul_a_reg[13]_3 ,
    \mul_a_reg[12]_0 ,
    \mul_a_reg[12]_1 ,
    \mul_a_reg[12]_2 ,
    \mul_a_reg[12]_3 ,
    \mul_a_reg[11]_0 ,
    \mul_a_reg[11]_1 ,
    \mul_a_reg[11]_2 ,
    \mul_a_reg[11]_3 ,
    \mul_a_reg[10]_0 ,
    \mul_a_reg[10]_1 ,
    \mul_a_reg[10]_2 ,
    \mul_a_reg[10]_3 ,
    \mul_a_reg[9]_0 ,
    \mul_a_reg[9]_1 ,
    \mul_a_reg[9]_2 ,
    \mul_a_reg[9]_3 ,
    \mul_a_reg[8]_0 ,
    \mul_a_reg[8]_1 ,
    \mul_a_reg[8]_2 ,
    \mul_a_reg[8]_3 ,
    \mul_a_reg[7]_0 ,
    \mul_a_reg[7]_1 ,
    \mul_a_reg[7]_2 ,
    \mul_a_reg[7]_3 ,
    \mul_a_reg[6]_0 ,
    \mul_a_reg[6]_1 ,
    \mul_a_reg[6]_2 ,
    \mul_a_reg[6]_3 ,
    \mul_a_reg[5]_0 ,
    \mul_a_reg[5]_1 ,
    \mul_a_reg[5]_2 ,
    \mul_a_reg[5]_3 ,
    \mul_a_reg[4]_0 ,
    \mul_a_reg[4]_1 ,
    \mul_a_reg[4]_2 ,
    \mul_a_reg[4]_3 ,
    \mul_a_reg[3]_0 ,
    \mul_a_reg[3]_1 ,
    \mul_a_reg[3]_2 ,
    \mul_a_reg[3]_3 ,
    \mul_a_reg[2]_0 ,
    \mul_a_reg[2]_1 ,
    \mul_a_reg[2]_2 ,
    \mul_a_reg[2]_3 ,
    \mul_a_reg[1]_0 ,
    \mul_a_reg[1]_1 ,
    \mul_a_reg[1]_2 ,
    \mul_a_reg[1]_3 ,
    \mul_a_reg[0]_0 ,
    \mul_a_reg[0]_1 ,
    \mul_a_reg[0]_2 ,
    \mul_a_reg[0]_3 ,
    \mul_a_reg[32] ,
    \mul_a_reg[32]_0 ,
    \mul_a_reg[32]_1 ,
    \mul_a_reg[32]_2 ,
    \mul_a_reg[32]_3 ,
    abus_sp,
    \mul_a_reg[30] ,
    \mul_a_reg[30]_0 ,
    \mul_a_reg[30]_1 ,
    \mul_a_reg[30]_2 ,
    \mul_a_reg[30]_3 ,
    \mul_a_reg[29] ,
    \mul_a_reg[29]_0 ,
    \mul_a_reg[29]_1 ,
    \mul_a_reg[29]_2 ,
    \mul_a_reg[29]_3 ,
    \mul_a_reg[28] ,
    \mul_a_reg[28]_0 ,
    \mul_a_reg[28]_1 ,
    \mul_a_reg[28]_2 ,
    \mul_a_reg[28]_3 ,
    \mul_a_reg[27] ,
    \mul_a_reg[27]_0 ,
    \mul_a_reg[27]_1 ,
    \mul_a_reg[27]_2 ,
    \mul_a_reg[27]_3 ,
    \mul_a_reg[26] ,
    \mul_a_reg[26]_0 ,
    \mul_a_reg[26]_1 ,
    \mul_a_reg[26]_2 ,
    \mul_a_reg[26]_3 ,
    \mul_a_reg[25] ,
    \mul_a_reg[25]_0 ,
    \mul_a_reg[25]_1 ,
    \mul_a_reg[25]_2 ,
    \mul_a_reg[25]_3 ,
    \mul_a_reg[24] ,
    \mul_a_reg[24]_0 ,
    \mul_a_reg[24]_1 ,
    \mul_a_reg[24]_2 ,
    \mul_a_reg[24]_3 ,
    \mul_a_reg[23] ,
    \mul_a_reg[23]_0 ,
    \mul_a_reg[23]_1 ,
    \mul_a_reg[23]_2 ,
    \mul_a_reg[23]_3 ,
    \mul_a_reg[22] ,
    \mul_a_reg[22]_0 ,
    \mul_a_reg[22]_1 ,
    \mul_a_reg[22]_2 ,
    \mul_a_reg[22]_3 ,
    \mul_a_reg[21] ,
    \mul_a_reg[21]_0 ,
    \mul_a_reg[21]_1 ,
    \mul_a_reg[21]_2 ,
    \mul_a_reg[21]_3 ,
    \mul_a_reg[20] ,
    \mul_a_reg[20]_0 ,
    \mul_a_reg[20]_1 ,
    \mul_a_reg[20]_2 ,
    \mul_a_reg[20]_3 ,
    \mul_a_reg[19] ,
    \mul_a_reg[19]_0 ,
    \mul_a_reg[19]_1 ,
    \mul_a_reg[19]_2 ,
    \mul_a_reg[19]_3 ,
    \mul_a_reg[18] ,
    \mul_a_reg[18]_0 ,
    \mul_a_reg[18]_1 ,
    \mul_a_reg[18]_2 ,
    \mul_a_reg[18]_3 ,
    \mul_a_reg[17] ,
    \mul_a_reg[17]_0 ,
    \mul_a_reg[17]_1 ,
    \mul_a_reg[17]_2 ,
    \mul_a_reg[17]_3 ,
    \mul_a_reg[16] ,
    \mul_a_reg[16]_0 ,
    \mul_a_reg[16]_1 ,
    \mul_a_reg[16]_2 ,
    \mul_a_reg[16]_3 ,
    \mul_a_reg[15]_4 ,
    rgf_pc,
    sp_dec_0);
  output [3:0]DI;
  output \sr_reg[15] ;
  output \sp_reg[15] ;
  output [3:0]\tr_reg[11] ;
  output [3:0]\tr_reg[7] ;
  output [3:0]\tr_reg[3] ;
  output \tr_reg[31] ;
  output \tr_reg[30] ;
  output \tr_reg[29] ;
  output \tr_reg[28] ;
  output \tr_reg[27] ;
  output \tr_reg[26] ;
  output \tr_reg[25] ;
  output \tr_reg[24] ;
  output \tr_reg[23] ;
  output \tr_reg[22] ;
  output \tr_reg[21] ;
  output \tr_reg[20] ;
  output \tr_reg[19] ;
  output \tr_reg[18] ;
  output \tr_reg[17] ;
  output \tr_reg[16] ;
  input \mul_a_reg[15] ;
  input [15:0]p_1_in;
  input [15:0]p_0_in;
  input \mul_a_reg[14] ;
  input \mul_a_reg[13] ;
  input \mul_a_reg[12] ;
  input \mul_a_reg[11] ;
  input \mul_a_reg[10] ;
  input \mul_a_reg[9] ;
  input \mul_a_reg[8] ;
  input \mul_a_reg[7] ;
  input \mul_a_reg[6] ;
  input \mul_a_reg[5] ;
  input \mul_a_reg[4] ;
  input \mul_a_reg[3] ;
  input \mul_a_reg[2] ;
  input \mul_a_reg[1] ;
  input \mul_a_reg[0] ;
  input [15:0]out;
  input [3:0]abus_sel_cr;
  input \mul_a_reg[15]_0 ;
  input \mul_a_reg[15]_1 ;
  input \mul_a_reg[15]_2 ;
  input \mul_a_reg[15]_3 ;
  input \mul_a_reg[14]_0 ;
  input \mul_a_reg[14]_1 ;
  input \mul_a_reg[14]_2 ;
  input \mul_a_reg[14]_3 ;
  input \mul_a_reg[13]_0 ;
  input \mul_a_reg[13]_1 ;
  input \mul_a_reg[13]_2 ;
  input \mul_a_reg[13]_3 ;
  input \mul_a_reg[12]_0 ;
  input \mul_a_reg[12]_1 ;
  input \mul_a_reg[12]_2 ;
  input \mul_a_reg[12]_3 ;
  input \mul_a_reg[11]_0 ;
  input \mul_a_reg[11]_1 ;
  input \mul_a_reg[11]_2 ;
  input \mul_a_reg[11]_3 ;
  input \mul_a_reg[10]_0 ;
  input \mul_a_reg[10]_1 ;
  input \mul_a_reg[10]_2 ;
  input \mul_a_reg[10]_3 ;
  input \mul_a_reg[9]_0 ;
  input \mul_a_reg[9]_1 ;
  input \mul_a_reg[9]_2 ;
  input \mul_a_reg[9]_3 ;
  input \mul_a_reg[8]_0 ;
  input \mul_a_reg[8]_1 ;
  input \mul_a_reg[8]_2 ;
  input \mul_a_reg[8]_3 ;
  input \mul_a_reg[7]_0 ;
  input \mul_a_reg[7]_1 ;
  input \mul_a_reg[7]_2 ;
  input \mul_a_reg[7]_3 ;
  input \mul_a_reg[6]_0 ;
  input \mul_a_reg[6]_1 ;
  input \mul_a_reg[6]_2 ;
  input \mul_a_reg[6]_3 ;
  input \mul_a_reg[5]_0 ;
  input \mul_a_reg[5]_1 ;
  input \mul_a_reg[5]_2 ;
  input \mul_a_reg[5]_3 ;
  input \mul_a_reg[4]_0 ;
  input \mul_a_reg[4]_1 ;
  input \mul_a_reg[4]_2 ;
  input \mul_a_reg[4]_3 ;
  input \mul_a_reg[3]_0 ;
  input \mul_a_reg[3]_1 ;
  input \mul_a_reg[3]_2 ;
  input \mul_a_reg[3]_3 ;
  input \mul_a_reg[2]_0 ;
  input \mul_a_reg[2]_1 ;
  input \mul_a_reg[2]_2 ;
  input \mul_a_reg[2]_3 ;
  input \mul_a_reg[1]_0 ;
  input \mul_a_reg[1]_1 ;
  input \mul_a_reg[1]_2 ;
  input \mul_a_reg[1]_3 ;
  input \mul_a_reg[0]_0 ;
  input \mul_a_reg[0]_1 ;
  input \mul_a_reg[0]_2 ;
  input \mul_a_reg[0]_3 ;
  input \mul_a_reg[32] ;
  input \mul_a_reg[32]_0 ;
  input \mul_a_reg[32]_1 ;
  input \mul_a_reg[32]_2 ;
  input \mul_a_reg[32]_3 ;
  input [15:0]abus_sp;
  input \mul_a_reg[30] ;
  input \mul_a_reg[30]_0 ;
  input \mul_a_reg[30]_1 ;
  input \mul_a_reg[30]_2 ;
  input \mul_a_reg[30]_3 ;
  input \mul_a_reg[29] ;
  input \mul_a_reg[29]_0 ;
  input \mul_a_reg[29]_1 ;
  input \mul_a_reg[29]_2 ;
  input \mul_a_reg[29]_3 ;
  input \mul_a_reg[28] ;
  input \mul_a_reg[28]_0 ;
  input \mul_a_reg[28]_1 ;
  input \mul_a_reg[28]_2 ;
  input \mul_a_reg[28]_3 ;
  input \mul_a_reg[27] ;
  input \mul_a_reg[27]_0 ;
  input \mul_a_reg[27]_1 ;
  input \mul_a_reg[27]_2 ;
  input \mul_a_reg[27]_3 ;
  input \mul_a_reg[26] ;
  input \mul_a_reg[26]_0 ;
  input \mul_a_reg[26]_1 ;
  input \mul_a_reg[26]_2 ;
  input \mul_a_reg[26]_3 ;
  input \mul_a_reg[25] ;
  input \mul_a_reg[25]_0 ;
  input \mul_a_reg[25]_1 ;
  input \mul_a_reg[25]_2 ;
  input \mul_a_reg[25]_3 ;
  input \mul_a_reg[24] ;
  input \mul_a_reg[24]_0 ;
  input \mul_a_reg[24]_1 ;
  input \mul_a_reg[24]_2 ;
  input \mul_a_reg[24]_3 ;
  input \mul_a_reg[23] ;
  input \mul_a_reg[23]_0 ;
  input \mul_a_reg[23]_1 ;
  input \mul_a_reg[23]_2 ;
  input \mul_a_reg[23]_3 ;
  input \mul_a_reg[22] ;
  input \mul_a_reg[22]_0 ;
  input \mul_a_reg[22]_1 ;
  input \mul_a_reg[22]_2 ;
  input \mul_a_reg[22]_3 ;
  input \mul_a_reg[21] ;
  input \mul_a_reg[21]_0 ;
  input \mul_a_reg[21]_1 ;
  input \mul_a_reg[21]_2 ;
  input \mul_a_reg[21]_3 ;
  input \mul_a_reg[20] ;
  input \mul_a_reg[20]_0 ;
  input \mul_a_reg[20]_1 ;
  input \mul_a_reg[20]_2 ;
  input \mul_a_reg[20]_3 ;
  input \mul_a_reg[19] ;
  input \mul_a_reg[19]_0 ;
  input \mul_a_reg[19]_1 ;
  input \mul_a_reg[19]_2 ;
  input \mul_a_reg[19]_3 ;
  input \mul_a_reg[18] ;
  input \mul_a_reg[18]_0 ;
  input \mul_a_reg[18]_1 ;
  input \mul_a_reg[18]_2 ;
  input \mul_a_reg[18]_3 ;
  input \mul_a_reg[17] ;
  input \mul_a_reg[17]_0 ;
  input \mul_a_reg[17]_1 ;
  input \mul_a_reg[17]_2 ;
  input \mul_a_reg[17]_3 ;
  input \mul_a_reg[16] ;
  input \mul_a_reg[16]_0 ;
  input \mul_a_reg[16]_1 ;
  input \mul_a_reg[16]_2 ;
  input \mul_a_reg[16]_3 ;
  input [15:0]\mul_a_reg[15]_4 ;
  input [15:0]rgf_pc;
  input [14:0]sp_dec_0;

  wire [3:0]DI;
  wire [3:0]abus_sel_cr;
  wire [15:0]abus_sp;
  wire \badr[0]_INST_0_i_5_n_0 ;
  wire \badr[0]_INST_0_i_6_n_0 ;
  wire \badr[10]_INST_0_i_5_n_0 ;
  wire \badr[10]_INST_0_i_6_n_0 ;
  wire \badr[11]_INST_0_i_5_n_0 ;
  wire \badr[11]_INST_0_i_6_n_0 ;
  wire \badr[12]_INST_0_i_5_n_0 ;
  wire \badr[12]_INST_0_i_6_n_0 ;
  wire \badr[13]_INST_0_i_5_n_0 ;
  wire \badr[13]_INST_0_i_6_n_0 ;
  wire \badr[14]_INST_0_i_5_n_0 ;
  wire \badr[14]_INST_0_i_6_n_0 ;
  wire \badr[1]_INST_0_i_5_n_0 ;
  wire \badr[1]_INST_0_i_6_n_0 ;
  wire \badr[2]_INST_0_i_5_n_0 ;
  wire \badr[2]_INST_0_i_6_n_0 ;
  wire \badr[3]_INST_0_i_5_n_0 ;
  wire \badr[3]_INST_0_i_6_n_0 ;
  wire \badr[4]_INST_0_i_5_n_0 ;
  wire \badr[4]_INST_0_i_6_n_0 ;
  wire \badr[5]_INST_0_i_5_n_0 ;
  wire \badr[5]_INST_0_i_6_n_0 ;
  wire \badr[6]_INST_0_i_5_n_0 ;
  wire \badr[6]_INST_0_i_6_n_0 ;
  wire \badr[7]_INST_0_i_5_n_0 ;
  wire \badr[7]_INST_0_i_6_n_0 ;
  wire \badr[8]_INST_0_i_5_n_0 ;
  wire \badr[8]_INST_0_i_6_n_0 ;
  wire \badr[9]_INST_0_i_5_n_0 ;
  wire \badr[9]_INST_0_i_6_n_0 ;
  wire \mul_a_reg[0] ;
  wire \mul_a_reg[0]_0 ;
  wire \mul_a_reg[0]_1 ;
  wire \mul_a_reg[0]_2 ;
  wire \mul_a_reg[0]_3 ;
  wire \mul_a_reg[10] ;
  wire \mul_a_reg[10]_0 ;
  wire \mul_a_reg[10]_1 ;
  wire \mul_a_reg[10]_2 ;
  wire \mul_a_reg[10]_3 ;
  wire \mul_a_reg[11] ;
  wire \mul_a_reg[11]_0 ;
  wire \mul_a_reg[11]_1 ;
  wire \mul_a_reg[11]_2 ;
  wire \mul_a_reg[11]_3 ;
  wire \mul_a_reg[12] ;
  wire \mul_a_reg[12]_0 ;
  wire \mul_a_reg[12]_1 ;
  wire \mul_a_reg[12]_2 ;
  wire \mul_a_reg[12]_3 ;
  wire \mul_a_reg[13] ;
  wire \mul_a_reg[13]_0 ;
  wire \mul_a_reg[13]_1 ;
  wire \mul_a_reg[13]_2 ;
  wire \mul_a_reg[13]_3 ;
  wire \mul_a_reg[14] ;
  wire \mul_a_reg[14]_0 ;
  wire \mul_a_reg[14]_1 ;
  wire \mul_a_reg[14]_2 ;
  wire \mul_a_reg[14]_3 ;
  wire \mul_a_reg[15] ;
  wire \mul_a_reg[15]_0 ;
  wire \mul_a_reg[15]_1 ;
  wire \mul_a_reg[15]_2 ;
  wire \mul_a_reg[15]_3 ;
  wire [15:0]\mul_a_reg[15]_4 ;
  wire \mul_a_reg[16] ;
  wire \mul_a_reg[16]_0 ;
  wire \mul_a_reg[16]_1 ;
  wire \mul_a_reg[16]_2 ;
  wire \mul_a_reg[16]_3 ;
  wire \mul_a_reg[17] ;
  wire \mul_a_reg[17]_0 ;
  wire \mul_a_reg[17]_1 ;
  wire \mul_a_reg[17]_2 ;
  wire \mul_a_reg[17]_3 ;
  wire \mul_a_reg[18] ;
  wire \mul_a_reg[18]_0 ;
  wire \mul_a_reg[18]_1 ;
  wire \mul_a_reg[18]_2 ;
  wire \mul_a_reg[18]_3 ;
  wire \mul_a_reg[19] ;
  wire \mul_a_reg[19]_0 ;
  wire \mul_a_reg[19]_1 ;
  wire \mul_a_reg[19]_2 ;
  wire \mul_a_reg[19]_3 ;
  wire \mul_a_reg[1] ;
  wire \mul_a_reg[1]_0 ;
  wire \mul_a_reg[1]_1 ;
  wire \mul_a_reg[1]_2 ;
  wire \mul_a_reg[1]_3 ;
  wire \mul_a_reg[20] ;
  wire \mul_a_reg[20]_0 ;
  wire \mul_a_reg[20]_1 ;
  wire \mul_a_reg[20]_2 ;
  wire \mul_a_reg[20]_3 ;
  wire \mul_a_reg[21] ;
  wire \mul_a_reg[21]_0 ;
  wire \mul_a_reg[21]_1 ;
  wire \mul_a_reg[21]_2 ;
  wire \mul_a_reg[21]_3 ;
  wire \mul_a_reg[22] ;
  wire \mul_a_reg[22]_0 ;
  wire \mul_a_reg[22]_1 ;
  wire \mul_a_reg[22]_2 ;
  wire \mul_a_reg[22]_3 ;
  wire \mul_a_reg[23] ;
  wire \mul_a_reg[23]_0 ;
  wire \mul_a_reg[23]_1 ;
  wire \mul_a_reg[23]_2 ;
  wire \mul_a_reg[23]_3 ;
  wire \mul_a_reg[24] ;
  wire \mul_a_reg[24]_0 ;
  wire \mul_a_reg[24]_1 ;
  wire \mul_a_reg[24]_2 ;
  wire \mul_a_reg[24]_3 ;
  wire \mul_a_reg[25] ;
  wire \mul_a_reg[25]_0 ;
  wire \mul_a_reg[25]_1 ;
  wire \mul_a_reg[25]_2 ;
  wire \mul_a_reg[25]_3 ;
  wire \mul_a_reg[26] ;
  wire \mul_a_reg[26]_0 ;
  wire \mul_a_reg[26]_1 ;
  wire \mul_a_reg[26]_2 ;
  wire \mul_a_reg[26]_3 ;
  wire \mul_a_reg[27] ;
  wire \mul_a_reg[27]_0 ;
  wire \mul_a_reg[27]_1 ;
  wire \mul_a_reg[27]_2 ;
  wire \mul_a_reg[27]_3 ;
  wire \mul_a_reg[28] ;
  wire \mul_a_reg[28]_0 ;
  wire \mul_a_reg[28]_1 ;
  wire \mul_a_reg[28]_2 ;
  wire \mul_a_reg[28]_3 ;
  wire \mul_a_reg[29] ;
  wire \mul_a_reg[29]_0 ;
  wire \mul_a_reg[29]_1 ;
  wire \mul_a_reg[29]_2 ;
  wire \mul_a_reg[29]_3 ;
  wire \mul_a_reg[2] ;
  wire \mul_a_reg[2]_0 ;
  wire \mul_a_reg[2]_1 ;
  wire \mul_a_reg[2]_2 ;
  wire \mul_a_reg[2]_3 ;
  wire \mul_a_reg[30] ;
  wire \mul_a_reg[30]_0 ;
  wire \mul_a_reg[30]_1 ;
  wire \mul_a_reg[30]_2 ;
  wire \mul_a_reg[30]_3 ;
  wire \mul_a_reg[32] ;
  wire \mul_a_reg[32]_0 ;
  wire \mul_a_reg[32]_1 ;
  wire \mul_a_reg[32]_2 ;
  wire \mul_a_reg[32]_3 ;
  wire \mul_a_reg[3] ;
  wire \mul_a_reg[3]_0 ;
  wire \mul_a_reg[3]_1 ;
  wire \mul_a_reg[3]_2 ;
  wire \mul_a_reg[3]_3 ;
  wire \mul_a_reg[4] ;
  wire \mul_a_reg[4]_0 ;
  wire \mul_a_reg[4]_1 ;
  wire \mul_a_reg[4]_2 ;
  wire \mul_a_reg[4]_3 ;
  wire \mul_a_reg[5] ;
  wire \mul_a_reg[5]_0 ;
  wire \mul_a_reg[5]_1 ;
  wire \mul_a_reg[5]_2 ;
  wire \mul_a_reg[5]_3 ;
  wire \mul_a_reg[6] ;
  wire \mul_a_reg[6]_0 ;
  wire \mul_a_reg[6]_1 ;
  wire \mul_a_reg[6]_2 ;
  wire \mul_a_reg[6]_3 ;
  wire \mul_a_reg[7] ;
  wire \mul_a_reg[7]_0 ;
  wire \mul_a_reg[7]_1 ;
  wire \mul_a_reg[7]_2 ;
  wire \mul_a_reg[7]_3 ;
  wire \mul_a_reg[8] ;
  wire \mul_a_reg[8]_0 ;
  wire \mul_a_reg[8]_1 ;
  wire \mul_a_reg[8]_2 ;
  wire \mul_a_reg[8]_3 ;
  wire \mul_a_reg[9] ;
  wire \mul_a_reg[9]_0 ;
  wire \mul_a_reg[9]_1 ;
  wire \mul_a_reg[9]_2 ;
  wire \mul_a_reg[9]_3 ;
  wire [15:0]out;
  wire [15:0]p_0_in;
  wire [15:0]p_1_in;
  wire [15:0]rgf_pc;
  wire [14:0]sp_dec_0;
  wire \sp_reg[15] ;
  wire \sr_reg[15] ;
  wire [3:0]\tr_reg[11] ;
  wire \tr_reg[16] ;
  wire \tr_reg[17] ;
  wire \tr_reg[18] ;
  wire \tr_reg[19] ;
  wire \tr_reg[20] ;
  wire \tr_reg[21] ;
  wire \tr_reg[22] ;
  wire \tr_reg[23] ;
  wire \tr_reg[24] ;
  wire \tr_reg[25] ;
  wire \tr_reg[26] ;
  wire \tr_reg[27] ;
  wire \tr_reg[28] ;
  wire \tr_reg[29] ;
  wire \tr_reg[30] ;
  wire \tr_reg[31] ;
  wire [3:0]\tr_reg[3] ;
  wire [3:0]\tr_reg[7] ;

  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[0]_INST_0_i_1 
       (.I0(\mul_a_reg[0] ),
        .I1(p_1_in[0]),
        .I2(p_0_in[0]),
        .I3(\badr[0]_INST_0_i_5_n_0 ),
        .I4(\badr[0]_INST_0_i_6_n_0 ),
        .O(\tr_reg[3] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[0]_INST_0_i_5 
       (.I0(out[0]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[0]_0 ),
        .I3(\mul_a_reg[0]_1 ),
        .I4(\mul_a_reg[0]_2 ),
        .I5(\mul_a_reg[0]_3 ),
        .O(\badr[0]_INST_0_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \badr[0]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(\mul_a_reg[15]_4 [0]),
        .I2(abus_sel_cr[2]),
        .I3(rgf_pc[0]),
        .I4(abus_sel_cr[1]),
        .O(\badr[0]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[10]_INST_0_i_1 
       (.I0(\mul_a_reg[10] ),
        .I1(p_1_in[10]),
        .I2(p_0_in[10]),
        .I3(\badr[10]_INST_0_i_5_n_0 ),
        .I4(\badr[10]_INST_0_i_6_n_0 ),
        .O(\tr_reg[11] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[10]_INST_0_i_5 
       (.I0(out[10]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[10]_0 ),
        .I3(\mul_a_reg[10]_1 ),
        .I4(\mul_a_reg[10]_2 ),
        .I5(\mul_a_reg[10]_3 ),
        .O(\badr[10]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[10]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[9]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [10]),
        .I4(rgf_pc[10]),
        .I5(abus_sel_cr[1]),
        .O(\badr[10]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[11]_INST_0_i_1 
       (.I0(\mul_a_reg[11] ),
        .I1(p_1_in[11]),
        .I2(p_0_in[11]),
        .I3(\badr[11]_INST_0_i_5_n_0 ),
        .I4(\badr[11]_INST_0_i_6_n_0 ),
        .O(\tr_reg[11] [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[11]_INST_0_i_5 
       (.I0(out[11]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[11]_0 ),
        .I3(\mul_a_reg[11]_1 ),
        .I4(\mul_a_reg[11]_2 ),
        .I5(\mul_a_reg[11]_3 ),
        .O(\badr[11]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[11]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[10]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [11]),
        .I4(rgf_pc[11]),
        .I5(abus_sel_cr[1]),
        .O(\badr[11]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[12]_INST_0_i_1 
       (.I0(\mul_a_reg[12] ),
        .I1(p_1_in[12]),
        .I2(p_0_in[12]),
        .I3(\badr[12]_INST_0_i_5_n_0 ),
        .I4(\badr[12]_INST_0_i_6_n_0 ),
        .O(DI[0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[12]_INST_0_i_5 
       (.I0(out[12]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[12]_0 ),
        .I3(\mul_a_reg[12]_1 ),
        .I4(\mul_a_reg[12]_2 ),
        .I5(\mul_a_reg[12]_3 ),
        .O(\badr[12]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[12]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[11]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [12]),
        .I4(rgf_pc[12]),
        .I5(abus_sel_cr[1]),
        .O(\badr[12]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[13]_INST_0_i_1 
       (.I0(\mul_a_reg[13] ),
        .I1(p_1_in[13]),
        .I2(p_0_in[13]),
        .I3(\badr[13]_INST_0_i_5_n_0 ),
        .I4(\badr[13]_INST_0_i_6_n_0 ),
        .O(DI[1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[13]_INST_0_i_5 
       (.I0(out[13]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[13]_0 ),
        .I3(\mul_a_reg[13]_1 ),
        .I4(\mul_a_reg[13]_2 ),
        .I5(\mul_a_reg[13]_3 ),
        .O(\badr[13]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[13]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[12]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [13]),
        .I4(rgf_pc[13]),
        .I5(abus_sel_cr[1]),
        .O(\badr[13]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[14]_INST_0_i_1 
       (.I0(\mul_a_reg[14] ),
        .I1(p_1_in[14]),
        .I2(p_0_in[14]),
        .I3(\badr[14]_INST_0_i_5_n_0 ),
        .I4(\badr[14]_INST_0_i_6_n_0 ),
        .O(DI[2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[14]_INST_0_i_5 
       (.I0(out[14]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[14]_0 ),
        .I3(\mul_a_reg[14]_1 ),
        .I4(\mul_a_reg[14]_2 ),
        .I5(\mul_a_reg[14]_3 ),
        .O(\badr[14]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[14]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[13]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [14]),
        .I4(rgf_pc[14]),
        .I5(abus_sel_cr[1]),
        .O(\badr[14]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[15]_INST_0_i_1 
       (.I0(\mul_a_reg[15] ),
        .I1(p_1_in[15]),
        .I2(p_0_in[15]),
        .I3(\sr_reg[15] ),
        .I4(\sp_reg[15] ),
        .O(DI[3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[15]_INST_0_i_5 
       (.I0(out[15]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[15]_0 ),
        .I3(\mul_a_reg[15]_1 ),
        .I4(\mul_a_reg[15]_2 ),
        .I5(\mul_a_reg[15]_3 ),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[15]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[14]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [15]),
        .I4(rgf_pc[15]),
        .I5(abus_sel_cr[1]),
        .O(\sp_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[16]_INST_0_i_1 
       (.I0(\mul_a_reg[16] ),
        .I1(\mul_a_reg[16]_0 ),
        .I2(\mul_a_reg[16]_1 ),
        .I3(\mul_a_reg[16]_2 ),
        .I4(\mul_a_reg[16]_3 ),
        .I5(abus_sp[0]),
        .O(\tr_reg[16] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[17]_INST_0_i_1 
       (.I0(\mul_a_reg[17] ),
        .I1(\mul_a_reg[17]_0 ),
        .I2(\mul_a_reg[17]_1 ),
        .I3(\mul_a_reg[17]_2 ),
        .I4(\mul_a_reg[17]_3 ),
        .I5(abus_sp[1]),
        .O(\tr_reg[17] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[18]_INST_0_i_1 
       (.I0(\mul_a_reg[18] ),
        .I1(\mul_a_reg[18]_0 ),
        .I2(\mul_a_reg[18]_1 ),
        .I3(\mul_a_reg[18]_2 ),
        .I4(\mul_a_reg[18]_3 ),
        .I5(abus_sp[2]),
        .O(\tr_reg[18] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[19]_INST_0_i_1 
       (.I0(\mul_a_reg[19] ),
        .I1(\mul_a_reg[19]_0 ),
        .I2(\mul_a_reg[19]_1 ),
        .I3(\mul_a_reg[19]_2 ),
        .I4(\mul_a_reg[19]_3 ),
        .I5(abus_sp[3]),
        .O(\tr_reg[19] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[1]_INST_0_i_1 
       (.I0(\mul_a_reg[1] ),
        .I1(p_1_in[1]),
        .I2(p_0_in[1]),
        .I3(\badr[1]_INST_0_i_5_n_0 ),
        .I4(\badr[1]_INST_0_i_6_n_0 ),
        .O(\tr_reg[3] [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[1]_INST_0_i_5 
       (.I0(out[1]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[1]_0 ),
        .I3(\mul_a_reg[1]_1 ),
        .I4(\mul_a_reg[1]_2 ),
        .I5(\mul_a_reg[1]_3 ),
        .O(\badr[1]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[1]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[0]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [1]),
        .I4(rgf_pc[1]),
        .I5(abus_sel_cr[1]),
        .O(\badr[1]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[20]_INST_0_i_1 
       (.I0(\mul_a_reg[20] ),
        .I1(\mul_a_reg[20]_0 ),
        .I2(\mul_a_reg[20]_1 ),
        .I3(\mul_a_reg[20]_2 ),
        .I4(\mul_a_reg[20]_3 ),
        .I5(abus_sp[4]),
        .O(\tr_reg[20] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[21]_INST_0_i_1 
       (.I0(\mul_a_reg[21] ),
        .I1(\mul_a_reg[21]_0 ),
        .I2(\mul_a_reg[21]_1 ),
        .I3(\mul_a_reg[21]_2 ),
        .I4(\mul_a_reg[21]_3 ),
        .I5(abus_sp[5]),
        .O(\tr_reg[21] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[22]_INST_0_i_1 
       (.I0(\mul_a_reg[22] ),
        .I1(\mul_a_reg[22]_0 ),
        .I2(\mul_a_reg[22]_1 ),
        .I3(\mul_a_reg[22]_2 ),
        .I4(\mul_a_reg[22]_3 ),
        .I5(abus_sp[6]),
        .O(\tr_reg[22] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[23]_INST_0_i_1 
       (.I0(\mul_a_reg[23] ),
        .I1(\mul_a_reg[23]_0 ),
        .I2(\mul_a_reg[23]_1 ),
        .I3(\mul_a_reg[23]_2 ),
        .I4(\mul_a_reg[23]_3 ),
        .I5(abus_sp[7]),
        .O(\tr_reg[23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[24]_INST_0_i_1 
       (.I0(\mul_a_reg[24] ),
        .I1(\mul_a_reg[24]_0 ),
        .I2(\mul_a_reg[24]_1 ),
        .I3(\mul_a_reg[24]_2 ),
        .I4(\mul_a_reg[24]_3 ),
        .I5(abus_sp[8]),
        .O(\tr_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[25]_INST_0_i_1 
       (.I0(\mul_a_reg[25] ),
        .I1(\mul_a_reg[25]_0 ),
        .I2(\mul_a_reg[25]_1 ),
        .I3(\mul_a_reg[25]_2 ),
        .I4(\mul_a_reg[25]_3 ),
        .I5(abus_sp[9]),
        .O(\tr_reg[25] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[26]_INST_0_i_1 
       (.I0(\mul_a_reg[26] ),
        .I1(\mul_a_reg[26]_0 ),
        .I2(\mul_a_reg[26]_1 ),
        .I3(\mul_a_reg[26]_2 ),
        .I4(\mul_a_reg[26]_3 ),
        .I5(abus_sp[10]),
        .O(\tr_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[27]_INST_0_i_1 
       (.I0(\mul_a_reg[27] ),
        .I1(\mul_a_reg[27]_0 ),
        .I2(\mul_a_reg[27]_1 ),
        .I3(\mul_a_reg[27]_2 ),
        .I4(\mul_a_reg[27]_3 ),
        .I5(abus_sp[11]),
        .O(\tr_reg[27] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[28]_INST_0_i_1 
       (.I0(\mul_a_reg[28] ),
        .I1(\mul_a_reg[28]_0 ),
        .I2(\mul_a_reg[28]_1 ),
        .I3(\mul_a_reg[28]_2 ),
        .I4(\mul_a_reg[28]_3 ),
        .I5(abus_sp[12]),
        .O(\tr_reg[28] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[29]_INST_0_i_1 
       (.I0(\mul_a_reg[29] ),
        .I1(\mul_a_reg[29]_0 ),
        .I2(\mul_a_reg[29]_1 ),
        .I3(\mul_a_reg[29]_2 ),
        .I4(\mul_a_reg[29]_3 ),
        .I5(abus_sp[13]),
        .O(\tr_reg[29] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[2]_INST_0_i_1 
       (.I0(\mul_a_reg[2] ),
        .I1(p_1_in[2]),
        .I2(p_0_in[2]),
        .I3(\badr[2]_INST_0_i_5_n_0 ),
        .I4(\badr[2]_INST_0_i_6_n_0 ),
        .O(\tr_reg[3] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[2]_INST_0_i_5 
       (.I0(out[2]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[2]_0 ),
        .I3(\mul_a_reg[2]_1 ),
        .I4(\mul_a_reg[2]_2 ),
        .I5(\mul_a_reg[2]_3 ),
        .O(\badr[2]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[2]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[1]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [2]),
        .I4(rgf_pc[2]),
        .I5(abus_sel_cr[1]),
        .O(\badr[2]_INST_0_i_6_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[30]_INST_0_i_1 
       (.I0(\mul_a_reg[30] ),
        .I1(\mul_a_reg[30]_0 ),
        .I2(\mul_a_reg[30]_1 ),
        .I3(\mul_a_reg[30]_2 ),
        .I4(\mul_a_reg[30]_3 ),
        .I5(abus_sp[14]),
        .O(\tr_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \badr[31]_INST_0_i_1 
       (.I0(\mul_a_reg[32] ),
        .I1(\mul_a_reg[32]_0 ),
        .I2(\mul_a_reg[32]_1 ),
        .I3(\mul_a_reg[32]_2 ),
        .I4(\mul_a_reg[32]_3 ),
        .I5(abus_sp[15]),
        .O(\tr_reg[31] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[3]_INST_0_i_1 
       (.I0(\mul_a_reg[3] ),
        .I1(p_1_in[3]),
        .I2(p_0_in[3]),
        .I3(\badr[3]_INST_0_i_5_n_0 ),
        .I4(\badr[3]_INST_0_i_6_n_0 ),
        .O(\tr_reg[3] [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[3]_INST_0_i_5 
       (.I0(out[3]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[3]_0 ),
        .I3(\mul_a_reg[3]_1 ),
        .I4(\mul_a_reg[3]_2 ),
        .I5(\mul_a_reg[3]_3 ),
        .O(\badr[3]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[3]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[2]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [3]),
        .I4(rgf_pc[3]),
        .I5(abus_sel_cr[1]),
        .O(\badr[3]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[4]_INST_0_i_1 
       (.I0(\mul_a_reg[4] ),
        .I1(p_1_in[4]),
        .I2(p_0_in[4]),
        .I3(\badr[4]_INST_0_i_5_n_0 ),
        .I4(\badr[4]_INST_0_i_6_n_0 ),
        .O(\tr_reg[7] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[4]_INST_0_i_5 
       (.I0(out[4]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[4]_0 ),
        .I3(\mul_a_reg[4]_1 ),
        .I4(\mul_a_reg[4]_2 ),
        .I5(\mul_a_reg[4]_3 ),
        .O(\badr[4]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[4]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[3]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [4]),
        .I4(rgf_pc[4]),
        .I5(abus_sel_cr[1]),
        .O(\badr[4]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[5]_INST_0_i_1 
       (.I0(\mul_a_reg[5] ),
        .I1(p_1_in[5]),
        .I2(p_0_in[5]),
        .I3(\badr[5]_INST_0_i_5_n_0 ),
        .I4(\badr[5]_INST_0_i_6_n_0 ),
        .O(\tr_reg[7] [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[5]_INST_0_i_5 
       (.I0(out[5]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[5]_0 ),
        .I3(\mul_a_reg[5]_1 ),
        .I4(\mul_a_reg[5]_2 ),
        .I5(\mul_a_reg[5]_3 ),
        .O(\badr[5]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[5]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[4]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [5]),
        .I4(rgf_pc[5]),
        .I5(abus_sel_cr[1]),
        .O(\badr[5]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[6]_INST_0_i_1 
       (.I0(\mul_a_reg[6] ),
        .I1(p_1_in[6]),
        .I2(p_0_in[6]),
        .I3(\badr[6]_INST_0_i_5_n_0 ),
        .I4(\badr[6]_INST_0_i_6_n_0 ),
        .O(\tr_reg[7] [2]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[6]_INST_0_i_5 
       (.I0(out[6]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[6]_0 ),
        .I3(\mul_a_reg[6]_1 ),
        .I4(\mul_a_reg[6]_2 ),
        .I5(\mul_a_reg[6]_3 ),
        .O(\badr[6]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[6]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[5]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [6]),
        .I4(rgf_pc[6]),
        .I5(abus_sel_cr[1]),
        .O(\badr[6]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[7]_INST_0_i_1 
       (.I0(\mul_a_reg[7] ),
        .I1(p_1_in[7]),
        .I2(p_0_in[7]),
        .I3(\badr[7]_INST_0_i_5_n_0 ),
        .I4(\badr[7]_INST_0_i_6_n_0 ),
        .O(\tr_reg[7] [3]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[7]_INST_0_i_5 
       (.I0(out[7]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[7]_0 ),
        .I3(\mul_a_reg[7]_1 ),
        .I4(\mul_a_reg[7]_2 ),
        .I5(\mul_a_reg[7]_3 ),
        .O(\badr[7]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[7]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[6]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [7]),
        .I4(rgf_pc[7]),
        .I5(abus_sel_cr[1]),
        .O(\badr[7]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[8]_INST_0_i_1 
       (.I0(\mul_a_reg[8] ),
        .I1(p_1_in[8]),
        .I2(p_0_in[8]),
        .I3(\badr[8]_INST_0_i_5_n_0 ),
        .I4(\badr[8]_INST_0_i_6_n_0 ),
        .O(\tr_reg[11] [0]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[8]_INST_0_i_5 
       (.I0(out[8]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[8]_0 ),
        .I3(\mul_a_reg[8]_1 ),
        .I4(\mul_a_reg[8]_2 ),
        .I5(\mul_a_reg[8]_3 ),
        .O(\badr[8]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[8]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[7]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [8]),
        .I4(rgf_pc[8]),
        .I5(abus_sel_cr[1]),
        .O(\badr[8]_INST_0_i_6_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \badr[9]_INST_0_i_1 
       (.I0(\mul_a_reg[9] ),
        .I1(p_1_in[9]),
        .I2(p_0_in[9]),
        .I3(\badr[9]_INST_0_i_5_n_0 ),
        .I4(\badr[9]_INST_0_i_6_n_0 ),
        .O(\tr_reg[11] [1]));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \badr[9]_INST_0_i_5 
       (.I0(out[9]),
        .I1(abus_sel_cr[0]),
        .I2(\mul_a_reg[9]_0 ),
        .I3(\mul_a_reg[9]_1 ),
        .I4(\mul_a_reg[9]_2 ),
        .I5(\mul_a_reg[9]_3 ),
        .O(\badr[9]_INST_0_i_5_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \badr[9]_INST_0_i_6 
       (.I0(abus_sel_cr[3]),
        .I1(sp_dec_0[8]),
        .I2(abus_sel_cr[2]),
        .I3(\mul_a_reg[15]_4 [9]),
        .I4(rgf_pc[9]),
        .I5(abus_sel_cr[1]),
        .O(\badr[9]_INST_0_i_6_n_0 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_bus" *) 
module niho_rgf_bus_1
   (\iv_reg[15] ,
    \iv_reg[14] ,
    \iv_reg[13] ,
    \iv_reg[12] ,
    \iv_reg[11] ,
    \iv_reg[10] ,
    \iv_reg[9] ,
    \iv_reg[8] ,
    \iv_reg[7] ,
    \iv_reg[6] ,
    \grn_reg[5] ,
    \tr_reg[5] ,
    \grn_reg[4] ,
    \grn_reg[3] ,
    \grn_reg[2] ,
    \grn_reg[1] ,
    \grn_reg[0] ,
    \tr_reg[0] ,
    \sr_reg[15] ,
    \sr_reg[14] ,
    \sr_reg[13] ,
    \sr_reg[12] ,
    \sr_reg[11] ,
    \sr_reg[10] ,
    \sr_reg[9] ,
    \sr_reg[8] ,
    \sr_reg[7] ,
    \sr_reg[6] ,
    \sp_reg[5] ,
    \sp_reg[5]_0 ,
    \sr_reg[5] ,
    \sr_reg[4] ,
    \sr_reg[3] ,
    \sr_reg[2] ,
    \sr_reg[1] ,
    \sp_reg[0] ,
    \sp_reg[31] ,
    \sp_reg[30] ,
    \sp_reg[29] ,
    \sp_reg[28] ,
    \sp_reg[27] ,
    \sp_reg[26] ,
    \sp_reg[25] ,
    \sp_reg[24] ,
    \sp_reg[23] ,
    \sp_reg[22] ,
    \sp_reg[21] ,
    \sp_reg[20] ,
    \sp_reg[19] ,
    \sp_reg[18] ,
    \sp_reg[17] ,
    \sp_reg[16] ,
    \tr_reg[31] ,
    \tr_reg[30] ,
    \tr_reg[29] ,
    \tr_reg[28] ,
    \tr_reg[27] ,
    \tr_reg[26] ,
    \tr_reg[25] ,
    \tr_reg[24] ,
    \tr_reg[23] ,
    \tr_reg[22] ,
    \tr_reg[21] ,
    \tr_reg[20] ,
    \tr_reg[19] ,
    \tr_reg[18] ,
    \tr_reg[17] ,
    \tr_reg[16] ,
    \sp_reg[1] ,
    \sp_reg[2] ,
    \sp_reg[3] ,
    \sp_reg[4] ,
    \mul_b_reg[15] ,
    \mul_b_reg[15]_0 ,
    bbus_sel_cr,
    \mul_b_reg[15]_1 ,
    \bdatw[31]_INST_0_i_1 ,
    \mul_b_reg[14] ,
    \mul_b_reg[14]_0 ,
    \mul_b_reg[13] ,
    \mul_b_reg[13]_0 ,
    \mul_b_reg[12] ,
    \mul_b_reg[12]_0 ,
    \mul_b_reg[11] ,
    \mul_b_reg[11]_0 ,
    \mul_b_reg[10] ,
    \mul_b_reg[10]_0 ,
    \mul_b_reg[9] ,
    \mul_b_reg[9]_0 ,
    \mul_b_reg[8] ,
    \mul_b_reg[8]_0 ,
    \mul_b_reg[7] ,
    \mul_b_reg[7]_0 ,
    \mul_b_reg[6] ,
    \mul_b_reg[6]_0 ,
    \iv[15]_i_56 ,
    \iv[15]_i_56_0 ,
    \iv[15]_i_56_1 ,
    \iv[15]_i_56_2 ,
    \mul_b_reg[4] ,
    \mul_b_reg[4]_0 ,
    \mul_b_reg[4]_1 ,
    \mul_b_reg[4]_2 ,
    \mul_b_reg[3] ,
    \mul_b_reg[3]_0 ,
    \mul_b_reg[3]_1 ,
    \mul_b_reg[3]_2 ,
    \mul_b_reg[2] ,
    \mul_b_reg[2]_0 ,
    \mul_b_reg[2]_1 ,
    \mul_b_reg[2]_2 ,
    \mul_b_reg[1] ,
    \mul_b_reg[1]_0 ,
    \mul_b_reg[1]_1 ,
    \mul_b_reg[1]_2 ,
    \iv[12]_i_51 ,
    \iv[12]_i_51_0 ,
    \iv[12]_i_51_1 ,
    \iv[12]_i_51_2 ,
    \mul_b_reg[15]_2 ,
    \mul_b_reg[15]_3 ,
    out,
    \mul_b_reg[14]_1 ,
    \mul_b_reg[14]_2 ,
    \mul_b_reg[13]_1 ,
    \mul_b_reg[13]_2 ,
    \mul_b_reg[12]_1 ,
    \mul_b_reg[12]_2 ,
    \mul_b_reg[11]_1 ,
    \mul_b_reg[11]_2 ,
    \mul_b_reg[10]_1 ,
    \mul_b_reg[10]_2 ,
    \mul_b_reg[9]_1 ,
    \mul_b_reg[9]_2 ,
    \mul_b_reg[8]_1 ,
    \mul_b_reg[8]_2 ,
    \mul_b_reg[7]_1 ,
    \mul_b_reg[7]_2 ,
    \mul_b_reg[6]_1 ,
    \mul_b_reg[6]_2 ,
    \mul_b_reg[5] ,
    \mul_b_reg[5]_0 ,
    \mul_b_reg[5]_1 ,
    \mul_b_reg[5]_2 ,
    bbus_sr,
    \mul_b_reg[4]_3 ,
    \mul_b_reg[4]_4 ,
    \mul_b_reg[4]_5 ,
    \mul_b_reg[4]_6 ,
    \mul_b_reg[3]_3 ,
    \mul_b_reg[3]_4 ,
    \mul_b_reg[3]_5 ,
    \mul_b_reg[3]_6 ,
    \mul_b_reg[2]_3 ,
    \mul_b_reg[2]_4 ,
    \mul_b_reg[2]_5 ,
    \mul_b_reg[2]_6 ,
    \mul_b_reg[1]_3 ,
    \mul_b_reg[1]_4 ,
    \mul_b_reg[1]_5 ,
    \mul_b_reg[1]_6 ,
    \mul_b_reg[0] ,
    \mul_b_reg[0]_0 ,
    \mul_b_reg[0]_1 ,
    \mul_b_reg[0]_2 ,
    sp_dec_0,
    \bdatw[31]_INST_0_i_1_0 ,
    \bdatw[31]_INST_0_i_1_1 ,
    \bdatw[31]_INST_0_i_1_2 ,
    \bdatw[30]_INST_0_i_1 ,
    \bdatw[30]_INST_0_i_1_0 ,
    \bdatw[29]_INST_0_i_1 ,
    \bdatw[29]_INST_0_i_1_0 ,
    \bdatw[28]_INST_0_i_1 ,
    \bdatw[28]_INST_0_i_1_0 ,
    \bdatw[27]_INST_0_i_1 ,
    \bdatw[27]_INST_0_i_1_0 ,
    \bdatw[26]_INST_0_i_1 ,
    \bdatw[26]_INST_0_i_1_0 ,
    \bdatw[25]_INST_0_i_1 ,
    \bdatw[25]_INST_0_i_1_0 ,
    \bdatw[24]_INST_0_i_1 ,
    \bdatw[24]_INST_0_i_1_0 ,
    \bdatw[23]_INST_0_i_1 ,
    \bdatw[23]_INST_0_i_1_0 ,
    \bdatw[22]_INST_0_i_1 ,
    \bdatw[22]_INST_0_i_1_0 ,
    \bdatw[21]_INST_0_i_1 ,
    \bdatw[21]_INST_0_i_1_0 ,
    \bdatw[20]_INST_0_i_1 ,
    \bdatw[20]_INST_0_i_1_0 ,
    \bdatw[19]_INST_0_i_1 ,
    \bdatw[19]_INST_0_i_1_0 ,
    \bdatw[18]_INST_0_i_1 ,
    \bdatw[18]_INST_0_i_1_0 ,
    \bdatw[17]_INST_0_i_1 ,
    \bdatw[17]_INST_0_i_1_0 ,
    \bdatw[16]_INST_0_i_1 ,
    \bdatw[16]_INST_0_i_1_0 ,
    \bdatw[31]_INST_0_i_1_3 ,
    \bdatw[31]_INST_0_i_1_4 ,
    \bdatw[31]_INST_0_i_1_5 ,
    \bdatw[31]_INST_0_i_1_6 ,
    \bdatw[30]_INST_0_i_1_1 ,
    \bdatw[30]_INST_0_i_1_2 ,
    \bdatw[30]_INST_0_i_1_3 ,
    \bdatw[30]_INST_0_i_1_4 ,
    \bdatw[29]_INST_0_i_1_1 ,
    \bdatw[29]_INST_0_i_1_2 ,
    \bdatw[29]_INST_0_i_1_3 ,
    \bdatw[29]_INST_0_i_1_4 ,
    \bdatw[28]_INST_0_i_1_1 ,
    \bdatw[28]_INST_0_i_1_2 ,
    \bdatw[28]_INST_0_i_1_3 ,
    \bdatw[28]_INST_0_i_1_4 ,
    \bdatw[27]_INST_0_i_1_1 ,
    \bdatw[27]_INST_0_i_1_2 ,
    \bdatw[27]_INST_0_i_1_3 ,
    \bdatw[27]_INST_0_i_1_4 ,
    \bdatw[26]_INST_0_i_1_1 ,
    \bdatw[26]_INST_0_i_1_2 ,
    \bdatw[26]_INST_0_i_1_3 ,
    \bdatw[26]_INST_0_i_1_4 ,
    \bdatw[25]_INST_0_i_1_1 ,
    \bdatw[25]_INST_0_i_1_2 ,
    \bdatw[25]_INST_0_i_1_3 ,
    \bdatw[25]_INST_0_i_1_4 ,
    \bdatw[24]_INST_0_i_1_1 ,
    \bdatw[24]_INST_0_i_1_2 ,
    \bdatw[24]_INST_0_i_1_3 ,
    \bdatw[24]_INST_0_i_1_4 ,
    \bdatw[23]_INST_0_i_1_1 ,
    \bdatw[23]_INST_0_i_1_2 ,
    \bdatw[23]_INST_0_i_1_3 ,
    \bdatw[23]_INST_0_i_1_4 ,
    \bdatw[22]_INST_0_i_1_1 ,
    \bdatw[22]_INST_0_i_1_2 ,
    \bdatw[22]_INST_0_i_1_3 ,
    \bdatw[22]_INST_0_i_1_4 ,
    \bdatw[21]_INST_0_i_1_1 ,
    \bdatw[21]_INST_0_i_1_2 ,
    \bdatw[21]_INST_0_i_1_3 ,
    \bdatw[21]_INST_0_i_1_4 ,
    \bdatw[20]_INST_0_i_1_1 ,
    \bdatw[20]_INST_0_i_1_2 ,
    \bdatw[20]_INST_0_i_1_3 ,
    \bdatw[20]_INST_0_i_1_4 ,
    \bdatw[19]_INST_0_i_1_1 ,
    \bdatw[19]_INST_0_i_1_2 ,
    \bdatw[19]_INST_0_i_1_3 ,
    \bdatw[19]_INST_0_i_1_4 ,
    \bdatw[18]_INST_0_i_1_1 ,
    \bdatw[18]_INST_0_i_1_2 ,
    \bdatw[18]_INST_0_i_1_3 ,
    \bdatw[18]_INST_0_i_1_4 ,
    \bdatw[17]_INST_0_i_1_1 ,
    \bdatw[17]_INST_0_i_1_2 ,
    \bdatw[17]_INST_0_i_1_3 ,
    \bdatw[17]_INST_0_i_1_4 ,
    \bdatw[16]_INST_0_i_1_1 ,
    \bdatw[16]_INST_0_i_1_2 ,
    \bdatw[16]_INST_0_i_1_3 ,
    \bdatw[16]_INST_0_i_1_4 ,
    \bdatw[15]_INST_0_i_9_0 );
  output \iv_reg[15] ;
  output \iv_reg[14] ;
  output \iv_reg[13] ;
  output \iv_reg[12] ;
  output \iv_reg[11] ;
  output \iv_reg[10] ;
  output \iv_reg[9] ;
  output \iv_reg[8] ;
  output \iv_reg[7] ;
  output \iv_reg[6] ;
  output \grn_reg[5] ;
  output \tr_reg[5] ;
  output \grn_reg[4] ;
  output \grn_reg[3] ;
  output \grn_reg[2] ;
  output \grn_reg[1] ;
  output \grn_reg[0] ;
  output \tr_reg[0] ;
  output \sr_reg[15] ;
  output \sr_reg[14] ;
  output \sr_reg[13] ;
  output \sr_reg[12] ;
  output \sr_reg[11] ;
  output \sr_reg[10] ;
  output \sr_reg[9] ;
  output \sr_reg[8] ;
  output \sr_reg[7] ;
  output \sr_reg[6] ;
  output \sp_reg[5] ;
  output \sp_reg[5]_0 ;
  output \sr_reg[5] ;
  output \sr_reg[4] ;
  output \sr_reg[3] ;
  output \sr_reg[2] ;
  output \sr_reg[1] ;
  output \sp_reg[0] ;
  output \sp_reg[31] ;
  output \sp_reg[30] ;
  output \sp_reg[29] ;
  output \sp_reg[28] ;
  output \sp_reg[27] ;
  output \sp_reg[26] ;
  output \sp_reg[25] ;
  output \sp_reg[24] ;
  output \sp_reg[23] ;
  output \sp_reg[22] ;
  output \sp_reg[21] ;
  output \sp_reg[20] ;
  output \sp_reg[19] ;
  output \sp_reg[18] ;
  output \sp_reg[17] ;
  output \sp_reg[16] ;
  output \tr_reg[31] ;
  output \tr_reg[30] ;
  output \tr_reg[29] ;
  output \tr_reg[28] ;
  output \tr_reg[27] ;
  output \tr_reg[26] ;
  output \tr_reg[25] ;
  output \tr_reg[24] ;
  output \tr_reg[23] ;
  output \tr_reg[22] ;
  output \tr_reg[21] ;
  output \tr_reg[20] ;
  output \tr_reg[19] ;
  output \tr_reg[18] ;
  output \tr_reg[17] ;
  output \tr_reg[16] ;
  output \sp_reg[1] ;
  output \sp_reg[2] ;
  output \sp_reg[3] ;
  output \sp_reg[4] ;
  input \mul_b_reg[15] ;
  input \mul_b_reg[15]_0 ;
  input [5:0]bbus_sel_cr;
  input [15:0]\mul_b_reg[15]_1 ;
  input [31:0]\bdatw[31]_INST_0_i_1 ;
  input \mul_b_reg[14] ;
  input \mul_b_reg[14]_0 ;
  input \mul_b_reg[13] ;
  input \mul_b_reg[13]_0 ;
  input \mul_b_reg[12] ;
  input \mul_b_reg[12]_0 ;
  input \mul_b_reg[11] ;
  input \mul_b_reg[11]_0 ;
  input \mul_b_reg[10] ;
  input \mul_b_reg[10]_0 ;
  input \mul_b_reg[9] ;
  input \mul_b_reg[9]_0 ;
  input \mul_b_reg[8] ;
  input \mul_b_reg[8]_0 ;
  input \mul_b_reg[7] ;
  input \mul_b_reg[7]_0 ;
  input \mul_b_reg[6] ;
  input \mul_b_reg[6]_0 ;
  input \iv[15]_i_56 ;
  input \iv[15]_i_56_0 ;
  input \iv[15]_i_56_1 ;
  input \iv[15]_i_56_2 ;
  input \mul_b_reg[4] ;
  input \mul_b_reg[4]_0 ;
  input \mul_b_reg[4]_1 ;
  input \mul_b_reg[4]_2 ;
  input \mul_b_reg[3] ;
  input \mul_b_reg[3]_0 ;
  input \mul_b_reg[3]_1 ;
  input \mul_b_reg[3]_2 ;
  input \mul_b_reg[2] ;
  input \mul_b_reg[2]_0 ;
  input \mul_b_reg[2]_1 ;
  input \mul_b_reg[2]_2 ;
  input \mul_b_reg[1] ;
  input \mul_b_reg[1]_0 ;
  input \mul_b_reg[1]_1 ;
  input \mul_b_reg[1]_2 ;
  input \iv[12]_i_51 ;
  input \iv[12]_i_51_0 ;
  input \iv[12]_i_51_1 ;
  input \iv[12]_i_51_2 ;
  input \mul_b_reg[15]_2 ;
  input \mul_b_reg[15]_3 ;
  input [14:0]out;
  input \mul_b_reg[14]_1 ;
  input \mul_b_reg[14]_2 ;
  input \mul_b_reg[13]_1 ;
  input \mul_b_reg[13]_2 ;
  input \mul_b_reg[12]_1 ;
  input \mul_b_reg[12]_2 ;
  input \mul_b_reg[11]_1 ;
  input \mul_b_reg[11]_2 ;
  input \mul_b_reg[10]_1 ;
  input \mul_b_reg[10]_2 ;
  input \mul_b_reg[9]_1 ;
  input \mul_b_reg[9]_2 ;
  input \mul_b_reg[8]_1 ;
  input \mul_b_reg[8]_2 ;
  input \mul_b_reg[7]_1 ;
  input \mul_b_reg[7]_2 ;
  input \mul_b_reg[6]_1 ;
  input \mul_b_reg[6]_2 ;
  input \mul_b_reg[5] ;
  input \mul_b_reg[5]_0 ;
  input \mul_b_reg[5]_1 ;
  input \mul_b_reg[5]_2 ;
  input [1:0]bbus_sr;
  input \mul_b_reg[4]_3 ;
  input \mul_b_reg[4]_4 ;
  input \mul_b_reg[4]_5 ;
  input \mul_b_reg[4]_6 ;
  input \mul_b_reg[3]_3 ;
  input \mul_b_reg[3]_4 ;
  input \mul_b_reg[3]_5 ;
  input \mul_b_reg[3]_6 ;
  input \mul_b_reg[2]_3 ;
  input \mul_b_reg[2]_4 ;
  input \mul_b_reg[2]_5 ;
  input \mul_b_reg[2]_6 ;
  input \mul_b_reg[1]_3 ;
  input \mul_b_reg[1]_4 ;
  input \mul_b_reg[1]_5 ;
  input \mul_b_reg[1]_6 ;
  input \mul_b_reg[0] ;
  input \mul_b_reg[0]_0 ;
  input \mul_b_reg[0]_1 ;
  input \mul_b_reg[0]_2 ;
  input [30:0]sp_dec_0;
  input [31:0]\bdatw[31]_INST_0_i_1_0 ;
  input \bdatw[31]_INST_0_i_1_1 ;
  input \bdatw[31]_INST_0_i_1_2 ;
  input \bdatw[30]_INST_0_i_1 ;
  input \bdatw[30]_INST_0_i_1_0 ;
  input \bdatw[29]_INST_0_i_1 ;
  input \bdatw[29]_INST_0_i_1_0 ;
  input \bdatw[28]_INST_0_i_1 ;
  input \bdatw[28]_INST_0_i_1_0 ;
  input \bdatw[27]_INST_0_i_1 ;
  input \bdatw[27]_INST_0_i_1_0 ;
  input \bdatw[26]_INST_0_i_1 ;
  input \bdatw[26]_INST_0_i_1_0 ;
  input \bdatw[25]_INST_0_i_1 ;
  input \bdatw[25]_INST_0_i_1_0 ;
  input \bdatw[24]_INST_0_i_1 ;
  input \bdatw[24]_INST_0_i_1_0 ;
  input \bdatw[23]_INST_0_i_1 ;
  input \bdatw[23]_INST_0_i_1_0 ;
  input \bdatw[22]_INST_0_i_1 ;
  input \bdatw[22]_INST_0_i_1_0 ;
  input \bdatw[21]_INST_0_i_1 ;
  input \bdatw[21]_INST_0_i_1_0 ;
  input \bdatw[20]_INST_0_i_1 ;
  input \bdatw[20]_INST_0_i_1_0 ;
  input \bdatw[19]_INST_0_i_1 ;
  input \bdatw[19]_INST_0_i_1_0 ;
  input \bdatw[18]_INST_0_i_1 ;
  input \bdatw[18]_INST_0_i_1_0 ;
  input \bdatw[17]_INST_0_i_1 ;
  input \bdatw[17]_INST_0_i_1_0 ;
  input \bdatw[16]_INST_0_i_1 ;
  input \bdatw[16]_INST_0_i_1_0 ;
  input \bdatw[31]_INST_0_i_1_3 ;
  input \bdatw[31]_INST_0_i_1_4 ;
  input \bdatw[31]_INST_0_i_1_5 ;
  input \bdatw[31]_INST_0_i_1_6 ;
  input \bdatw[30]_INST_0_i_1_1 ;
  input \bdatw[30]_INST_0_i_1_2 ;
  input \bdatw[30]_INST_0_i_1_3 ;
  input \bdatw[30]_INST_0_i_1_4 ;
  input \bdatw[29]_INST_0_i_1_1 ;
  input \bdatw[29]_INST_0_i_1_2 ;
  input \bdatw[29]_INST_0_i_1_3 ;
  input \bdatw[29]_INST_0_i_1_4 ;
  input \bdatw[28]_INST_0_i_1_1 ;
  input \bdatw[28]_INST_0_i_1_2 ;
  input \bdatw[28]_INST_0_i_1_3 ;
  input \bdatw[28]_INST_0_i_1_4 ;
  input \bdatw[27]_INST_0_i_1_1 ;
  input \bdatw[27]_INST_0_i_1_2 ;
  input \bdatw[27]_INST_0_i_1_3 ;
  input \bdatw[27]_INST_0_i_1_4 ;
  input \bdatw[26]_INST_0_i_1_1 ;
  input \bdatw[26]_INST_0_i_1_2 ;
  input \bdatw[26]_INST_0_i_1_3 ;
  input \bdatw[26]_INST_0_i_1_4 ;
  input \bdatw[25]_INST_0_i_1_1 ;
  input \bdatw[25]_INST_0_i_1_2 ;
  input \bdatw[25]_INST_0_i_1_3 ;
  input \bdatw[25]_INST_0_i_1_4 ;
  input \bdatw[24]_INST_0_i_1_1 ;
  input \bdatw[24]_INST_0_i_1_2 ;
  input \bdatw[24]_INST_0_i_1_3 ;
  input \bdatw[24]_INST_0_i_1_4 ;
  input \bdatw[23]_INST_0_i_1_1 ;
  input \bdatw[23]_INST_0_i_1_2 ;
  input \bdatw[23]_INST_0_i_1_3 ;
  input \bdatw[23]_INST_0_i_1_4 ;
  input \bdatw[22]_INST_0_i_1_1 ;
  input \bdatw[22]_INST_0_i_1_2 ;
  input \bdatw[22]_INST_0_i_1_3 ;
  input \bdatw[22]_INST_0_i_1_4 ;
  input \bdatw[21]_INST_0_i_1_1 ;
  input \bdatw[21]_INST_0_i_1_2 ;
  input \bdatw[21]_INST_0_i_1_3 ;
  input \bdatw[21]_INST_0_i_1_4 ;
  input \bdatw[20]_INST_0_i_1_1 ;
  input \bdatw[20]_INST_0_i_1_2 ;
  input \bdatw[20]_INST_0_i_1_3 ;
  input \bdatw[20]_INST_0_i_1_4 ;
  input \bdatw[19]_INST_0_i_1_1 ;
  input \bdatw[19]_INST_0_i_1_2 ;
  input \bdatw[19]_INST_0_i_1_3 ;
  input \bdatw[19]_INST_0_i_1_4 ;
  input \bdatw[18]_INST_0_i_1_1 ;
  input \bdatw[18]_INST_0_i_1_2 ;
  input \bdatw[18]_INST_0_i_1_3 ;
  input \bdatw[18]_INST_0_i_1_4 ;
  input \bdatw[17]_INST_0_i_1_1 ;
  input \bdatw[17]_INST_0_i_1_2 ;
  input \bdatw[17]_INST_0_i_1_3 ;
  input \bdatw[17]_INST_0_i_1_4 ;
  input \bdatw[16]_INST_0_i_1_1 ;
  input \bdatw[16]_INST_0_i_1_2 ;
  input \bdatw[16]_INST_0_i_1_3 ;
  input \bdatw[16]_INST_0_i_1_4 ;
  input [15:0]\bdatw[15]_INST_0_i_9_0 ;

  wire [5:0]bbus_sel_cr;
  wire [1:0]bbus_sr;
  wire \bdatw[10]_INST_0_i_15_n_0 ;
  wire \bdatw[10]_INST_0_i_22_n_0 ;
  wire \bdatw[11]_INST_0_i_14_n_0 ;
  wire \bdatw[11]_INST_0_i_22_n_0 ;
  wire \bdatw[12]_INST_0_i_16_n_0 ;
  wire \bdatw[12]_INST_0_i_26_n_0 ;
  wire \bdatw[13]_INST_0_i_30_n_0 ;
  wire \bdatw[14]_INST_0_i_12_n_0 ;
  wire \bdatw[14]_INST_0_i_17_n_0 ;
  wire \bdatw[15]_INST_0_i_19_n_0 ;
  wire \bdatw[15]_INST_0_i_25_n_0 ;
  wire [15:0]\bdatw[15]_INST_0_i_9_0 ;
  wire \bdatw[16]_INST_0_i_1 ;
  wire \bdatw[16]_INST_0_i_1_0 ;
  wire \bdatw[16]_INST_0_i_1_1 ;
  wire \bdatw[16]_INST_0_i_1_2 ;
  wire \bdatw[16]_INST_0_i_1_3 ;
  wire \bdatw[16]_INST_0_i_1_4 ;
  wire \bdatw[17]_INST_0_i_1 ;
  wire \bdatw[17]_INST_0_i_1_0 ;
  wire \bdatw[17]_INST_0_i_1_1 ;
  wire \bdatw[17]_INST_0_i_1_2 ;
  wire \bdatw[17]_INST_0_i_1_3 ;
  wire \bdatw[17]_INST_0_i_1_4 ;
  wire \bdatw[18]_INST_0_i_1 ;
  wire \bdatw[18]_INST_0_i_1_0 ;
  wire \bdatw[18]_INST_0_i_1_1 ;
  wire \bdatw[18]_INST_0_i_1_2 ;
  wire \bdatw[18]_INST_0_i_1_3 ;
  wire \bdatw[18]_INST_0_i_1_4 ;
  wire \bdatw[19]_INST_0_i_1 ;
  wire \bdatw[19]_INST_0_i_1_0 ;
  wire \bdatw[19]_INST_0_i_1_1 ;
  wire \bdatw[19]_INST_0_i_1_2 ;
  wire \bdatw[19]_INST_0_i_1_3 ;
  wire \bdatw[19]_INST_0_i_1_4 ;
  wire \bdatw[20]_INST_0_i_1 ;
  wire \bdatw[20]_INST_0_i_1_0 ;
  wire \bdatw[20]_INST_0_i_1_1 ;
  wire \bdatw[20]_INST_0_i_1_2 ;
  wire \bdatw[20]_INST_0_i_1_3 ;
  wire \bdatw[20]_INST_0_i_1_4 ;
  wire \bdatw[21]_INST_0_i_1 ;
  wire \bdatw[21]_INST_0_i_1_0 ;
  wire \bdatw[21]_INST_0_i_1_1 ;
  wire \bdatw[21]_INST_0_i_1_2 ;
  wire \bdatw[21]_INST_0_i_1_3 ;
  wire \bdatw[21]_INST_0_i_1_4 ;
  wire \bdatw[22]_INST_0_i_1 ;
  wire \bdatw[22]_INST_0_i_1_0 ;
  wire \bdatw[22]_INST_0_i_1_1 ;
  wire \bdatw[22]_INST_0_i_1_2 ;
  wire \bdatw[22]_INST_0_i_1_3 ;
  wire \bdatw[22]_INST_0_i_1_4 ;
  wire \bdatw[23]_INST_0_i_1 ;
  wire \bdatw[23]_INST_0_i_1_0 ;
  wire \bdatw[23]_INST_0_i_1_1 ;
  wire \bdatw[23]_INST_0_i_1_2 ;
  wire \bdatw[23]_INST_0_i_1_3 ;
  wire \bdatw[23]_INST_0_i_1_4 ;
  wire \bdatw[24]_INST_0_i_1 ;
  wire \bdatw[24]_INST_0_i_1_0 ;
  wire \bdatw[24]_INST_0_i_1_1 ;
  wire \bdatw[24]_INST_0_i_1_2 ;
  wire \bdatw[24]_INST_0_i_1_3 ;
  wire \bdatw[24]_INST_0_i_1_4 ;
  wire \bdatw[25]_INST_0_i_1 ;
  wire \bdatw[25]_INST_0_i_1_0 ;
  wire \bdatw[25]_INST_0_i_1_1 ;
  wire \bdatw[25]_INST_0_i_1_2 ;
  wire \bdatw[25]_INST_0_i_1_3 ;
  wire \bdatw[25]_INST_0_i_1_4 ;
  wire \bdatw[26]_INST_0_i_1 ;
  wire \bdatw[26]_INST_0_i_1_0 ;
  wire \bdatw[26]_INST_0_i_1_1 ;
  wire \bdatw[26]_INST_0_i_1_2 ;
  wire \bdatw[26]_INST_0_i_1_3 ;
  wire \bdatw[26]_INST_0_i_1_4 ;
  wire \bdatw[27]_INST_0_i_1 ;
  wire \bdatw[27]_INST_0_i_1_0 ;
  wire \bdatw[27]_INST_0_i_1_1 ;
  wire \bdatw[27]_INST_0_i_1_2 ;
  wire \bdatw[27]_INST_0_i_1_3 ;
  wire \bdatw[27]_INST_0_i_1_4 ;
  wire \bdatw[28]_INST_0_i_1 ;
  wire \bdatw[28]_INST_0_i_1_0 ;
  wire \bdatw[28]_INST_0_i_1_1 ;
  wire \bdatw[28]_INST_0_i_1_2 ;
  wire \bdatw[28]_INST_0_i_1_3 ;
  wire \bdatw[28]_INST_0_i_1_4 ;
  wire \bdatw[29]_INST_0_i_1 ;
  wire \bdatw[29]_INST_0_i_1_0 ;
  wire \bdatw[29]_INST_0_i_1_1 ;
  wire \bdatw[29]_INST_0_i_1_2 ;
  wire \bdatw[29]_INST_0_i_1_3 ;
  wire \bdatw[29]_INST_0_i_1_4 ;
  wire \bdatw[30]_INST_0_i_1 ;
  wire \bdatw[30]_INST_0_i_1_0 ;
  wire \bdatw[30]_INST_0_i_1_1 ;
  wire \bdatw[30]_INST_0_i_1_2 ;
  wire \bdatw[30]_INST_0_i_1_3 ;
  wire \bdatw[30]_INST_0_i_1_4 ;
  wire [31:0]\bdatw[31]_INST_0_i_1 ;
  wire [31:0]\bdatw[31]_INST_0_i_1_0 ;
  wire \bdatw[31]_INST_0_i_1_1 ;
  wire \bdatw[31]_INST_0_i_1_2 ;
  wire \bdatw[31]_INST_0_i_1_3 ;
  wire \bdatw[31]_INST_0_i_1_4 ;
  wire \bdatw[31]_INST_0_i_1_5 ;
  wire \bdatw[31]_INST_0_i_1_6 ;
  wire \bdatw[8]_INST_0_i_16_n_0 ;
  wire \bdatw[8]_INST_0_i_24_n_0 ;
  wire \bdatw[9]_INST_0_i_15_n_0 ;
  wire \bdatw[9]_INST_0_i_23_n_0 ;
  wire \grn_reg[0] ;
  wire \grn_reg[1] ;
  wire \grn_reg[2] ;
  wire \grn_reg[3] ;
  wire \grn_reg[4] ;
  wire \grn_reg[5] ;
  wire \iv[12]_i_51 ;
  wire \iv[12]_i_51_0 ;
  wire \iv[12]_i_51_1 ;
  wire \iv[12]_i_51_2 ;
  wire \iv[15]_i_56 ;
  wire \iv[15]_i_56_0 ;
  wire \iv[15]_i_56_1 ;
  wire \iv[15]_i_56_2 ;
  wire \iv_reg[10] ;
  wire \iv_reg[11] ;
  wire \iv_reg[12] ;
  wire \iv_reg[13] ;
  wire \iv_reg[14] ;
  wire \iv_reg[15] ;
  wire \iv_reg[6] ;
  wire \iv_reg[7] ;
  wire \iv_reg[8] ;
  wire \iv_reg[9] ;
  wire \mul_b_reg[0] ;
  wire \mul_b_reg[0]_0 ;
  wire \mul_b_reg[0]_1 ;
  wire \mul_b_reg[0]_2 ;
  wire \mul_b_reg[10] ;
  wire \mul_b_reg[10]_0 ;
  wire \mul_b_reg[10]_1 ;
  wire \mul_b_reg[10]_2 ;
  wire \mul_b_reg[11] ;
  wire \mul_b_reg[11]_0 ;
  wire \mul_b_reg[11]_1 ;
  wire \mul_b_reg[11]_2 ;
  wire \mul_b_reg[12] ;
  wire \mul_b_reg[12]_0 ;
  wire \mul_b_reg[12]_1 ;
  wire \mul_b_reg[12]_2 ;
  wire \mul_b_reg[13] ;
  wire \mul_b_reg[13]_0 ;
  wire \mul_b_reg[13]_1 ;
  wire \mul_b_reg[13]_2 ;
  wire \mul_b_reg[14] ;
  wire \mul_b_reg[14]_0 ;
  wire \mul_b_reg[14]_1 ;
  wire \mul_b_reg[14]_2 ;
  wire \mul_b_reg[15] ;
  wire \mul_b_reg[15]_0 ;
  wire [15:0]\mul_b_reg[15]_1 ;
  wire \mul_b_reg[15]_2 ;
  wire \mul_b_reg[15]_3 ;
  wire \mul_b_reg[1] ;
  wire \mul_b_reg[1]_0 ;
  wire \mul_b_reg[1]_1 ;
  wire \mul_b_reg[1]_2 ;
  wire \mul_b_reg[1]_3 ;
  wire \mul_b_reg[1]_4 ;
  wire \mul_b_reg[1]_5 ;
  wire \mul_b_reg[1]_6 ;
  wire \mul_b_reg[2] ;
  wire \mul_b_reg[2]_0 ;
  wire \mul_b_reg[2]_1 ;
  wire \mul_b_reg[2]_2 ;
  wire \mul_b_reg[2]_3 ;
  wire \mul_b_reg[2]_4 ;
  wire \mul_b_reg[2]_5 ;
  wire \mul_b_reg[2]_6 ;
  wire \mul_b_reg[3] ;
  wire \mul_b_reg[3]_0 ;
  wire \mul_b_reg[3]_1 ;
  wire \mul_b_reg[3]_2 ;
  wire \mul_b_reg[3]_3 ;
  wire \mul_b_reg[3]_4 ;
  wire \mul_b_reg[3]_5 ;
  wire \mul_b_reg[3]_6 ;
  wire \mul_b_reg[4] ;
  wire \mul_b_reg[4]_0 ;
  wire \mul_b_reg[4]_1 ;
  wire \mul_b_reg[4]_2 ;
  wire \mul_b_reg[4]_3 ;
  wire \mul_b_reg[4]_4 ;
  wire \mul_b_reg[4]_5 ;
  wire \mul_b_reg[4]_6 ;
  wire \mul_b_reg[5] ;
  wire \mul_b_reg[5]_0 ;
  wire \mul_b_reg[5]_1 ;
  wire \mul_b_reg[5]_2 ;
  wire \mul_b_reg[6] ;
  wire \mul_b_reg[6]_0 ;
  wire \mul_b_reg[6]_1 ;
  wire \mul_b_reg[6]_2 ;
  wire \mul_b_reg[7] ;
  wire \mul_b_reg[7]_0 ;
  wire \mul_b_reg[7]_1 ;
  wire \mul_b_reg[7]_2 ;
  wire \mul_b_reg[8] ;
  wire \mul_b_reg[8]_0 ;
  wire \mul_b_reg[8]_1 ;
  wire \mul_b_reg[8]_2 ;
  wire \mul_b_reg[9] ;
  wire \mul_b_reg[9]_0 ;
  wire \mul_b_reg[9]_1 ;
  wire \mul_b_reg[9]_2 ;
  wire [14:0]out;
  wire [30:0]sp_dec_0;
  wire \sp_reg[0] ;
  wire \sp_reg[16] ;
  wire \sp_reg[17] ;
  wire \sp_reg[18] ;
  wire \sp_reg[19] ;
  wire \sp_reg[1] ;
  wire \sp_reg[20] ;
  wire \sp_reg[21] ;
  wire \sp_reg[22] ;
  wire \sp_reg[23] ;
  wire \sp_reg[24] ;
  wire \sp_reg[25] ;
  wire \sp_reg[26] ;
  wire \sp_reg[27] ;
  wire \sp_reg[28] ;
  wire \sp_reg[29] ;
  wire \sp_reg[2] ;
  wire \sp_reg[30] ;
  wire \sp_reg[31] ;
  wire \sp_reg[3] ;
  wire \sp_reg[4] ;
  wire \sp_reg[5] ;
  wire \sp_reg[5]_0 ;
  wire \sr_reg[10] ;
  wire \sr_reg[11] ;
  wire \sr_reg[12] ;
  wire \sr_reg[13] ;
  wire \sr_reg[14] ;
  wire \sr_reg[15] ;
  wire \sr_reg[1] ;
  wire \sr_reg[2] ;
  wire \sr_reg[3] ;
  wire \sr_reg[4] ;
  wire \sr_reg[5] ;
  wire \sr_reg[6] ;
  wire \sr_reg[7] ;
  wire \sr_reg[8] ;
  wire \sr_reg[9] ;
  wire \tr_reg[0] ;
  wire \tr_reg[16] ;
  wire \tr_reg[17] ;
  wire \tr_reg[18] ;
  wire \tr_reg[19] ;
  wire \tr_reg[20] ;
  wire \tr_reg[21] ;
  wire \tr_reg[22] ;
  wire \tr_reg[23] ;
  wire \tr_reg[24] ;
  wire \tr_reg[25] ;
  wire \tr_reg[26] ;
  wire \tr_reg[27] ;
  wire \tr_reg[28] ;
  wire \tr_reg[29] ;
  wire \tr_reg[30] ;
  wire \tr_reg[31] ;
  wire \tr_reg[5] ;

  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[10]_INST_0_i_15 
       (.I0(\bdatw[31]_INST_0_i_1 [2]),
        .I1(bbus_sel_cr[4]),
        .I2(\mul_b_reg[15]_1 [2]),
        .I3(bbus_sel_cr[3]),
        .O(\bdatw[10]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_22 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[9]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [10]),
        .I4(\bdatw[15]_INST_0_i_9_0 [10]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[10]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[10]_INST_0_i_4 
       (.I0(\mul_b_reg[2] ),
        .I1(\mul_b_reg[2]_0 ),
        .I2(\mul_b_reg[2]_1 ),
        .I3(\mul_b_reg[2]_2 ),
        .I4(\bdatw[10]_INST_0_i_15_n_0 ),
        .O(\grn_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[10]_INST_0_i_5 
       (.I0(out[1]),
        .I1(bbus_sel_cr[0]),
        .I2(\mul_b_reg[2]_3 ),
        .I3(\mul_b_reg[2]_4 ),
        .I4(\mul_b_reg[2]_5 ),
        .I5(\mul_b_reg[2]_6 ),
        .O(\sr_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[10]_INST_0_i_6 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[1]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [2]),
        .I4(\bdatw[15]_INST_0_i_9_0 [2]),
        .I5(bbus_sel_cr[1]),
        .O(\sp_reg[2] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[10]_INST_0_i_8 
       (.I0(\mul_b_reg[10] ),
        .I1(\mul_b_reg[10]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [10]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [10]),
        .O(\iv_reg[10] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[10]_INST_0_i_9 
       (.I0(\bdatw[10]_INST_0_i_22_n_0 ),
        .I1(\mul_b_reg[10]_1 ),
        .I2(\mul_b_reg[10]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[9]),
        .O(\sr_reg[10] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[11]_INST_0_i_14 
       (.I0(\bdatw[31]_INST_0_i_1 [3]),
        .I1(bbus_sel_cr[4]),
        .I2(\mul_b_reg[15]_1 [3]),
        .I3(bbus_sel_cr[3]),
        .O(\bdatw[11]_INST_0_i_14_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_22 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[10]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [11]),
        .I4(\bdatw[15]_INST_0_i_9_0 [11]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[11]_INST_0_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[11]_INST_0_i_3 
       (.I0(\mul_b_reg[3] ),
        .I1(\mul_b_reg[3]_0 ),
        .I2(\mul_b_reg[3]_1 ),
        .I3(\mul_b_reg[3]_2 ),
        .I4(\bdatw[11]_INST_0_i_14_n_0 ),
        .O(\grn_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[11]_INST_0_i_4 
       (.I0(out[2]),
        .I1(bbus_sel_cr[0]),
        .I2(\mul_b_reg[3]_3 ),
        .I3(\mul_b_reg[3]_4 ),
        .I4(\mul_b_reg[3]_5 ),
        .I5(\mul_b_reg[3]_6 ),
        .O(\sr_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[11]_INST_0_i_5 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[2]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [3]),
        .I4(\bdatw[15]_INST_0_i_9_0 [3]),
        .I5(bbus_sel_cr[1]),
        .O(\sp_reg[3] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[11]_INST_0_i_8 
       (.I0(\mul_b_reg[11] ),
        .I1(\mul_b_reg[11]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [11]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [11]),
        .O(\iv_reg[11] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[11]_INST_0_i_9 
       (.I0(\bdatw[11]_INST_0_i_22_n_0 ),
        .I1(\mul_b_reg[11]_1 ),
        .I2(\mul_b_reg[11]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[10]),
        .O(\sr_reg[11] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[12]_INST_0_i_10 
       (.I0(\mul_b_reg[12] ),
        .I1(\mul_b_reg[12]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [12]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [12]),
        .O(\iv_reg[12] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[12]_INST_0_i_11 
       (.I0(\bdatw[12]_INST_0_i_26_n_0 ),
        .I1(\mul_b_reg[12]_1 ),
        .I2(\mul_b_reg[12]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[11]),
        .O(\sr_reg[12] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[12]_INST_0_i_16 
       (.I0(\bdatw[31]_INST_0_i_1 [4]),
        .I1(bbus_sel_cr[4]),
        .I2(\mul_b_reg[15]_1 [4]),
        .I3(bbus_sel_cr[3]),
        .O(\bdatw[12]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_26 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[11]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [12]),
        .I4(\bdatw[15]_INST_0_i_9_0 [12]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[12]_INST_0_i_26_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[12]_INST_0_i_5 
       (.I0(\mul_b_reg[4] ),
        .I1(\mul_b_reg[4]_0 ),
        .I2(\mul_b_reg[4]_1 ),
        .I3(\mul_b_reg[4]_2 ),
        .I4(\bdatw[12]_INST_0_i_16_n_0 ),
        .O(\grn_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[12]_INST_0_i_6 
       (.I0(out[3]),
        .I1(bbus_sel_cr[0]),
        .I2(\mul_b_reg[4]_3 ),
        .I3(\mul_b_reg[4]_4 ),
        .I4(\mul_b_reg[4]_5 ),
        .I5(\mul_b_reg[4]_6 ),
        .O(\sr_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[12]_INST_0_i_7 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[3]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [4]),
        .I4(\bdatw[15]_INST_0_i_9_0 [4]),
        .I5(bbus_sel_cr[1]),
        .O(\sp_reg[4] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[13]_INST_0_i_10 
       (.I0(\mul_b_reg[13] ),
        .I1(\mul_b_reg[13]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [13]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [13]),
        .O(\iv_reg[13] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[13]_INST_0_i_11 
       (.I0(\bdatw[13]_INST_0_i_30_n_0 ),
        .I1(\mul_b_reg[13]_1 ),
        .I2(\mul_b_reg[13]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[12]),
        .O(\sr_reg[13] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_21 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[4]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [5]),
        .I4(\bdatw[15]_INST_0_i_9_0 [5]),
        .I5(bbus_sel_cr[1]),
        .O(\sp_reg[5]_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[13]_INST_0_i_30 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[12]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [13]),
        .I4(\bdatw[15]_INST_0_i_9_0 [13]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[13]_INST_0_i_30_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[13]_INST_0_i_5 
       (.I0(\bdatw[31]_INST_0_i_1 [5]),
        .I1(bbus_sel_cr[4]),
        .I2(\mul_b_reg[15]_1 [5]),
        .I3(bbus_sel_cr[3]),
        .O(\tr_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[13]_INST_0_i_8 
       (.I0(\sp_reg[5]_0 ),
        .I1(\mul_b_reg[5] ),
        .I2(\mul_b_reg[5]_0 ),
        .I3(\mul_b_reg[5]_1 ),
        .I4(\mul_b_reg[5]_2 ),
        .I5(bbus_sr[1]),
        .O(\sp_reg[5] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_12 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[5]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [6]),
        .I4(\bdatw[15]_INST_0_i_9_0 [6]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[14]_INST_0_i_12_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[14]_INST_0_i_17 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[13]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [14]),
        .I4(\bdatw[15]_INST_0_i_9_0 [14]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[14]_INST_0_i_17_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[14]_INST_0_i_4 
       (.I0(\mul_b_reg[6] ),
        .I1(\mul_b_reg[6]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [6]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [6]),
        .O(\iv_reg[6] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[14]_INST_0_i_5 
       (.I0(\bdatw[14]_INST_0_i_12_n_0 ),
        .I1(\mul_b_reg[6]_1 ),
        .I2(\mul_b_reg[6]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[5]),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[14]_INST_0_i_7 
       (.I0(\mul_b_reg[14] ),
        .I1(\mul_b_reg[14]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [14]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [14]),
        .O(\iv_reg[14] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[14]_INST_0_i_8 
       (.I0(\bdatw[14]_INST_0_i_17_n_0 ),
        .I1(\mul_b_reg[14]_1 ),
        .I2(\mul_b_reg[14]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[13]),
        .O(\sr_reg[14] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_19 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[6]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [7]),
        .I4(\bdatw[15]_INST_0_i_9_0 [7]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[15]_INST_0_i_19_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[15]_INST_0_i_25 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[14]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [15]),
        .I4(\bdatw[15]_INST_0_i_9_0 [15]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[15]_INST_0_i_25_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[15]_INST_0_i_5 
       (.I0(\mul_b_reg[7] ),
        .I1(\mul_b_reg[7]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [7]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [7]),
        .O(\iv_reg[7] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[15]_INST_0_i_6 
       (.I0(\bdatw[15]_INST_0_i_19_n_0 ),
        .I1(\mul_b_reg[7]_1 ),
        .I2(\mul_b_reg[7]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[6]),
        .O(\sr_reg[7] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[15]_INST_0_i_8 
       (.I0(\mul_b_reg[15] ),
        .I1(\mul_b_reg[15]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [15]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [15]),
        .O(\iv_reg[15] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[15]_INST_0_i_9 
       (.I0(\bdatw[15]_INST_0_i_25_n_0 ),
        .I1(\mul_b_reg[15]_2 ),
        .I2(\mul_b_reg[15]_3 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[14]),
        .O(\sr_reg[15] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[16]_INST_0_i_2 
       (.I0(\bdatw[16]_INST_0_i_1_1 ),
        .I1(\bdatw[16]_INST_0_i_1_2 ),
        .I2(\bdatw[16]_INST_0_i_1_3 ),
        .I3(\bdatw[16]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [16]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[16] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[16]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[15]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [16]),
        .I4(\bdatw[16]_INST_0_i_1 ),
        .I5(\bdatw[16]_INST_0_i_1_0 ),
        .O(\sp_reg[16] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[17]_INST_0_i_2 
       (.I0(\bdatw[17]_INST_0_i_1_1 ),
        .I1(\bdatw[17]_INST_0_i_1_2 ),
        .I2(\bdatw[17]_INST_0_i_1_3 ),
        .I3(\bdatw[17]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [17]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[17] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[17]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[16]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [17]),
        .I4(\bdatw[17]_INST_0_i_1 ),
        .I5(\bdatw[17]_INST_0_i_1_0 ),
        .O(\sp_reg[17] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[18]_INST_0_i_2 
       (.I0(\bdatw[18]_INST_0_i_1_1 ),
        .I1(\bdatw[18]_INST_0_i_1_2 ),
        .I2(\bdatw[18]_INST_0_i_1_3 ),
        .I3(\bdatw[18]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [18]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[18] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[18]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[17]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [18]),
        .I4(\bdatw[18]_INST_0_i_1 ),
        .I5(\bdatw[18]_INST_0_i_1_0 ),
        .O(\sp_reg[18] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[19]_INST_0_i_2 
       (.I0(\bdatw[19]_INST_0_i_1_1 ),
        .I1(\bdatw[19]_INST_0_i_1_2 ),
        .I2(\bdatw[19]_INST_0_i_1_3 ),
        .I3(\bdatw[19]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [19]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[19] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[19]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[18]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [19]),
        .I4(\bdatw[19]_INST_0_i_1 ),
        .I5(\bdatw[19]_INST_0_i_1_0 ),
        .O(\sp_reg[19] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[20]_INST_0_i_2 
       (.I0(\bdatw[20]_INST_0_i_1_1 ),
        .I1(\bdatw[20]_INST_0_i_1_2 ),
        .I2(\bdatw[20]_INST_0_i_1_3 ),
        .I3(\bdatw[20]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [20]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[20] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[20]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[19]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [20]),
        .I4(\bdatw[20]_INST_0_i_1 ),
        .I5(\bdatw[20]_INST_0_i_1_0 ),
        .O(\sp_reg[20] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[21]_INST_0_i_2 
       (.I0(\bdatw[21]_INST_0_i_1_1 ),
        .I1(\bdatw[21]_INST_0_i_1_2 ),
        .I2(\bdatw[21]_INST_0_i_1_3 ),
        .I3(\bdatw[21]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [21]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[21] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[21]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[20]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [21]),
        .I4(\bdatw[21]_INST_0_i_1 ),
        .I5(\bdatw[21]_INST_0_i_1_0 ),
        .O(\sp_reg[21] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[22]_INST_0_i_2 
       (.I0(\bdatw[22]_INST_0_i_1_1 ),
        .I1(\bdatw[22]_INST_0_i_1_2 ),
        .I2(\bdatw[22]_INST_0_i_1_3 ),
        .I3(\bdatw[22]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [22]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[22] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[22]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[21]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [22]),
        .I4(\bdatw[22]_INST_0_i_1 ),
        .I5(\bdatw[22]_INST_0_i_1_0 ),
        .O(\sp_reg[22] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[23]_INST_0_i_2 
       (.I0(\bdatw[23]_INST_0_i_1_1 ),
        .I1(\bdatw[23]_INST_0_i_1_2 ),
        .I2(\bdatw[23]_INST_0_i_1_3 ),
        .I3(\bdatw[23]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [23]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[23]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[22]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [23]),
        .I4(\bdatw[23]_INST_0_i_1 ),
        .I5(\bdatw[23]_INST_0_i_1_0 ),
        .O(\sp_reg[23] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[24]_INST_0_i_2 
       (.I0(\bdatw[24]_INST_0_i_1_1 ),
        .I1(\bdatw[24]_INST_0_i_1_2 ),
        .I2(\bdatw[24]_INST_0_i_1_3 ),
        .I3(\bdatw[24]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [24]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[24]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[23]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [24]),
        .I4(\bdatw[24]_INST_0_i_1 ),
        .I5(\bdatw[24]_INST_0_i_1_0 ),
        .O(\sp_reg[24] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[25]_INST_0_i_2 
       (.I0(\bdatw[25]_INST_0_i_1_1 ),
        .I1(\bdatw[25]_INST_0_i_1_2 ),
        .I2(\bdatw[25]_INST_0_i_1_3 ),
        .I3(\bdatw[25]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [25]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[25] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[25]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[24]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [25]),
        .I4(\bdatw[25]_INST_0_i_1 ),
        .I5(\bdatw[25]_INST_0_i_1_0 ),
        .O(\sp_reg[25] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[26]_INST_0_i_2 
       (.I0(\bdatw[26]_INST_0_i_1_1 ),
        .I1(\bdatw[26]_INST_0_i_1_2 ),
        .I2(\bdatw[26]_INST_0_i_1_3 ),
        .I3(\bdatw[26]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [26]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[26]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[25]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [26]),
        .I4(\bdatw[26]_INST_0_i_1 ),
        .I5(\bdatw[26]_INST_0_i_1_0 ),
        .O(\sp_reg[26] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[27]_INST_0_i_2 
       (.I0(\bdatw[27]_INST_0_i_1_1 ),
        .I1(\bdatw[27]_INST_0_i_1_2 ),
        .I2(\bdatw[27]_INST_0_i_1_3 ),
        .I3(\bdatw[27]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [27]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[27] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[27]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[26]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [27]),
        .I4(\bdatw[27]_INST_0_i_1 ),
        .I5(\bdatw[27]_INST_0_i_1_0 ),
        .O(\sp_reg[27] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[28]_INST_0_i_2 
       (.I0(\bdatw[28]_INST_0_i_1_1 ),
        .I1(\bdatw[28]_INST_0_i_1_2 ),
        .I2(\bdatw[28]_INST_0_i_1_3 ),
        .I3(\bdatw[28]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [28]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[28] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[28]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[27]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [28]),
        .I4(\bdatw[28]_INST_0_i_1 ),
        .I5(\bdatw[28]_INST_0_i_1_0 ),
        .O(\sp_reg[28] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[29]_INST_0_i_2 
       (.I0(\bdatw[29]_INST_0_i_1_1 ),
        .I1(\bdatw[29]_INST_0_i_1_2 ),
        .I2(\bdatw[29]_INST_0_i_1_3 ),
        .I3(\bdatw[29]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [29]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[29] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[29]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[28]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [29]),
        .I4(\bdatw[29]_INST_0_i_1 ),
        .I5(\bdatw[29]_INST_0_i_1_0 ),
        .O(\sp_reg[29] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[30]_INST_0_i_2 
       (.I0(\bdatw[30]_INST_0_i_1_1 ),
        .I1(\bdatw[30]_INST_0_i_1_2 ),
        .I2(\bdatw[30]_INST_0_i_1_3 ),
        .I3(\bdatw[30]_INST_0_i_1_4 ),
        .I4(\bdatw[31]_INST_0_i_1 [30]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[30]_INST_0_i_3 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[29]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [30]),
        .I4(\bdatw[30]_INST_0_i_1 ),
        .I5(\bdatw[30]_INST_0_i_1_0 ),
        .O(\sp_reg[30] ));
  LUT6 #(
    .INIT(64'hFFFFFFFEFFFEFFFE)) 
    \bdatw[31]_INST_0_i_4 
       (.I0(\bdatw[31]_INST_0_i_1_3 ),
        .I1(\bdatw[31]_INST_0_i_1_4 ),
        .I2(\bdatw[31]_INST_0_i_1_5 ),
        .I3(\bdatw[31]_INST_0_i_1_6 ),
        .I4(\bdatw[31]_INST_0_i_1 [31]),
        .I5(bbus_sel_cr[4]),
        .O(\tr_reg[31] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFF888)) 
    \bdatw[31]_INST_0_i_5 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[30]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [31]),
        .I4(\bdatw[31]_INST_0_i_1_1 ),
        .I5(\bdatw[31]_INST_0_i_1_2 ),
        .O(\sp_reg[31] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[8]_INST_0_i_10 
       (.I0(\mul_b_reg[8] ),
        .I1(\mul_b_reg[8]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [8]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [8]),
        .O(\iv_reg[8] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[8]_INST_0_i_11 
       (.I0(\bdatw[8]_INST_0_i_24_n_0 ),
        .I1(\mul_b_reg[8]_1 ),
        .I2(\mul_b_reg[8]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[7]),
        .O(\sr_reg[8] ));
  LUT5 #(
    .INIT(32'hFFC8C8C8)) 
    \bdatw[8]_INST_0_i_16 
       (.I0(bbus_sel_cr[5]),
        .I1(\bdatw[31]_INST_0_i_1_0 [0]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[15]_INST_0_i_9_0 [0]),
        .I4(bbus_sel_cr[1]),
        .O(\bdatw[8]_INST_0_i_16_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[8]_INST_0_i_24 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[7]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [8]),
        .I4(\bdatw[15]_INST_0_i_9_0 [8]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[8]_INST_0_i_24_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[8]_INST_0_i_5 
       (.I0(\bdatw[31]_INST_0_i_1 [0]),
        .I1(bbus_sel_cr[4]),
        .I2(\mul_b_reg[15]_1 [0]),
        .I3(bbus_sel_cr[3]),
        .O(\tr_reg[0] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \bdatw[8]_INST_0_i_8 
       (.I0(\bdatw[8]_INST_0_i_16_n_0 ),
        .I1(\mul_b_reg[0] ),
        .I2(\mul_b_reg[0]_0 ),
        .I3(\mul_b_reg[0]_1 ),
        .I4(\mul_b_reg[0]_2 ),
        .I5(bbus_sr[0]),
        .O(\sp_reg[0] ));
  LUT4 #(
    .INIT(16'hF888)) 
    \bdatw[9]_INST_0_i_15 
       (.I0(\bdatw[31]_INST_0_i_1 [1]),
        .I1(bbus_sel_cr[4]),
        .I2(\mul_b_reg[15]_1 [1]),
        .I3(bbus_sel_cr[3]),
        .O(\bdatw[9]_INST_0_i_15_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_23 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[8]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [9]),
        .I4(\bdatw[15]_INST_0_i_9_0 [9]),
        .I5(bbus_sel_cr[1]),
        .O(\bdatw[9]_INST_0_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \bdatw[9]_INST_0_i_4 
       (.I0(\mul_b_reg[1] ),
        .I1(\mul_b_reg[1]_0 ),
        .I2(\mul_b_reg[1]_1 ),
        .I3(\mul_b_reg[1]_2 ),
        .I4(\bdatw[9]_INST_0_i_15_n_0 ),
        .O(\grn_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \bdatw[9]_INST_0_i_5 
       (.I0(out[0]),
        .I1(bbus_sel_cr[0]),
        .I2(\mul_b_reg[1]_3 ),
        .I3(\mul_b_reg[1]_4 ),
        .I4(\mul_b_reg[1]_5 ),
        .I5(\mul_b_reg[1]_6 ),
        .O(\sr_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFF888F888F888)) 
    \bdatw[9]_INST_0_i_6 
       (.I0(bbus_sel_cr[5]),
        .I1(sp_dec_0[0]),
        .I2(bbus_sel_cr[2]),
        .I3(\bdatw[31]_INST_0_i_1_0 [1]),
        .I4(\bdatw[15]_INST_0_i_9_0 [1]),
        .I5(bbus_sel_cr[1]),
        .O(\sp_reg[1] ));
  LUT6 #(
    .INIT(64'hFFFFFEEEFEEEFEEE)) 
    \bdatw[9]_INST_0_i_8 
       (.I0(\mul_b_reg[9] ),
        .I1(\mul_b_reg[9]_0 ),
        .I2(bbus_sel_cr[3]),
        .I3(\mul_b_reg[15]_1 [9]),
        .I4(bbus_sel_cr[4]),
        .I5(\bdatw[31]_INST_0_i_1 [9]),
        .O(\iv_reg[9] ));
  LUT5 #(
    .INIT(32'hFFFEFEFE)) 
    \bdatw[9]_INST_0_i_9 
       (.I0(\bdatw[9]_INST_0_i_23_n_0 ),
        .I1(\mul_b_reg[9]_1 ),
        .I2(\mul_b_reg[9]_2 ),
        .I3(bbus_sel_cr[0]),
        .I4(out[8]),
        .O(\sr_reg[9] ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFF8)) 
    \iv[15]_i_98 
       (.I0(out[4]),
        .I1(bbus_sel_cr[0]),
        .I2(\mul_b_reg[5]_2 ),
        .I3(\mul_b_reg[5]_1 ),
        .I4(\mul_b_reg[5]_0 ),
        .I5(\mul_b_reg[5] ),
        .O(\sr_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \iv[15]_i_99 
       (.I0(\iv[15]_i_56 ),
        .I1(\iv[15]_i_56_0 ),
        .I2(\iv[15]_i_56_1 ),
        .I3(\iv[15]_i_56_2 ),
        .I4(\tr_reg[5] ),
        .O(\grn_reg[5] ));
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \sr[7]_i_54 
       (.I0(\iv[12]_i_51 ),
        .I1(\iv[12]_i_51_0 ),
        .I2(\iv[12]_i_51_1 ),
        .I3(\iv[12]_i_51_2 ),
        .I4(\tr_reg[0] ),
        .O(\grn_reg[0] ));
endmodule

module niho_rgf_ctl
   (bank_sel,
    out);
  output [0:0]bank_sel;
  input [2:0]out;

  wire [0:0]bank_sel;
  wire [2:0]out;

  LUT3 #(
    .INIT(8'h45)) 
    bank_sel__0
       (.I0(out[0]),
        .I1(out[2]),
        .I2(out[1]),
        .O(bank_sel));
endmodule

module niho_rgf_grn
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_10
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_11
   (Q,
    SR,
    \grn_reg[0]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_12
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_13
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_14
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_15
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_16
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_17
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_18
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_19
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_20
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_21
   (SR,
    Q,
    rst_n,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [0:0]SR;
  output [15:0]Q;
  input rst_n;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire rst_n;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT1 #(
    .INIT(2'h1)) 
    \sr[11]_i_1 
       (.I0(rst_n),
        .O(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_27
   (Q,
    SR,
    E,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]E;
  input [15:0]cbus;
  input clk;

  wire [0:0]E;
  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(E),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(E),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(E),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(E),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(E),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(E),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(E),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(E),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(E),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(E),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(E),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(E),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(E),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(E),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(E),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(E),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_28
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_29
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_30
   (Q,
    SR,
    \grn_reg[0]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_31
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_32
   (Q,
    SR,
    \grn_reg[0]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_33
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_34
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_35
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_36
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_37
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_38
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_39
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_40
   (Q,
    SR,
    \grn_reg[0]_0 ,
    \grn_reg[15]_0 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[0]_0 ;
  input [15:0]\grn_reg[15]_0 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[0]_0 ;
  wire [15:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[0]_0 ),
        .D(\grn_reg[15]_0 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_41
   (Q,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_42
   (\bdatw[8]_INST_0_i_2 ,
    \iv[7]_i_33 ,
    \sr_reg[8] ,
    \sr[7]_i_20 ,
    \sr_reg[8]_0 ,
    \sr_reg[8]_1 ,
    \sr_reg[8]_2 ,
    \iv[1]_i_15 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \iv[2]_i_15 ,
    \iv[2]_i_26 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    \sr_reg[8]_12 ,
    \iv[5]_i_28 ,
    \sr_reg[8]_13 ,
    \iv[4]_i_29 ,
    \sr_reg[8]_14 ,
    \sr_reg[8]_15 ,
    \sr_reg[8]_16 ,
    \sr_reg[8]_17 ,
    \iv[9]_i_36 ,
    \iv[7]_i_17 ,
    \iv[15]_i_94 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \iv[10]_i_10 ,
    \iv[9]_i_11 ,
    \sr_reg[8]_22 ,
    \bdatw[12]_INST_0_i_1 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \sr_reg[8]_28 ,
    \bdatw[12]_INST_0_i_1_0 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \sr_reg[8]_33 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \sr_reg[8]_36 ,
    \iv[7]_i_25 ,
    \sr_reg[8]_37 ,
    \iv[0]_i_25 ,
    \sr_reg[8]_38 ,
    \sr_reg[8]_39 ,
    \sr_reg[6] ,
    \iv[14]_i_49 ,
    \sr_reg[8]_40 ,
    \sr_reg[8]_41 ,
    \iv[5]_i_23 ,
    \sr_reg[8]_42 ,
    \sr_reg[8]_43 ,
    \sr_reg[8]_44 ,
    \sr_reg[8]_45 ,
    \badr[5]_INST_0_i_1 ,
    \niho_dsp_a[15]_INST_0_i_3 ,
    \sr_reg[8]_46 ,
    \sr_reg[6]_0 ,
    \sr_reg[6]_1 ,
    \sr_reg[6]_2 ,
    \sr_reg[6]_3 ,
    \sr_reg[8]_47 ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    \sr_reg[8]_50 ,
    Q,
    \iv[8]_i_9 ,
    \iv[0]_i_7 ,
    \sr[4]_i_146 ,
    \sr[4]_i_82 ,
    \iv[0]_i_7_0 ,
    bbus_0,
    \iv[9]_i_4_0 ,
    \iv[7]_i_7 ,
    \iv[7]_i_7_0 ,
    DI,
    \iv[7]_i_7_1 ,
    \iv[7]_i_7_2 ,
    \niho_dsp_a[32] ,
    \iv[5]_i_7 ,
    \iv[7]_i_9_0 ,
    \iv[9]_i_4_1 ,
    \iv[7]_i_9_1 ,
    \iv[11]_i_2 ,
    \iv[8]_i_5_0 ,
    \iv[11]_i_5_0 ,
    \iv[11]_i_5_1 ,
    \tr_reg[1] ,
    \tr_reg[1]_0 ,
    \iv[1]_i_3_0 ,
    \iv[2]_i_3_0 ,
    \sr[4]_i_47 ,
    \sr[4]_i_47_0 ,
    \iv[3]_i_3 ,
    \sr[4]_i_46 ,
    \sr[4]_i_46_0 ,
    \sr[4]_i_46_1 ,
    \iv[13]_i_2 ,
    \iv[13]_i_2_0 ,
    \iv[12]_i_2 ,
    \iv[12]_i_2_0 ,
    \iv[10]_i_2 ,
    \iv[10]_i_2_0 ,
    \iv[5]_i_3 ,
    \sr[4]_i_33 ,
    \sr[4]_i_33_0 ,
    \sr[4]_i_33_1 ,
    \iv[4]_i_3 ,
    \sr[4]_i_31 ,
    \sr[4]_i_31_0 ,
    \iv[8]_i_2 ,
    \iv[8]_i_5_1 ,
    \iv[8]_i_5_2 ,
    \iv[8]_i_2_0 ,
    \iv[14]_i_2 ,
    \iv[14]_i_5_0 ,
    \iv[14]_i_5_1 ,
    \iv[9]_i_2 ,
    \iv[9]_i_5_0 ,
    \iv[9]_i_5_1 ,
    \iv[9]_i_2_0 ,
    \iv[7]_i_3 ,
    \iv[9]_i_4_2 ,
    \iv[9]_i_4_3 ,
    \sr[4]_i_19 ,
    \sr[4]_i_21 ,
    \iv[10]_i_2_1 ,
    \iv[10]_i_2_2 ,
    \iv[9]_i_2_1 ,
    \iv[1]_i_9_0 ,
    \iv[1]_i_9_1 ,
    \iv[13]_i_5_0 ,
    \iv[13]_i_5_1 ,
    \iv[12]_i_5_0 ,
    \iv[12]_i_5_1 ,
    \iv[10]_i_5_0 ,
    \iv[10]_i_5_1 ,
    \iv[1]_i_10_0 ,
    \iv[1]_i_10_1 ,
    \iv[1]_i_10_2 ,
    \iv[3]_i_3_0 ,
    \iv[3]_i_10_0 ,
    \iv[3]_i_10_1 ,
    \iv[3]_i_10_2 ,
    \iv[4]_i_14 ,
    \iv[4]_i_14_0 ,
    \iv[5]_i_10_0 ,
    \iv[13]_i_6 ,
    \iv[3]_i_15 ,
    \iv[4]_i_10_0 ,
    \iv[12]_i_6 ,
    \iv[1]_i_15_0 ,
    \iv[2]_i_10_0 ,
    \iv[10]_i_6 ,
    \iv[5]_i_3_0 ,
    \iv[6]_i_10 ,
    \iv[6]_i_10_0 ,
    \iv[6]_i_10_1 ,
    \iv[6]_i_9 ,
    \iv[7]_i_9_2 ,
    \iv[7]_i_9_3 ,
    \iv[11]_i_5_2 ,
    \iv[11]_i_5_3 ,
    \iv[11]_i_5_4 ,
    \iv[1]_i_9_2 ,
    \iv[1]_i_9_3 ,
    \iv[1]_i_9_4 ,
    \iv[2]_i_9_0 ,
    \iv[2]_i_9_1 ,
    \iv[2]_i_9_2 ,
    \iv[3]_i_9_0 ,
    \iv[3]_i_9_1 ,
    \iv[3]_i_9_2 ,
    \iv[13]_i_5_2 ,
    \iv[13]_i_5_3 ,
    \iv[13]_i_5_4 ,
    \iv[12]_i_5_2 ,
    \iv[12]_i_5_3 ,
    \iv[12]_i_5_4 ,
    \iv[10]_i_5_2 ,
    \iv[10]_i_5_3 ,
    \iv[10]_i_5_4 ,
    \iv[5]_i_9_0 ,
    \iv[5]_i_9_1 ,
    \iv[5]_i_9_2 ,
    \iv[4]_i_9_0 ,
    \iv[4]_i_9_1 ,
    \iv[4]_i_9_2 ,
    \iv[8]_i_5_3 ,
    \iv[8]_i_5_4 ,
    \iv[8]_i_5_5 ,
    \iv[14]_i_5_2 ,
    \iv[14]_i_5_3 ,
    \iv[14]_i_5_4 ,
    \iv[9]_i_5_2 ,
    \iv[9]_i_5_3 ,
    \iv[9]_i_5_4 ,
    \iv[6]_i_9_0 ,
    \iv[6]_i_9_1 ,
    \iv[6]_i_9_2 ,
    \iv[4]_i_10_1 ,
    \sr[4]_i_31_1 ,
    \iv[4]_i_17_0 ,
    \iv[11]_i_6_0 ,
    \iv[1]_i_10_3 ,
    \iv[7]_i_3_0 ,
    \iv[7]_i_9_4 ,
    \iv[7]_i_3_1 ,
    \iv[12]_i_9 ,
    \iv[8]_i_6_0 ,
    \iv[8]_i_6_1 ,
    \iv[3]_i_20 ,
    \iv[12]_i_15 ,
    \iv[8]_i_10 ,
    \iv[8]_i_10_0 ,
    \iv[12]_i_21 ,
    \iv[12]_i_21_0 ,
    \iv[12]_i_21_1 ,
    \tr[25]_i_7 ,
    \iv[1]_i_20_0 ,
    \iv[13]_i_15 ,
    \tr[25]_i_7_0 ,
    \sr[4]_i_135 ,
    \sr[4]_i_135_0 ,
    \iv[6]_i_15 ,
    \iv[6]_i_15_0 ,
    \sr[4]_i_135_1 ,
    \sr[4]_i_135_2 ,
    \iv[5]_i_10_1 ,
    \iv[5]_i_14 ,
    \tr[17]_i_9 ,
    \iv[11]_i_18 ,
    \iv[1]_i_32 ,
    \iv[1]_i_23_0 ,
    \iv[1]_i_23_1 ,
    \iv[7]_i_17_0 ,
    \sr[4]_i_88 ,
    \sr[4]_i_88_0 ,
    \iv[7]_i_17_1 ,
    \sr[4]_i_146_0 ,
    \sr[4]_i_114 ,
    \sr[4]_i_114_0 ,
    \iv[0]_i_7_1 ,
    \iv[14]_i_19 ,
    \niho_dsp_a[32]_0 ,
    \niho_dsp_a[32]_1 ,
    p_0_in,
    p_1_in,
    \niho_dsp_a[32]_2 ,
    \tr[23]_i_10 ,
    \iv[4]_i_10_2 ,
    \iv[5]_i_10_2 ,
    \iv[2]_i_15_0 ,
    \iv[2]_i_10_1 ,
    \iv[11]_i_18_0 ,
    \sr[4]_i_146_1 ,
    \iv[3]_i_15_0 ,
    \iv[9]_i_11_0 ,
    \iv[14]_i_6 ,
    \iv[2]_i_15_1 ,
    \iv[2]_i_15_2 ,
    \iv[13]_i_15_0 ,
    \iv[4]_i_14_1 ,
    \iv[12]_i_15_0 ,
    SR,
    \grn_reg[15]_0 ,
    \grn_reg[15]_1 ,
    clk);
  output \bdatw[8]_INST_0_i_2 ;
  output \iv[7]_i_33 ;
  output \sr_reg[8] ;
  output \sr[7]_i_20 ;
  output \sr_reg[8]_0 ;
  output \sr_reg[8]_1 ;
  output \sr_reg[8]_2 ;
  output \iv[1]_i_15 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \iv[2]_i_15 ;
  output \iv[2]_i_26 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output \sr_reg[8]_12 ;
  output \iv[5]_i_28 ;
  output \sr_reg[8]_13 ;
  output \iv[4]_i_29 ;
  output \sr_reg[8]_14 ;
  output \sr_reg[8]_15 ;
  output \sr_reg[8]_16 ;
  output \sr_reg[8]_17 ;
  output \iv[9]_i_36 ;
  output \iv[7]_i_17 ;
  output \iv[15]_i_94 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \iv[10]_i_10 ;
  output \iv[9]_i_11 ;
  output \sr_reg[8]_22 ;
  output \bdatw[12]_INST_0_i_1 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \sr_reg[8]_28 ;
  output \bdatw[12]_INST_0_i_1_0 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \sr_reg[8]_33 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \sr_reg[8]_36 ;
  output \iv[7]_i_25 ;
  output \sr_reg[8]_37 ;
  output \iv[0]_i_25 ;
  output \sr_reg[8]_38 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[6] ;
  output \iv[14]_i_49 ;
  output \sr_reg[8]_40 ;
  output \sr_reg[8]_41 ;
  output \iv[5]_i_23 ;
  output \sr_reg[8]_42 ;
  output \sr_reg[8]_43 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[8]_45 ;
  output \badr[5]_INST_0_i_1 ;
  output \niho_dsp_a[15]_INST_0_i_3 ;
  output \sr_reg[8]_46 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[6]_1 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[8]_47 ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output \sr_reg[8]_50 ;
  output [15:0]Q;
  input \iv[8]_i_9 ;
  input \iv[0]_i_7 ;
  input \sr[4]_i_146 ;
  input \sr[4]_i_82 ;
  input [0:0]\iv[0]_i_7_0 ;
  input [1:0]bbus_0;
  input \iv[9]_i_4_0 ;
  input [1:0]\iv[7]_i_7 ;
  input \iv[7]_i_7_0 ;
  input [1:0]DI;
  input \iv[7]_i_7_1 ;
  input \iv[7]_i_7_2 ;
  input [1:0]\niho_dsp_a[32] ;
  input \iv[5]_i_7 ;
  input \iv[7]_i_9_0 ;
  input \iv[9]_i_4_1 ;
  input \iv[7]_i_9_1 ;
  input \iv[11]_i_2 ;
  input \iv[8]_i_5_0 ;
  input \iv[11]_i_5_0 ;
  input \iv[11]_i_5_1 ;
  input \tr_reg[1] ;
  input \tr_reg[1]_0 ;
  input \iv[1]_i_3_0 ;
  input \iv[2]_i_3_0 ;
  input \sr[4]_i_47 ;
  input \sr[4]_i_47_0 ;
  input \iv[3]_i_3 ;
  input \sr[4]_i_46 ;
  input \sr[4]_i_46_0 ;
  input \sr[4]_i_46_1 ;
  input \iv[13]_i_2 ;
  input \iv[13]_i_2_0 ;
  input \iv[12]_i_2 ;
  input \iv[12]_i_2_0 ;
  input \iv[10]_i_2 ;
  input \iv[10]_i_2_0 ;
  input \iv[5]_i_3 ;
  input \sr[4]_i_33 ;
  input \sr[4]_i_33_0 ;
  input \sr[4]_i_33_1 ;
  input \iv[4]_i_3 ;
  input \sr[4]_i_31 ;
  input \sr[4]_i_31_0 ;
  input \iv[8]_i_2 ;
  input \iv[8]_i_5_1 ;
  input \iv[8]_i_5_2 ;
  input \iv[8]_i_2_0 ;
  input \iv[14]_i_2 ;
  input \iv[14]_i_5_0 ;
  input \iv[14]_i_5_1 ;
  input \iv[9]_i_2 ;
  input \iv[9]_i_5_0 ;
  input \iv[9]_i_5_1 ;
  input \iv[9]_i_2_0 ;
  input \iv[7]_i_3 ;
  input \iv[9]_i_4_2 ;
  input \iv[9]_i_4_3 ;
  input \sr[4]_i_19 ;
  input \sr[4]_i_21 ;
  input \iv[10]_i_2_1 ;
  input \iv[10]_i_2_2 ;
  input \iv[9]_i_2_1 ;
  input \iv[1]_i_9_0 ;
  input \iv[1]_i_9_1 ;
  input \iv[13]_i_5_0 ;
  input \iv[13]_i_5_1 ;
  input \iv[12]_i_5_0 ;
  input \iv[12]_i_5_1 ;
  input \iv[10]_i_5_0 ;
  input \iv[10]_i_5_1 ;
  input \iv[1]_i_10_0 ;
  input \iv[1]_i_10_1 ;
  input \iv[1]_i_10_2 ;
  input \iv[3]_i_3_0 ;
  input \iv[3]_i_10_0 ;
  input \iv[3]_i_10_1 ;
  input \iv[3]_i_10_2 ;
  input \iv[4]_i_14 ;
  input \iv[4]_i_14_0 ;
  input \iv[5]_i_10_0 ;
  input \iv[13]_i_6 ;
  input \iv[3]_i_15 ;
  input \iv[4]_i_10_0 ;
  input \iv[12]_i_6 ;
  input \iv[1]_i_15_0 ;
  input \iv[2]_i_10_0 ;
  input \iv[10]_i_6 ;
  input \iv[5]_i_3_0 ;
  input \iv[6]_i_10 ;
  input \iv[6]_i_10_0 ;
  input \iv[6]_i_10_1 ;
  input \iv[6]_i_9 ;
  input \iv[7]_i_9_2 ;
  input \iv[7]_i_9_3 ;
  input \iv[11]_i_5_2 ;
  input \iv[11]_i_5_3 ;
  input \iv[11]_i_5_4 ;
  input \iv[1]_i_9_2 ;
  input \iv[1]_i_9_3 ;
  input \iv[1]_i_9_4 ;
  input \iv[2]_i_9_0 ;
  input \iv[2]_i_9_1 ;
  input \iv[2]_i_9_2 ;
  input \iv[3]_i_9_0 ;
  input \iv[3]_i_9_1 ;
  input \iv[3]_i_9_2 ;
  input \iv[13]_i_5_2 ;
  input \iv[13]_i_5_3 ;
  input \iv[13]_i_5_4 ;
  input \iv[12]_i_5_2 ;
  input \iv[12]_i_5_3 ;
  input \iv[12]_i_5_4 ;
  input \iv[10]_i_5_2 ;
  input \iv[10]_i_5_3 ;
  input \iv[10]_i_5_4 ;
  input \iv[5]_i_9_0 ;
  input \iv[5]_i_9_1 ;
  input \iv[5]_i_9_2 ;
  input \iv[4]_i_9_0 ;
  input \iv[4]_i_9_1 ;
  input \iv[4]_i_9_2 ;
  input \iv[8]_i_5_3 ;
  input \iv[8]_i_5_4 ;
  input \iv[8]_i_5_5 ;
  input \iv[14]_i_5_2 ;
  input \iv[14]_i_5_3 ;
  input \iv[14]_i_5_4 ;
  input \iv[9]_i_5_2 ;
  input \iv[9]_i_5_3 ;
  input \iv[9]_i_5_4 ;
  input \iv[6]_i_9_0 ;
  input \iv[6]_i_9_1 ;
  input \iv[6]_i_9_2 ;
  input \iv[4]_i_10_1 ;
  input \sr[4]_i_31_1 ;
  input \iv[4]_i_17_0 ;
  input \iv[11]_i_6_0 ;
  input \iv[1]_i_10_3 ;
  input \iv[7]_i_3_0 ;
  input \iv[7]_i_9_4 ;
  input \iv[7]_i_3_1 ;
  input \iv[12]_i_9 ;
  input \iv[8]_i_6_0 ;
  input \iv[8]_i_6_1 ;
  input \iv[3]_i_20 ;
  input \iv[12]_i_15 ;
  input \iv[8]_i_10 ;
  input \iv[8]_i_10_0 ;
  input \iv[12]_i_21 ;
  input \iv[12]_i_21_0 ;
  input \iv[12]_i_21_1 ;
  input \tr[25]_i_7 ;
  input \iv[1]_i_20_0 ;
  input \iv[13]_i_15 ;
  input \tr[25]_i_7_0 ;
  input \sr[4]_i_135 ;
  input \sr[4]_i_135_0 ;
  input \iv[6]_i_15 ;
  input \iv[6]_i_15_0 ;
  input \sr[4]_i_135_1 ;
  input \sr[4]_i_135_2 ;
  input \iv[5]_i_10_1 ;
  input \iv[5]_i_14 ;
  input \tr[17]_i_9 ;
  input \iv[11]_i_18 ;
  input \iv[1]_i_32 ;
  input \iv[1]_i_23_0 ;
  input \iv[1]_i_23_1 ;
  input \iv[7]_i_17_0 ;
  input \sr[4]_i_88 ;
  input \sr[4]_i_88_0 ;
  input \iv[7]_i_17_1 ;
  input \sr[4]_i_146_0 ;
  input \sr[4]_i_114 ;
  input \sr[4]_i_114_0 ;
  input \iv[0]_i_7_1 ;
  input [0:0]\iv[14]_i_19 ;
  input \niho_dsp_a[32]_0 ;
  input \niho_dsp_a[32]_1 ;
  input [0:0]p_0_in;
  input [0:0]p_1_in;
  input \niho_dsp_a[32]_2 ;
  input \tr[23]_i_10 ;
  input \iv[4]_i_10_2 ;
  input \iv[5]_i_10_2 ;
  input \iv[2]_i_15_0 ;
  input \iv[2]_i_10_1 ;
  input \iv[11]_i_18_0 ;
  input \sr[4]_i_146_1 ;
  input \iv[3]_i_15_0 ;
  input \iv[9]_i_11_0 ;
  input \iv[14]_i_6 ;
  input \iv[2]_i_15_1 ;
  input \iv[2]_i_15_2 ;
  input \iv[13]_i_15_0 ;
  input \iv[4]_i_14_1 ;
  input \iv[12]_i_15_0 ;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]\grn_reg[15]_1 ;
  input clk;

  wire [1:0]DI;
  wire [15:0]Q;
  wire [0:0]SR;
  wire \badr[5]_INST_0_i_1 ;
  wire [1:0]bbus_0;
  wire \bdatw[12]_INST_0_i_1 ;
  wire \bdatw[12]_INST_0_i_1_0 ;
  wire \bdatw[8]_INST_0_i_2 ;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;
  wire [15:0]\grn_reg[15]_1 ;
  wire \iv[0]_i_25 ;
  wire \iv[0]_i_7 ;
  wire [0:0]\iv[0]_i_7_0 ;
  wire \iv[0]_i_7_1 ;
  wire \iv[10]_i_10 ;
  wire \iv[10]_i_12_n_0 ;
  wire \iv[10]_i_14_n_0 ;
  wire \iv[10]_i_2 ;
  wire \iv[10]_i_2_0 ;
  wire \iv[10]_i_2_1 ;
  wire \iv[10]_i_2_2 ;
  wire \iv[10]_i_5_0 ;
  wire \iv[10]_i_5_1 ;
  wire \iv[10]_i_5_2 ;
  wire \iv[10]_i_5_3 ;
  wire \iv[10]_i_5_4 ;
  wire \iv[10]_i_6 ;
  wire \iv[11]_i_12_n_0 ;
  wire \iv[11]_i_14_n_0 ;
  wire \iv[11]_i_16_n_0 ;
  wire \iv[11]_i_18 ;
  wire \iv[11]_i_18_0 ;
  wire \iv[11]_i_2 ;
  wire \iv[11]_i_5_0 ;
  wire \iv[11]_i_5_1 ;
  wire \iv[11]_i_5_2 ;
  wire \iv[11]_i_5_3 ;
  wire \iv[11]_i_5_4 ;
  wire \iv[11]_i_6_0 ;
  wire \iv[12]_i_11_n_0 ;
  wire \iv[12]_i_14_n_0 ;
  wire \iv[12]_i_15 ;
  wire \iv[12]_i_15_0 ;
  wire \iv[12]_i_2 ;
  wire \iv[12]_i_21 ;
  wire \iv[12]_i_21_0 ;
  wire \iv[12]_i_21_1 ;
  wire \iv[12]_i_2_0 ;
  wire \iv[12]_i_5_0 ;
  wire \iv[12]_i_5_1 ;
  wire \iv[12]_i_5_2 ;
  wire \iv[12]_i_5_3 ;
  wire \iv[12]_i_5_4 ;
  wire \iv[12]_i_6 ;
  wire \iv[12]_i_9 ;
  wire \iv[13]_i_11_n_0 ;
  wire \iv[13]_i_14_n_0 ;
  wire \iv[13]_i_15 ;
  wire \iv[13]_i_15_0 ;
  wire \iv[13]_i_2 ;
  wire \iv[13]_i_2_0 ;
  wire \iv[13]_i_5_0 ;
  wire \iv[13]_i_5_1 ;
  wire \iv[13]_i_5_2 ;
  wire \iv[13]_i_5_3 ;
  wire \iv[13]_i_5_4 ;
  wire \iv[13]_i_6 ;
  wire \iv[14]_i_12_n_0 ;
  wire \iv[14]_i_14_n_0 ;
  wire [0:0]\iv[14]_i_19 ;
  wire \iv[14]_i_2 ;
  wire \iv[14]_i_49 ;
  wire \iv[14]_i_5_0 ;
  wire \iv[14]_i_5_1 ;
  wire \iv[14]_i_5_2 ;
  wire \iv[14]_i_5_3 ;
  wire \iv[14]_i_5_4 ;
  wire \iv[14]_i_6 ;
  wire \iv[15]_i_94 ;
  wire \iv[1]_i_10_0 ;
  wire \iv[1]_i_10_1 ;
  wire \iv[1]_i_10_2 ;
  wire \iv[1]_i_10_3 ;
  wire \iv[1]_i_10_n_0 ;
  wire \iv[1]_i_14_n_0 ;
  wire \iv[1]_i_15 ;
  wire \iv[1]_i_15_0 ;
  wire \iv[1]_i_17_n_0 ;
  wire \iv[1]_i_19_n_0 ;
  wire \iv[1]_i_20_0 ;
  wire \iv[1]_i_20_n_0 ;
  wire \iv[1]_i_21_n_0 ;
  wire \iv[1]_i_23_0 ;
  wire \iv[1]_i_23_1 ;
  wire \iv[1]_i_31_n_0 ;
  wire \iv[1]_i_32 ;
  wire \iv[1]_i_3_0 ;
  wire \iv[1]_i_9_0 ;
  wire \iv[1]_i_9_1 ;
  wire \iv[1]_i_9_2 ;
  wire \iv[1]_i_9_3 ;
  wire \iv[1]_i_9_4 ;
  wire \iv[1]_i_9_n_0 ;
  wire \iv[2]_i_10_0 ;
  wire \iv[2]_i_10_1 ;
  wire \iv[2]_i_10_n_0 ;
  wire \iv[2]_i_14_n_0 ;
  wire \iv[2]_i_15 ;
  wire \iv[2]_i_15_0 ;
  wire \iv[2]_i_15_1 ;
  wire \iv[2]_i_15_2 ;
  wire \iv[2]_i_18_n_0 ;
  wire \iv[2]_i_20_n_0 ;
  wire \iv[2]_i_25_n_0 ;
  wire \iv[2]_i_26 ;
  wire \iv[2]_i_3_0 ;
  wire \iv[2]_i_9_0 ;
  wire \iv[2]_i_9_1 ;
  wire \iv[2]_i_9_2 ;
  wire \iv[2]_i_9_n_0 ;
  wire \iv[3]_i_10_0 ;
  wire \iv[3]_i_10_1 ;
  wire \iv[3]_i_10_2 ;
  wire \iv[3]_i_15 ;
  wire \iv[3]_i_15_0 ;
  wire \iv[3]_i_19_n_0 ;
  wire \iv[3]_i_20 ;
  wire \iv[3]_i_21_n_0 ;
  wire \iv[3]_i_3 ;
  wire \iv[3]_i_3_0 ;
  wire \iv[3]_i_9_0 ;
  wire \iv[3]_i_9_1 ;
  wire \iv[3]_i_9_2 ;
  wire \iv[4]_i_10_0 ;
  wire \iv[4]_i_10_1 ;
  wire \iv[4]_i_10_2 ;
  wire \iv[4]_i_14 ;
  wire \iv[4]_i_14_0 ;
  wire \iv[4]_i_14_1 ;
  wire \iv[4]_i_17_0 ;
  wire \iv[4]_i_19_n_0 ;
  wire \iv[4]_i_21_n_0 ;
  wire \iv[4]_i_28_n_0 ;
  wire \iv[4]_i_29 ;
  wire \iv[4]_i_3 ;
  wire \iv[4]_i_9_0 ;
  wire \iv[4]_i_9_1 ;
  wire \iv[4]_i_9_2 ;
  wire \iv[5]_i_10_0 ;
  wire \iv[5]_i_10_1 ;
  wire \iv[5]_i_10_2 ;
  wire \iv[5]_i_14 ;
  wire \iv[5]_i_19_n_0 ;
  wire \iv[5]_i_21_n_0 ;
  wire \iv[5]_i_23 ;
  wire \iv[5]_i_28 ;
  wire \iv[5]_i_3 ;
  wire \iv[5]_i_3_0 ;
  wire \iv[5]_i_7 ;
  wire \iv[5]_i_9_0 ;
  wire \iv[5]_i_9_1 ;
  wire \iv[5]_i_9_2 ;
  wire \iv[6]_i_10 ;
  wire \iv[6]_i_10_0 ;
  wire \iv[6]_i_10_1 ;
  wire \iv[6]_i_15 ;
  wire \iv[6]_i_15_0 ;
  wire \iv[6]_i_9 ;
  wire \iv[6]_i_9_0 ;
  wire \iv[6]_i_9_1 ;
  wire \iv[6]_i_9_2 ;
  wire \iv[7]_i_16_n_0 ;
  wire \iv[7]_i_17 ;
  wire \iv[7]_i_17_0 ;
  wire \iv[7]_i_17_1 ;
  wire \iv[7]_i_18_n_0 ;
  wire \iv[7]_i_19_n_0 ;
  wire \iv[7]_i_20_n_0 ;
  wire \iv[7]_i_25 ;
  wire \iv[7]_i_3 ;
  wire \iv[7]_i_33 ;
  wire \iv[7]_i_3_0 ;
  wire \iv[7]_i_3_1 ;
  wire [1:0]\iv[7]_i_7 ;
  wire \iv[7]_i_7_0 ;
  wire \iv[7]_i_7_1 ;
  wire \iv[7]_i_7_2 ;
  wire \iv[7]_i_9_0 ;
  wire \iv[7]_i_9_1 ;
  wire \iv[7]_i_9_2 ;
  wire \iv[7]_i_9_3 ;
  wire \iv[7]_i_9_4 ;
  wire \iv[8]_i_10 ;
  wire \iv[8]_i_10_0 ;
  wire \iv[8]_i_12_n_0 ;
  wire \iv[8]_i_14_n_0 ;
  wire \iv[8]_i_16_n_0 ;
  wire \iv[8]_i_2 ;
  wire \iv[8]_i_2_0 ;
  wire \iv[8]_i_5_0 ;
  wire \iv[8]_i_5_1 ;
  wire \iv[8]_i_5_2 ;
  wire \iv[8]_i_5_3 ;
  wire \iv[8]_i_5_4 ;
  wire \iv[8]_i_5_5 ;
  wire \iv[8]_i_6_0 ;
  wire \iv[8]_i_6_1 ;
  wire \iv[8]_i_9 ;
  wire \iv[9]_i_10_n_0 ;
  wire \iv[9]_i_11 ;
  wire \iv[9]_i_11_0 ;
  wire \iv[9]_i_12_n_0 ;
  wire \iv[9]_i_14_n_0 ;
  wire \iv[9]_i_17_n_0 ;
  wire \iv[9]_i_2 ;
  wire \iv[9]_i_2_0 ;
  wire \iv[9]_i_2_1 ;
  wire \iv[9]_i_36 ;
  wire \iv[9]_i_44_n_0 ;
  wire \iv[9]_i_4_0 ;
  wire \iv[9]_i_4_1 ;
  wire \iv[9]_i_4_2 ;
  wire \iv[9]_i_4_3 ;
  wire \iv[9]_i_5_0 ;
  wire \iv[9]_i_5_1 ;
  wire \iv[9]_i_5_2 ;
  wire \iv[9]_i_5_3 ;
  wire \iv[9]_i_5_4 ;
  wire \niho_dsp_a[15]_INST_0_i_3 ;
  wire [1:0]\niho_dsp_a[32] ;
  wire \niho_dsp_a[32]_0 ;
  wire \niho_dsp_a[32]_1 ;
  wire \niho_dsp_a[32]_2 ;
  wire [0:0]p_0_in;
  wire [0:0]p_1_in;
  wire \sr[4]_i_114 ;
  wire \sr[4]_i_114_0 ;
  wire \sr[4]_i_135 ;
  wire \sr[4]_i_135_0 ;
  wire \sr[4]_i_135_1 ;
  wire \sr[4]_i_135_2 ;
  wire \sr[4]_i_146 ;
  wire \sr[4]_i_146_0 ;
  wire \sr[4]_i_146_1 ;
  wire \sr[4]_i_19 ;
  wire \sr[4]_i_21 ;
  wire \sr[4]_i_31 ;
  wire \sr[4]_i_31_0 ;
  wire \sr[4]_i_31_1 ;
  wire \sr[4]_i_33 ;
  wire \sr[4]_i_33_0 ;
  wire \sr[4]_i_33_1 ;
  wire \sr[4]_i_46 ;
  wire \sr[4]_i_46_0 ;
  wire \sr[4]_i_46_1 ;
  wire \sr[4]_i_47 ;
  wire \sr[4]_i_47_0 ;
  wire \sr[4]_i_82 ;
  wire \sr[4]_i_88 ;
  wire \sr[4]_i_88_0 ;
  wire \sr[7]_i_20 ;
  wire \sr_reg[6] ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[8] ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_9 ;
  wire \tr[17]_i_9 ;
  wire \tr[23]_i_10 ;
  wire \tr[25]_i_7 ;
  wire \tr[25]_i_7_0 ;
  wire \tr_reg[1] ;
  wire \tr_reg[1]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(\grn_reg[15]_1 [9]),
        .Q(Q[9]),
        .R(SR));
  LUT5 #(
    .INIT(32'h44777474)) 
    \iv[0]_i_12 
       (.I0(\sr[4]_i_146 ),
        .I1(\iv[0]_i_7 ),
        .I2(\iv[14]_i_19 ),
        .I3(\iv[0]_i_7_0 ),
        .I4(\iv[0]_i_7_1 ),
        .O(\niho_dsp_a[15]_INST_0_i_3 ));
  LUT4 #(
    .INIT(16'h1F11)) 
    \iv[10]_i_12 
       (.I0(\iv[10]_i_5_0 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\iv[10]_i_5_1 ),
        .I3(\sr_reg[8]_6 ),
        .O(\iv[10]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[10]_i_14 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[10]_i_5_2 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[10]_i_5_3 ),
        .I4(\iv[10]_i_5_4 ),
        .O(\iv[10]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[10]_i_16 
       (.I0(\sr_reg[8]_5 ),
        .I1(\iv[1]_i_15_0 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\iv[2]_i_10_0 ),
        .I4(\iv[10]_i_6 ),
        .O(\sr_reg[8]_26 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_32 
       (.I0(\sr_reg[8]_39 ),
        .I1(\iv[3]_i_20 ),
        .I2(\sr_reg[6] ),
        .O(\sr_reg[8]_36 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[10]_i_4 
       (.I0(\iv[9]_i_2_0 ),
        .I1(\iv[10]_i_2_1 ),
        .I2(\iv[10]_i_2_2 ),
        .O(\iv[10]_i_10 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_46 
       (.I0(\sr[4]_i_114 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\sr[4]_i_114_0 ),
        .O(\sr_reg[8]_39 ));
  LUT5 #(
    .INIT(32'h2AFF2A00)) 
    \iv[10]_i_47 
       (.I0(\sr[4]_i_135 ),
        .I1(\niho_dsp_a[32] [0]),
        .I2(\sr[4]_i_146 ),
        .I3(\iv[12]_i_21_0 ),
        .I4(\sr[4]_i_135_0 ),
        .O(\sr_reg[6] ));
  LUT6 #(
    .INIT(64'hCF00CF00DDDDDD00)) 
    \iv[10]_i_5 
       (.I0(\iv[10]_i_2 ),
        .I1(\iv[10]_i_12_n_0 ),
        .I2(\iv[10]_i_2_0 ),
        .I3(\iv[10]_i_14_n_0 ),
        .I4(\niho_dsp_a[32] [1]),
        .I5(\iv[5]_i_7 ),
        .O(\sr_reg[8]_11 ));
  LUT6 #(
    .INIT(64'h0001F00100F1F0F1)) 
    \iv[11]_i_12 
       (.I0(\sr_reg[8]_1 ),
        .I1(\iv[5]_i_7 ),
        .I2(\sr[4]_i_82 ),
        .I3(\iv[8]_i_5_0 ),
        .I4(\iv[11]_i_5_0 ),
        .I5(\iv[11]_i_5_1 ),
        .O(\iv[11]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[11]_i_14 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[11]_i_5_2 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[11]_i_5_3 ),
        .I4(\iv[11]_i_5_4 ),
        .O(\iv[11]_i_14_n_0 ));
  LUT4 #(
    .INIT(16'hBBB8)) 
    \iv[11]_i_15 
       (.I0(\iv[11]_i_6_0 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\iv[3]_i_20 ),
        .I3(\sr_reg[8]_45 ),
        .O(\sr_reg[8]_1 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[11]_i_16 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[11]_i_6_0 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\sr_reg[8]_45 ),
        .I4(\sr_reg[6]_3 ),
        .O(\iv[11]_i_16_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_34 
       (.I0(\tr[17]_i_9 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\sr[4]_i_146_0 ),
        .O(\sr_reg[8]_45 ));
  LUT5 #(
    .INIT(32'hF044F077)) 
    \iv[11]_i_35 
       (.I0(DI[1]),
        .I1(\sr[4]_i_146 ),
        .I2(\sr[4]_i_146_1 ),
        .I3(\iv[12]_i_21_0 ),
        .I4(\niho_dsp_a[32] [0]),
        .O(\sr_reg[6]_3 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_36 
       (.I0(\iv[1]_i_23_1 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\iv[11]_i_18 ),
        .O(\sr_reg[8]_44 ));
  LUT5 #(
    .INIT(32'hF011F0DD)) 
    \iv[11]_i_37 
       (.I0(DI[1]),
        .I1(\sr[4]_i_146 ),
        .I2(\iv[11]_i_18_0 ),
        .I3(\iv[12]_i_21_0 ),
        .I4(\niho_dsp_a[32] [0]),
        .O(\sr_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[11]_i_5 
       (.I0(\iv[11]_i_12_n_0 ),
        .I1(\iv[11]_i_2 ),
        .I2(\iv[11]_i_14_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8]_0 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[11]_i_6 
       (.I0(\iv[11]_i_2 ),
        .I1(bbus_0[0]),
        .I2(\sr_reg[8]_1 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[9]_i_4_1 ),
        .I5(\iv[11]_i_16_n_0 ),
        .O(\sr_reg[8]_31 ));
  LUT4 #(
    .INIT(16'h444F)) 
    \iv[12]_i_11 
       (.I0(\iv[12]_i_5_0 ),
        .I1(\sr_reg[8]_6 ),
        .I2(\iv[12]_i_5_1 ),
        .I3(\sr_reg[8]_5 ),
        .O(\iv[12]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[12]_i_14 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[12]_i_5_2 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[12]_i_5_3 ),
        .I4(\iv[12]_i_5_4 ),
        .O(\iv[12]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[12]_i_16 
       (.I0(\sr_reg[8]_5 ),
        .I1(\iv[3]_i_15 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\iv[4]_i_10_0 ),
        .I4(\iv[12]_i_6 ),
        .O(\sr_reg[8]_25 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[12]_i_32 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[12]_i_15_0 ),
        .I2(\iv[12]_i_15 ),
        .O(\sr_reg[8]_35 ));
  LUT6 #(
    .INIT(64'hAF00AF00BBBBBB00)) 
    \iv[12]_i_5 
       (.I0(\iv[12]_i_11_n_0 ),
        .I1(\iv[12]_i_2 ),
        .I2(\iv[12]_i_2_0 ),
        .I3(\iv[12]_i_14_n_0 ),
        .I4(\niho_dsp_a[32] [1]),
        .I5(\iv[5]_i_7 ),
        .O(\sr_reg[8]_10 ));
  LUT4 #(
    .INIT(16'h1F11)) 
    \iv[13]_i_11 
       (.I0(\iv[13]_i_5_0 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\iv[13]_i_5_1 ),
        .I3(\sr_reg[8]_6 ),
        .O(\iv[13]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[13]_i_14 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[13]_i_5_2 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[13]_i_5_3 ),
        .I4(\iv[13]_i_5_4 ),
        .O(\iv[13]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'h0000ABFB)) 
    \iv[13]_i_16 
       (.I0(\sr_reg[8]_5 ),
        .I1(\iv[4]_i_14 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\iv[5]_i_10_0 ),
        .I4(\iv[13]_i_6 ),
        .O(\sr_reg[8]_24 ));
  LUT4 #(
    .INIT(16'h60CC)) 
    \iv[13]_i_21 
       (.I0(\iv[5]_i_7 ),
        .I1(bbus_0[0]),
        .I2(\niho_dsp_a[32] [1]),
        .I3(\iv[12]_i_9 ),
        .O(\sr_reg[8]_37 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[13]_i_27 
       (.I0(\iv[8]_i_5_0 ),
        .I1(\sr[4]_i_82 ),
        .O(\sr_reg[8]_6 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[13]_i_34 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[13]_i_15_0 ),
        .I2(\iv[13]_i_15 ),
        .O(\sr_reg[8]_49 ));
  LUT6 #(
    .INIT(64'hAF00AF00BBBBBB00)) 
    \iv[13]_i_5 
       (.I0(\iv[13]_i_11_n_0 ),
        .I1(\iv[13]_i_2 ),
        .I2(\iv[13]_i_2_0 ),
        .I3(\iv[13]_i_14_n_0 ),
        .I4(\niho_dsp_a[32] [1]),
        .I5(\iv[5]_i_7 ),
        .O(\sr_reg[8]_9 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[14]_i_10 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[14]_i_6 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\sr_reg[8]_41 ),
        .I4(\sr_reg[8]_40 ),
        .O(\sr_reg[8]_16 ));
  LUT6 #(
    .INIT(64'h350035003500350F)) 
    \iv[14]_i_12 
       (.I0(\iv[14]_i_5_0 ),
        .I1(\iv[14]_i_5_1 ),
        .I2(\iv[8]_i_5_0 ),
        .I3(\sr[4]_i_82 ),
        .I4(\sr_reg[8]_16 ),
        .I5(\iv[5]_i_7 ),
        .O(\iv[14]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[14]_i_14 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[14]_i_5_2 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[14]_i_5_3 ),
        .I4(\iv[14]_i_5_4 ),
        .O(\iv[14]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_25 
       (.I0(\sr[4]_i_135_1 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\sr[4]_i_135_2 ),
        .O(\sr_reg[8]_41 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_26 
       (.I0(\sr[4]_i_135 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\sr[4]_i_135_0 ),
        .O(\sr_reg[8]_40 ));
  LUT5 #(
    .INIT(32'h47FF4700)) 
    \iv[14]_i_36 
       (.I0(\iv[14]_i_19 ),
        .I1(\sr[4]_i_146 ),
        .I2(\niho_dsp_a[32] [0]),
        .I3(\iv[12]_i_21_0 ),
        .I4(\iv[12]_i_21 ),
        .O(\sr_reg[6]_2 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[14]_i_5 
       (.I0(\iv[14]_i_12_n_0 ),
        .I1(\iv[14]_i_2 ),
        .I2(\iv[14]_i_14_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8]_15 ));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[1]_i_10 
       (.I0(\iv[1]_i_20_n_0 ),
        .I1(\iv[1]_i_3_0 ),
        .I2(\iv[1]_i_21_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(bbus_0[0]),
        .O(\iv[1]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'hF444F4F4F4444444)) 
    \iv[1]_i_14 
       (.I0(\sr_reg[8]_18 ),
        .I1(\iv[9]_i_4_3 ),
        .I2(\iv[9]_i_4_2 ),
        .I3(\iv[9]_i_4_0 ),
        .I4(\iv[9]_i_4_1 ),
        .I5(\sr_reg[8]_19 ),
        .O(\iv[1]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[1]_i_16 
       (.I0(\iv[9]_i_4_1 ),
        .I1(\sr[4]_i_82 ),
        .I2(\sr_reg[8]_18 ),
        .O(\sr_reg[8]_3 ));
  LUT4 #(
    .INIT(16'h444F)) 
    \iv[1]_i_17 
       (.I0(\iv[1]_i_9_0 ),
        .I1(\sr_reg[8]_6 ),
        .I2(\iv[1]_i_9_1 ),
        .I3(\sr_reg[8]_5 ),
        .O(\iv[1]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[1]_i_19 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[1]_i_9_2 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[1]_i_9_3 ),
        .I4(\iv[1]_i_9_4 ),
        .O(\iv[1]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[1]_i_20 
       (.I0(\iv[1]_i_31_n_0 ),
        .I1(\iv[4]_i_10_1 ),
        .I2(\iv[1]_i_10_3 ),
        .I3(\sr[4]_i_82 ),
        .I4(\sr_reg[8]_3 ),
        .I5(bbus_0[0]),
        .O(\iv[1]_i_20_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \iv[1]_i_21 
       (.I0(\sr_reg[8]_5 ),
        .I1(\iv[1]_i_10_0 ),
        .I2(\iv[1]_i_10_1 ),
        .I3(\iv[8]_i_5_0 ),
        .I4(\iv[1]_i_10_2 ),
        .I5(\niho_dsp_a[32] [1]),
        .O(\iv[1]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'hFEFF)) 
    \iv[1]_i_22 
       (.I0(\iv[12]_i_21_0 ),
        .I1(\tr[17]_i_9 ),
        .I2(\iv[3]_i_20 ),
        .I3(\iv[4]_i_14_0 ),
        .O(\sr_reg[8]_18 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[1]_i_23 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[1]_i_15_0 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\sr_reg[8]_43 ),
        .I4(\iv[9]_i_44_n_0 ),
        .O(\sr_reg[8]_19 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[1]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\iv[1]_i_15 ),
        .I2(\iv[1]_i_9_n_0 ),
        .I3(\iv[1]_i_10_n_0 ),
        .I4(\tr_reg[1]_0 ),
        .O(\sr_reg[8]_2 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[1]_i_31 
       (.I0(\iv[1]_i_20_0 ),
        .I1(\iv[3]_i_20 ),
        .I2(\iv[13]_i_15 ),
        .O(\iv[1]_i_31_n_0 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[1]_i_8 
       (.I0(\iv[9]_i_2_0 ),
        .I1(\iv[1]_i_14_n_0 ),
        .I2(\sr[4]_i_19 ),
        .O(\iv[1]_i_15 ));
  LUT6 #(
    .INIT(64'hCF00CF00DDDDDD00)) 
    \iv[1]_i_9 
       (.I0(\sr_reg[8]_3 ),
        .I1(\iv[1]_i_17_n_0 ),
        .I2(\iv[1]_i_3_0 ),
        .I3(\iv[1]_i_19_n_0 ),
        .I4(\niho_dsp_a[32] [1]),
        .I5(\iv[5]_i_7 ),
        .O(\iv[1]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[2]_i_10 
       (.I0(\bdatw[12]_INST_0_i_1 ),
        .I1(\iv[2]_i_3_0 ),
        .I2(\iv[2]_i_20_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(bbus_0[0]),
        .O(\iv[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[2]_i_14 
       (.I0(\iv[9]_i_4_2 ),
        .I1(\iv[9]_i_4_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\sr_reg[8]_20 ),
        .I4(\sr_reg[8]_21 ),
        .I5(\iv[9]_i_4_3 ),
        .O(\iv[2]_i_14_n_0 ));
  LUT6 #(
    .INIT(64'h111F111FFFFF111F)) 
    \iv[2]_i_16 
       (.I0(\sr[4]_i_47 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\iv[5]_i_7 ),
        .I3(\iv[2]_i_25_n_0 ),
        .I4(\sr_reg[8]_6 ),
        .I5(\sr[4]_i_47_0 ),
        .O(\iv[2]_i_26 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[2]_i_18 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[2]_i_9_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[2]_i_9_1 ),
        .I4(\iv[2]_i_9_2 ),
        .O(\iv[2]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[2]_i_19 
       (.I0(\sr_reg[8]_36 ),
        .I1(\iv[4]_i_10_1 ),
        .I2(\iv[11]_i_6_0 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[2]_i_25_n_0 ),
        .I5(bbus_0[0]),
        .O(\bdatw[12]_INST_0_i_1 ));
  LUT5 #(
    .INIT(32'h0000F2F7)) 
    \iv[2]_i_20 
       (.I0(\iv[4]_i_10_1 ),
        .I1(\iv[2]_i_15_0 ),
        .I2(\sr_reg[8]_5 ),
        .I3(\iv[2]_i_10_0 ),
        .I4(\iv[2]_i_10_1 ),
        .O(\iv[2]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[2]_i_21 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[2]_i_15_0 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\iv[2]_i_15_1 ),
        .I4(\iv[2]_i_15_2 ),
        .O(\sr_reg[8]_20 ));
  LUT5 #(
    .INIT(32'hFFB8FFFF)) 
    \iv[2]_i_22 
       (.I0(\sr[4]_i_135 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\sr[4]_i_135_0 ),
        .I3(\iv[3]_i_20 ),
        .I4(\iv[4]_i_14_0 ),
        .O(\sr_reg[8]_21 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[2]_i_25 
       (.I0(\iv[9]_i_4_1 ),
        .I1(\sr[4]_i_82 ),
        .I2(\sr_reg[8]_21 ),
        .O(\iv[2]_i_25_n_0 ));
  LUT5 #(
    .INIT(32'hA8AA8888)) 
    \iv[2]_i_3 
       (.I0(\tr_reg[1] ),
        .I1(\iv[2]_i_15 ),
        .I2(\iv[2]_i_9_n_0 ),
        .I3(\iv[2]_i_10_n_0 ),
        .I4(\tr_reg[1]_0 ),
        .O(\sr_reg[8]_4 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[2]_i_8 
       (.I0(\iv[9]_i_2_0 ),
        .I1(\iv[2]_i_14_n_0 ),
        .I2(\sr[4]_i_21 ),
        .O(\iv[2]_i_15 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[2]_i_9 
       (.I0(\iv[2]_i_26 ),
        .I1(\iv[2]_i_3_0 ),
        .I2(\iv[2]_i_18_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\iv[2]_i_9_n_0 ));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[3]_i_10 
       (.I0(\iv[3]_i_3_0 ),
        .I1(\iv[3]_i_3 ),
        .I2(\iv[3]_i_21_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(bbus_0[0]),
        .O(\sr_reg[8]_23 ));
  LUT6 #(
    .INIT(64'h550000035500FF03)) 
    \iv[3]_i_17 
       (.I0(\sr[4]_i_46 ),
        .I1(\iv[5]_i_7 ),
        .I2(\sr[4]_i_46_0 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[9]_i_4_1 ),
        .I5(\sr[4]_i_46_1 ),
        .O(\sr_reg[8]_8 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[3]_i_19 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[3]_i_9_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[3]_i_9_1 ),
        .I4(\iv[3]_i_9_2 ),
        .O(\iv[3]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \iv[3]_i_21 
       (.I0(\sr_reg[8]_5 ),
        .I1(\iv[3]_i_10_0 ),
        .I2(\iv[3]_i_10_1 ),
        .I3(\iv[8]_i_5_0 ),
        .I4(\iv[3]_i_10_2 ),
        .I5(\niho_dsp_a[32] [1]),
        .O(\iv[3]_i_21_n_0 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[3]_i_28 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[3]_i_15 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\sr_reg[8]_44 ),
        .I4(\iv[3]_i_15_0 ),
        .O(\sr_reg[8]_48 ));
  LUT3 #(
    .INIT(8'hE4)) 
    \iv[3]_i_36 
       (.I0(\iv[3]_i_20 ),
        .I1(\sr_reg[8]_45 ),
        .I2(\sr_reg[6]_3 ),
        .O(\sr_reg[8]_47 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[3]_i_9 
       (.I0(\sr_reg[8]_8 ),
        .I1(\iv[3]_i_3 ),
        .I2(\iv[3]_i_19_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8]_7 ));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[4]_i_10 
       (.I0(\bdatw[12]_INST_0_i_1_0 ),
        .I1(\iv[4]_i_3 ),
        .I2(\iv[4]_i_21_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(bbus_0[0]),
        .O(\sr_reg[8]_28 ));
  LUT5 #(
    .INIT(32'h3A3F3035)) 
    \iv[4]_i_16 
       (.I0(\iv[3]_i_20 ),
        .I1(\iv[4]_i_14 ),
        .I2(\iv[4]_i_14_0 ),
        .I3(\sr_reg[8]_38 ),
        .I4(\iv[4]_i_14_1 ),
        .O(\sr_reg[8]_50 ));
  LUT6 #(
    .INIT(64'h444F444F444FFFFF)) 
    \iv[4]_i_17 
       (.I0(\sr[4]_i_31 ),
        .I1(\sr_reg[8]_6 ),
        .I2(\iv[5]_i_7 ),
        .I3(\iv[4]_i_28_n_0 ),
        .I4(\sr_reg[8]_5 ),
        .I5(\sr[4]_i_31_0 ),
        .O(\iv[4]_i_29 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[4]_i_19 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[4]_i_9_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[4]_i_9_1 ),
        .I4(\iv[4]_i_9_2 ),
        .O(\iv[4]_i_19_n_0 ));
  LUT6 #(
    .INIT(64'h470047004700FFFF)) 
    \iv[4]_i_20 
       (.I0(\sr_reg[8]_35 ),
        .I1(\iv[4]_i_10_1 ),
        .I2(\sr[4]_i_31_1 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[4]_i_28_n_0 ),
        .I5(bbus_0[0]),
        .O(\bdatw[12]_INST_0_i_1_0 ));
  LUT5 #(
    .INIT(32'h0000F2F7)) 
    \iv[4]_i_21 
       (.I0(\iv[4]_i_10_1 ),
        .I1(\iv[4]_i_14 ),
        .I2(\sr_reg[8]_5 ),
        .I3(\iv[4]_i_10_0 ),
        .I4(\iv[4]_i_10_2 ),
        .O(\iv[4]_i_21_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_25 
       (.I0(\iv[12]_i_21 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\iv[12]_i_21_1 ),
        .O(\sr_reg[8]_38 ));
  LUT3 #(
    .INIT(8'hFE)) 
    \iv[4]_i_28 
       (.I0(\iv[9]_i_4_1 ),
        .I1(\sr[4]_i_82 ),
        .I2(\iv[4]_i_17_0 ),
        .O(\iv[4]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[4]_i_9 
       (.I0(\iv[4]_i_29 ),
        .I1(\iv[4]_i_3 ),
        .I2(\iv[4]_i_19_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8]_13 ));
  LUT5 #(
    .INIT(32'h4F4F5F55)) 
    \iv[5]_i_10 
       (.I0(\iv[5]_i_3_0 ),
        .I1(\iv[5]_i_3 ),
        .I2(\iv[5]_i_21_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(bbus_0[0]),
        .O(\sr_reg[8]_27 ));
  LUT5 #(
    .INIT(32'h47774744)) 
    \iv[5]_i_12 
       (.I0(\iv[5]_i_7 ),
        .I1(\iv[0]_i_7 ),
        .I2(DI[0]),
        .I3(\iv[0]_i_7_1 ),
        .I4(\iv[7]_i_7 [0]),
        .O(\badr[5]_INST_0_i_1 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[5]_i_15 
       (.I0(\iv[5]_i_10_1 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\iv[5]_i_14 ),
        .O(\iv[5]_i_23 ));
  LUT6 #(
    .INIT(64'h111F111FFFFF111F)) 
    \iv[5]_i_17 
       (.I0(\sr[4]_i_33 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\iv[5]_i_7 ),
        .I3(\sr[4]_i_33_0 ),
        .I4(\sr_reg[8]_6 ),
        .I5(\sr[4]_i_33_1 ),
        .O(\iv[5]_i_28 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[5]_i_19 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[5]_i_9_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[5]_i_9_1 ),
        .I4(\iv[5]_i_9_2 ),
        .O(\iv[5]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h0000F2F7)) 
    \iv[5]_i_21 
       (.I0(\iv[4]_i_10_1 ),
        .I1(\iv[5]_i_10_1 ),
        .I2(\sr_reg[8]_5 ),
        .I3(\iv[5]_i_10_0 ),
        .I4(\iv[5]_i_10_2 ),
        .O(\iv[5]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \iv[5]_i_25 
       (.I0(\iv[12]_i_21_0 ),
        .I1(\tr[17]_i_9 ),
        .O(\sr_reg[8]_42 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[5]_i_9 
       (.I0(\iv[5]_i_28 ),
        .I1(\iv[5]_i_3 ),
        .I2(\iv[5]_i_19_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8]_12 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[6]_i_19 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[6]_i_9_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[6]_i_9_1 ),
        .I4(\iv[6]_i_9_2 ),
        .O(\sr_reg[8]_34 ));
  LUT6 #(
    .INIT(64'h00000000FEFE00FE)) 
    \iv[6]_i_22 
       (.I0(\sr_reg[8]_5 ),
        .I1(\iv[6]_i_10 ),
        .I2(\iv[6]_i_10_0 ),
        .I3(\iv[8]_i_5_0 ),
        .I4(\iv[6]_i_10_1 ),
        .I5(\niho_dsp_a[32] [1]),
        .O(\sr_reg[8]_29 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[6]_i_23 
       (.I0(\iv[6]_i_15 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\iv[6]_i_15_0 ),
        .O(\iv[14]_i_49 ));
  LUT6 #(
    .INIT(64'h00000000AFAFEFE0)) 
    \iv[7]_i_10 
       (.I0(\iv[7]_i_3_0 ),
        .I1(\sr_reg[8]_30 ),
        .I2(bbus_0[0]),
        .I3(\sr[7]_i_20 ),
        .I4(\iv[7]_i_9_4 ),
        .I5(\iv[7]_i_3_1 ),
        .O(\iv[7]_i_25 ));
  LUT6 #(
    .INIT(64'h505F30305F5F3F3F)) 
    \iv[7]_i_13 
       (.I0(\iv[9]_i_4_0 ),
        .I1(\iv[7]_i_7 [1]),
        .I2(\iv[7]_i_7_0 ),
        .I3(DI[1]),
        .I4(\iv[7]_i_7_1 ),
        .I5(\iv[7]_i_7_2 ),
        .O(\iv[7]_i_33 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[7]_i_16 
       (.I0(\iv[9]_i_4_2 ),
        .I1(\iv[9]_i_4_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\iv[15]_i_94 ),
        .I4(\sr[7]_i_20 ),
        .I5(\iv[9]_i_4_3 ),
        .O(\iv[7]_i_16_n_0 ));
  LUT6 #(
    .INIT(64'h550000035500FF03)) 
    \iv[7]_i_18 
       (.I0(\iv[7]_i_9_0 ),
        .I1(\iv[5]_i_7 ),
        .I2(\sr[7]_i_20 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[9]_i_4_1 ),
        .I5(\iv[7]_i_9_1 ),
        .O(\iv[7]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h00A2)) 
    \iv[7]_i_19 
       (.I0(\iv[5]_i_7 ),
        .I1(\sr_reg[8]_30 ),
        .I2(\iv[7]_i_9_4 ),
        .I3(\iv[7]_i_3_0 ),
        .O(\iv[7]_i_19_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[7]_i_20 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[7]_i_9_2 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\sr_reg[8]_30 ),
        .I4(\iv[7]_i_9_3 ),
        .O(\iv[7]_i_20_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[7]_i_22 
       (.I0(\iv[7]_i_17_0 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\sr[4]_i_88 ),
        .I3(\iv[3]_i_20 ),
        .I4(\sr[4]_i_88_0 ),
        .O(\sr_reg[8]_30 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[7]_i_23 
       (.I0(\tr[23]_i_10 ),
        .I1(\iv[4]_i_14_0 ),
        .O(\sr[7]_i_20 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[7]_i_35 
       (.I0(\iv[7]_i_17_0 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\iv[7]_i_17_1 ),
        .O(\iv[15]_i_94 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[7]_i_8 
       (.I0(\iv[9]_i_2_0 ),
        .I1(\iv[7]_i_16_n_0 ),
        .I2(\iv[7]_i_3 ),
        .O(\iv[7]_i_17 ));
  LUT5 #(
    .INIT(32'hE0E0EEE0)) 
    \iv[7]_i_9 
       (.I0(\iv[7]_i_18_n_0 ),
        .I1(\iv[7]_i_19_n_0 ),
        .I2(\iv[7]_i_20_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8] ));
  LUT6 #(
    .INIT(64'hA300A300A300A30F)) 
    \iv[8]_i_12 
       (.I0(\iv[8]_i_5_1 ),
        .I1(\iv[8]_i_5_2 ),
        .I2(\iv[8]_i_5_0 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[8]_i_2_0 ),
        .I5(\iv[5]_i_7 ),
        .O(\iv[8]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[8]_i_14 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[8]_i_5_3 ),
        .I2(\iv[8]_i_5_0 ),
        .I3(\iv[8]_i_5_4 ),
        .I4(\iv[8]_i_5_5 ),
        .O(\iv[8]_i_14_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[8]_i_16 
       (.I0(\iv[8]_i_6_0 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\iv[8]_i_6_1 ),
        .I3(\iv[3]_i_20 ),
        .I4(\iv[12]_i_15 ),
        .O(\iv[8]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'hB)) 
    \iv[8]_i_20 
       (.I0(\iv[8]_i_5_0 ),
        .I1(\sr[4]_i_82 ),
        .O(\sr_reg[8]_5 ));
  LUT6 #(
    .INIT(64'h1DFF1D331D331DFF)) 
    \iv[8]_i_21 
       (.I0(\iv[8]_i_9 ),
        .I1(\iv[0]_i_7 ),
        .I2(\sr[4]_i_146 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[0]_i_7_0 ),
        .I5(bbus_0[1]),
        .O(\bdatw[8]_INST_0_i_2 ));
  LUT3 #(
    .INIT(8'h74)) 
    \iv[8]_i_24 
       (.I0(\iv[8]_i_10 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\iv[8]_i_10_0 ),
        .O(\iv[0]_i_25 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[8]_i_5 
       (.I0(\iv[8]_i_12_n_0 ),
        .I1(\iv[8]_i_2 ),
        .I2(\iv[8]_i_14_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8]_14 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[8]_i_6 
       (.I0(\iv[8]_i_2 ),
        .I1(bbus_0[0]),
        .I2(\iv[8]_i_2_0 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[9]_i_4_1 ),
        .I5(\iv[8]_i_16_n_0 ),
        .O(\sr_reg[8]_32 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[9]_i_10 
       (.I0(\iv[9]_i_4_2 ),
        .I1(\iv[9]_i_4_0 ),
        .I2(\iv[9]_i_4_1 ),
        .I3(\sr_reg[8]_22 ),
        .I4(\iv[9]_i_36 ),
        .I5(\iv[9]_i_4_3 ),
        .O(\iv[9]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h0001F00100F1F0F1)) 
    \iv[9]_i_12 
       (.I0(\iv[9]_i_36 ),
        .I1(\iv[5]_i_7 ),
        .I2(\sr[4]_i_82 ),
        .I3(\iv[8]_i_5_0 ),
        .I4(\iv[9]_i_5_0 ),
        .I5(\iv[9]_i_5_1 ),
        .O(\iv[9]_i_12_n_0 ));
  LUT5 #(
    .INIT(32'h0000BABF)) 
    \iv[9]_i_14 
       (.I0(\iv[6]_i_9 ),
        .I1(\iv[9]_i_5_2 ),
        .I2(\iv[8]_i_5_0 ),
        .I3(\iv[9]_i_5_3 ),
        .I4(\iv[9]_i_5_4 ),
        .O(\iv[9]_i_14_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_15 
       (.I0(\tr[25]_i_7 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\tr[25]_i_7_0 ),
        .O(\iv[9]_i_36 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_17 
       (.I0(\tr[25]_i_7 ),
        .I1(\iv[4]_i_14_0 ),
        .I2(\iv[1]_i_20_0 ),
        .I3(\iv[3]_i_20 ),
        .I4(\iv[13]_i_15 ),
        .O(\iv[9]_i_17_n_0 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[9]_i_25 
       (.I0(\iv[3]_i_20 ),
        .I1(\sr_reg[8]_43 ),
        .I2(\iv[9]_i_44_n_0 ),
        .I3(\iv[4]_i_14_0 ),
        .I4(\iv[9]_i_11_0 ),
        .O(\sr_reg[8]_22 ));
  LUT5 #(
    .INIT(32'h1DFF1D00)) 
    \iv[9]_i_39 
       (.I0(DI[1]),
        .I1(\sr[4]_i_146 ),
        .I2(\niho_dsp_a[32] [0]),
        .I3(\iv[12]_i_21_0 ),
        .I4(\iv[1]_i_23_1 ),
        .O(\sr_reg[6]_1 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[9]_i_4 
       (.I0(\iv[9]_i_2_0 ),
        .I1(\iv[9]_i_10_n_0 ),
        .I2(\iv[9]_i_2_1 ),
        .O(\iv[9]_i_11 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_40 
       (.I0(\iv[11]_i_18 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\iv[1]_i_32 ),
        .O(\sr_reg[8]_43 ));
  LUT3 #(
    .INIT(8'h8B)) 
    \iv[9]_i_44 
       (.I0(\iv[1]_i_23_0 ),
        .I1(\iv[12]_i_21_0 ),
        .I2(\iv[1]_i_23_1 ),
        .O(\iv[9]_i_44_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[9]_i_5 
       (.I0(\iv[9]_i_12_n_0 ),
        .I1(\iv[9]_i_2 ),
        .I2(\iv[9]_i_14_n_0 ),
        .I3(\niho_dsp_a[32] [1]),
        .I4(\iv[5]_i_7 ),
        .O(\sr_reg[8]_17 ));
  LUT6 #(
    .INIT(64'hBBBBBBB800BB00B8)) 
    \iv[9]_i_6 
       (.I0(\iv[9]_i_2 ),
        .I1(bbus_0[0]),
        .I2(\iv[9]_i_36 ),
        .I3(\sr[4]_i_82 ),
        .I4(\iv[8]_i_5_0 ),
        .I5(\iv[9]_i_17_n_0 ),
        .O(\sr_reg[8]_33 ));
  LUT6 #(
    .INIT(64'h00000000FFFFFFFE)) 
    \niho_dsp_a[32]_INST_0_i_2 
       (.I0(\niho_dsp_a[32]_0 ),
        .I1(\niho_dsp_a[32]_1 ),
        .I2(p_0_in),
        .I3(p_1_in),
        .I4(\niho_dsp_a[32]_2 ),
        .I5(\niho_dsp_a[32] [1]),
        .O(\sr_reg[8]_46 ));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_7
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_8
   (Q,
    SR,
    \grn_reg[15]_0 ,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]\grn_reg[15]_0 ;
  input [15:0]cbus;
  input clk;

  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  wire [0:0]\grn_reg[15]_0 ;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(\grn_reg[15]_0 ),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

(* ORIG_REF_NAME = "niho_rgf_grn" *) 
module niho_rgf_grn_9
   (Q,
    SR,
    E,
    cbus,
    clk);
  output [15:0]Q;
  input [0:0]SR;
  input [0:0]E;
  input [15:0]cbus;
  input clk;

  wire [0:0]E;
  wire [15:0]Q;
  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;

  FDRE \grn_reg[0] 
       (.C(clk),
        .CE(E),
        .D(cbus[0]),
        .Q(Q[0]),
        .R(SR));
  FDRE \grn_reg[10] 
       (.C(clk),
        .CE(E),
        .D(cbus[10]),
        .Q(Q[10]),
        .R(SR));
  FDRE \grn_reg[11] 
       (.C(clk),
        .CE(E),
        .D(cbus[11]),
        .Q(Q[11]),
        .R(SR));
  FDRE \grn_reg[12] 
       (.C(clk),
        .CE(E),
        .D(cbus[12]),
        .Q(Q[12]),
        .R(SR));
  FDRE \grn_reg[13] 
       (.C(clk),
        .CE(E),
        .D(cbus[13]),
        .Q(Q[13]),
        .R(SR));
  FDRE \grn_reg[14] 
       (.C(clk),
        .CE(E),
        .D(cbus[14]),
        .Q(Q[14]),
        .R(SR));
  FDRE \grn_reg[15] 
       (.C(clk),
        .CE(E),
        .D(cbus[15]),
        .Q(Q[15]),
        .R(SR));
  FDRE \grn_reg[1] 
       (.C(clk),
        .CE(E),
        .D(cbus[1]),
        .Q(Q[1]),
        .R(SR));
  FDRE \grn_reg[2] 
       (.C(clk),
        .CE(E),
        .D(cbus[2]),
        .Q(Q[2]),
        .R(SR));
  FDRE \grn_reg[3] 
       (.C(clk),
        .CE(E),
        .D(cbus[3]),
        .Q(Q[3]),
        .R(SR));
  FDRE \grn_reg[4] 
       (.C(clk),
        .CE(E),
        .D(cbus[4]),
        .Q(Q[4]),
        .R(SR));
  FDRE \grn_reg[5] 
       (.C(clk),
        .CE(E),
        .D(cbus[5]),
        .Q(Q[5]),
        .R(SR));
  FDRE \grn_reg[6] 
       (.C(clk),
        .CE(E),
        .D(cbus[6]),
        .Q(Q[6]),
        .R(SR));
  FDRE \grn_reg[7] 
       (.C(clk),
        .CE(E),
        .D(cbus[7]),
        .Q(Q[7]),
        .R(SR));
  FDRE \grn_reg[8] 
       (.C(clk),
        .CE(E),
        .D(cbus[8]),
        .Q(Q[8]),
        .R(SR));
  FDRE \grn_reg[9] 
       (.C(clk),
        .CE(E),
        .D(cbus[9]),
        .Q(Q[9]),
        .R(SR));
endmodule

module niho_rgf_ivec
   (.\iv_reg[15]_0 ({iv[15],iv[14],iv[13],iv[12],iv[11],iv[10],iv[9],iv[8],iv[7],iv[6],iv[5],iv[4],iv[3],iv[2],iv[1],iv[0]}),
    SR,
    \iv_reg[0]_0 ,
    cbus,
    clk);
  input [0:0]SR;
  input [0:0]\iv_reg[0]_0 ;
  input [15:0]cbus;
  input clk;
     output [15:0]iv;

  wire [0:0]SR;
  wire [15:0]cbus;
  wire clk;
  (* DONT_TOUCH *) wire [15:0]iv;
  wire [0:0]\iv_reg[0]_0 ;

  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[0] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[0]),
        .Q(iv[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[10] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[10]),
        .Q(iv[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[11] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[11]),
        .Q(iv[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[12] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[12]),
        .Q(iv[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[13] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[13]),
        .Q(iv[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[14] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[14]),
        .Q(iv[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[15] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[15]),
        .Q(iv[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[1] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[1]),
        .Q(iv[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[2] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[2]),
        .Q(iv[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[3] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[3]),
        .Q(iv[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[4] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[4]),
        .Q(iv[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[5] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[5]),
        .Q(iv[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[6] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[6]),
        .Q(iv[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[7] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[7]),
        .Q(iv[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[8] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[8]),
        .Q(iv[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \iv_reg[9] 
       (.C(clk),
        .CE(\iv_reg[0]_0 ),
        .D(cbus[9]),
        .Q(iv[9]),
        .R(SR));
endmodule

module niho_rgf_pcnt
   (.out({pc[15],pc[14],pc[13],pc[12],pc[11],pc[10],pc[9],pc[8],pc[7],pc[6],pc[5],pc[4],pc[3],pc[2],pc[1],pc[0]}),
    fch_pc,
    S,
    SR,
    \pc_reg[15]_0 ,
    clk);
  output [15:0]fch_pc;
  input [0:0]S;
  input [0:0]SR;
  input [15:0]\pc_reg[15]_0 ;
  input clk;
     output [15:0]pc;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]S;
  wire [0:0]SR;
  wire clk;
  wire [15:0]fch_pc;
  (* DONT_TOUCH *) wire [15:0]pc;
  wire \pc_reg[11]_i_2_n_0 ;
  wire \pc_reg[11]_i_2_n_1 ;
  wire \pc_reg[11]_i_2_n_2 ;
  wire \pc_reg[11]_i_2_n_3 ;
  wire [15:0]\pc_reg[15]_0 ;
  wire \pc_reg[15]_i_3_n_1 ;
  wire \pc_reg[15]_i_3_n_2 ;
  wire \pc_reg[15]_i_3_n_3 ;
  wire \pc_reg[3]_i_2_n_0 ;
  wire \pc_reg[3]_i_2_n_1 ;
  wire \pc_reg[3]_i_2_n_2 ;
  wire \pc_reg[3]_i_2_n_3 ;
  wire \pc_reg[7]_i_2_n_0 ;
  wire \pc_reg[7]_i_2_n_1 ;
  wire \pc_reg[7]_i_2_n_2 ;
  wire \pc_reg[7]_i_2_n_3 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [0]),
        .Q(pc[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [10]),
        .Q(pc[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [11]),
        .Q(pc[11]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[11]_i_2 
       (.CI(\pc_reg[7]_i_2_n_0 ),
        .CO({\pc_reg[11]_i_2_n_0 ,\pc_reg[11]_i_2_n_1 ,\pc_reg[11]_i_2_n_2 ,\pc_reg[11]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(fch_pc[11:8]),
        .S(pc[11:8]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [12]),
        .Q(pc[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [13]),
        .Q(pc[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [14]),
        .Q(pc[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [15]),
        .Q(pc[15]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[15]_i_3 
       (.CI(\pc_reg[11]_i_2_n_0 ),
        .CO({\pc_reg[15]_i_3_n_1 ,\pc_reg[15]_i_3_n_2 ,\pc_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(fch_pc[15:12]),
        .S(pc[15:12]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [1]),
        .Q(pc[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [2]),
        .Q(pc[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [3]),
        .Q(pc[3]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[3]_i_2 
       (.CI(\<const0> ),
        .CO({\pc_reg[3]_i_2_n_0 ,\pc_reg[3]_i_2_n_1 ,\pc_reg[3]_i_2_n_2 ,\pc_reg[3]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,pc[1],\<const0> }),
        .O(fch_pc[3:0]),
        .S({pc[3:2],S,pc[0]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [4]),
        .Q(pc[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [5]),
        .Q(pc[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [6]),
        .Q(pc[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [7]),
        .Q(pc[7]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \pc_reg[7]_i_2 
       (.CI(\pc_reg[3]_i_2_n_0 ),
        .CO({\pc_reg[7]_i_2_n_0 ,\pc_reg[7]_i_2_n_1 ,\pc_reg[7]_i_2_n_2 ,\pc_reg[7]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O(fch_pc[7:4]),
        .S(pc[7:4]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [8]),
        .Q(pc[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \pc_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\pc_reg[15]_0 [9]),
        .Q(pc[9]),
        .R(SR));
endmodule

module niho_rgf_sptr
   (.out({sp[31],sp[30],sp[29],sp[28],sp[27],sp[26],sp[25],sp[24],sp[23],sp[22],sp[21],sp[20],sp[19],sp[18],sp[17],sp[16],sp[15],sp[14],sp[13],sp[12],sp[11],sp[10],sp[9],sp[8],sp[7],sp[6],sp[5],sp[4],sp[3],sp[2],sp[1],sp[0]}),
    abus_sp,
    sp_dec_0,
    \sp_reg[1]_0 ,
    \sp_reg[2]_0 ,
    \sp_reg[3]_0 ,
    \sp_reg[4]_0 ,
    \sp_reg[5]_0 ,
    \sp_reg[6]_0 ,
    \sp_reg[7]_0 ,
    \sp_reg[8]_0 ,
    \sp_reg[9]_0 ,
    \sp_reg[10]_0 ,
    \sp_reg[11]_0 ,
    \sp_reg[12]_0 ,
    \sp_reg[13]_0 ,
    \sp_reg[14]_0 ,
    \sp_reg[15]_0 ,
    \sp_reg[16]_0 ,
    \sp_reg[17]_0 ,
    \sp_reg[18]_0 ,
    \sp_reg[19]_0 ,
    \sp_reg[20]_0 ,
    \sp_reg[21]_0 ,
    \sp_reg[22]_0 ,
    \sp_reg[23]_0 ,
    \sp_reg[24]_0 ,
    \sp_reg[25]_0 ,
    \sp_reg[26]_0 ,
    \sp_reg[27]_0 ,
    \sp_reg[28]_0 ,
    \sp_reg[29]_0 ,
    \sp_reg[30]_0 ,
    \sp_reg[31]_0 ,
    O,
    abus_sel_cr,
    ctl_sp_id4,
    ctl_sp_inc,
    ctl_sp_dec,
    SR,
    \sp_reg[31]_1 ,
    clk);
  output [15:0]abus_sp;
  output [30:0]sp_dec_0;
  output \sp_reg[1]_0 ;
  output \sp_reg[2]_0 ;
  output \sp_reg[3]_0 ;
  output \sp_reg[4]_0 ;
  output \sp_reg[5]_0 ;
  output \sp_reg[6]_0 ;
  output \sp_reg[7]_0 ;
  output \sp_reg[8]_0 ;
  output \sp_reg[9]_0 ;
  output \sp_reg[10]_0 ;
  output \sp_reg[11]_0 ;
  output \sp_reg[12]_0 ;
  output \sp_reg[13]_0 ;
  output \sp_reg[14]_0 ;
  output \sp_reg[15]_0 ;
  output \sp_reg[16]_0 ;
  output \sp_reg[17]_0 ;
  output \sp_reg[18]_0 ;
  output \sp_reg[19]_0 ;
  output \sp_reg[20]_0 ;
  output \sp_reg[21]_0 ;
  output \sp_reg[22]_0 ;
  output \sp_reg[23]_0 ;
  output \sp_reg[24]_0 ;
  output \sp_reg[25]_0 ;
  output \sp_reg[26]_0 ;
  output \sp_reg[27]_0 ;
  output \sp_reg[28]_0 ;
  output \sp_reg[29]_0 ;
  output \sp_reg[30]_0 ;
  output \sp_reg[31]_0 ;
  output [0:0]O;
  input [1:0]abus_sel_cr;
  input ctl_sp_id4;
  input ctl_sp_inc;
  input ctl_sp_dec;
  input [0:0]SR;
  input [31:0]\sp_reg[31]_1 ;
  input clk;
     output [31:0]sp;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]O;
  wire [0:0]SR;
  wire [1:0]abus_sel_cr;
  wire [15:0]abus_sp;
  wire \badr[12]_INST_0_i_15_n_0 ;
  wire \badr[12]_INST_0_i_15_n_1 ;
  wire \badr[12]_INST_0_i_15_n_2 ;
  wire \badr[12]_INST_0_i_15_n_3 ;
  wire \badr[12]_INST_0_i_22_n_0 ;
  wire \badr[12]_INST_0_i_23_n_0 ;
  wire \badr[12]_INST_0_i_24_n_0 ;
  wire \badr[12]_INST_0_i_25_n_0 ;
  wire \badr[16]_INST_0_i_12_n_0 ;
  wire \badr[16]_INST_0_i_12_n_1 ;
  wire \badr[16]_INST_0_i_12_n_2 ;
  wire \badr[16]_INST_0_i_12_n_3 ;
  wire \badr[16]_INST_0_i_13_n_0 ;
  wire \badr[16]_INST_0_i_14_n_0 ;
  wire \badr[16]_INST_0_i_15_n_0 ;
  wire \badr[16]_INST_0_i_16_n_0 ;
  wire \badr[20]_INST_0_i_12_n_0 ;
  wire \badr[20]_INST_0_i_12_n_1 ;
  wire \badr[20]_INST_0_i_12_n_2 ;
  wire \badr[20]_INST_0_i_12_n_3 ;
  wire \badr[20]_INST_0_i_13_n_0 ;
  wire \badr[20]_INST_0_i_14_n_0 ;
  wire \badr[20]_INST_0_i_15_n_0 ;
  wire \badr[20]_INST_0_i_16_n_0 ;
  wire \badr[24]_INST_0_i_12_n_0 ;
  wire \badr[24]_INST_0_i_12_n_1 ;
  wire \badr[24]_INST_0_i_12_n_2 ;
  wire \badr[24]_INST_0_i_12_n_3 ;
  wire \badr[24]_INST_0_i_13_n_0 ;
  wire \badr[24]_INST_0_i_14_n_0 ;
  wire \badr[24]_INST_0_i_15_n_0 ;
  wire \badr[24]_INST_0_i_16_n_0 ;
  wire \badr[28]_INST_0_i_12_n_0 ;
  wire \badr[28]_INST_0_i_12_n_1 ;
  wire \badr[28]_INST_0_i_12_n_2 ;
  wire \badr[28]_INST_0_i_12_n_3 ;
  wire \badr[28]_INST_0_i_13_n_0 ;
  wire \badr[28]_INST_0_i_14_n_0 ;
  wire \badr[28]_INST_0_i_15_n_0 ;
  wire \badr[28]_INST_0_i_16_n_0 ;
  wire \badr[31]_INST_0_i_27_n_2 ;
  wire \badr[31]_INST_0_i_27_n_3 ;
  wire \badr[31]_INST_0_i_45_n_0 ;
  wire \badr[31]_INST_0_i_46_n_0 ;
  wire \badr[31]_INST_0_i_47_n_0 ;
  wire \badr[4]_INST_0_i_15_n_0 ;
  wire \badr[4]_INST_0_i_15_n_1 ;
  wire \badr[4]_INST_0_i_15_n_2 ;
  wire \badr[4]_INST_0_i_15_n_3 ;
  wire \badr[4]_INST_0_i_22_n_0 ;
  wire \badr[4]_INST_0_i_23_n_0 ;
  wire \badr[4]_INST_0_i_24_n_0 ;
  wire \badr[4]_INST_0_i_25_n_0 ;
  wire \badr[4]_INST_0_i_26_n_0 ;
  wire \badr[4]_INST_0_i_27_n_0 ;
  wire \badr[8]_INST_0_i_15_n_0 ;
  wire \badr[8]_INST_0_i_15_n_1 ;
  wire \badr[8]_INST_0_i_15_n_2 ;
  wire \badr[8]_INST_0_i_15_n_3 ;
  wire \badr[8]_INST_0_i_22_n_0 ;
  wire \badr[8]_INST_0_i_23_n_0 ;
  wire \badr[8]_INST_0_i_24_n_0 ;
  wire \badr[8]_INST_0_i_25_n_0 ;
  wire clk;
  wire ctl_sp_dec;
  wire ctl_sp_id4;
  wire ctl_sp_inc;
  (* DONT_TOUCH *) wire [31:0]sp;
  wire \sp[0]_i_4_n_0 ;
  wire \sp[0]_i_5_n_0 ;
  wire [30:0]sp_dec_0;
  wire \sp_reg[0]_i_2_n_0 ;
  wire \sp_reg[0]_i_2_n_1 ;
  wire \sp_reg[0]_i_2_n_2 ;
  wire \sp_reg[0]_i_2_n_3 ;
  wire \sp_reg[0]_i_2_n_4 ;
  wire \sp_reg[0]_i_2_n_5 ;
  wire \sp_reg[0]_i_2_n_6 ;
  wire \sp_reg[10]_0 ;
  wire \sp_reg[11]_0 ;
  wire \sp_reg[11]_i_3_n_0 ;
  wire \sp_reg[11]_i_3_n_1 ;
  wire \sp_reg[11]_i_3_n_2 ;
  wire \sp_reg[11]_i_3_n_3 ;
  wire \sp_reg[11]_i_3_n_4 ;
  wire \sp_reg[11]_i_3_n_5 ;
  wire \sp_reg[11]_i_3_n_6 ;
  wire \sp_reg[11]_i_3_n_7 ;
  wire \sp_reg[12]_0 ;
  wire \sp_reg[13]_0 ;
  wire \sp_reg[14]_0 ;
  wire \sp_reg[15]_0 ;
  wire \sp_reg[15]_i_3_n_0 ;
  wire \sp_reg[15]_i_3_n_1 ;
  wire \sp_reg[15]_i_3_n_2 ;
  wire \sp_reg[15]_i_3_n_3 ;
  wire \sp_reg[15]_i_3_n_4 ;
  wire \sp_reg[15]_i_3_n_5 ;
  wire \sp_reg[15]_i_3_n_6 ;
  wire \sp_reg[15]_i_3_n_7 ;
  wire \sp_reg[16]_0 ;
  wire \sp_reg[17]_0 ;
  wire \sp_reg[18]_0 ;
  wire \sp_reg[19]_0 ;
  wire \sp_reg[19]_i_3_n_0 ;
  wire \sp_reg[19]_i_3_n_1 ;
  wire \sp_reg[19]_i_3_n_2 ;
  wire \sp_reg[19]_i_3_n_3 ;
  wire \sp_reg[19]_i_3_n_4 ;
  wire \sp_reg[19]_i_3_n_5 ;
  wire \sp_reg[19]_i_3_n_6 ;
  wire \sp_reg[19]_i_3_n_7 ;
  wire \sp_reg[1]_0 ;
  wire \sp_reg[20]_0 ;
  wire \sp_reg[21]_0 ;
  wire \sp_reg[22]_0 ;
  wire \sp_reg[23]_0 ;
  wire \sp_reg[23]_i_3_n_0 ;
  wire \sp_reg[23]_i_3_n_1 ;
  wire \sp_reg[23]_i_3_n_2 ;
  wire \sp_reg[23]_i_3_n_3 ;
  wire \sp_reg[23]_i_3_n_4 ;
  wire \sp_reg[23]_i_3_n_5 ;
  wire \sp_reg[23]_i_3_n_6 ;
  wire \sp_reg[23]_i_3_n_7 ;
  wire \sp_reg[24]_0 ;
  wire \sp_reg[25]_0 ;
  wire \sp_reg[26]_0 ;
  wire \sp_reg[27]_0 ;
  wire \sp_reg[27]_i_3_n_0 ;
  wire \sp_reg[27]_i_3_n_1 ;
  wire \sp_reg[27]_i_3_n_2 ;
  wire \sp_reg[27]_i_3_n_3 ;
  wire \sp_reg[27]_i_3_n_4 ;
  wire \sp_reg[27]_i_3_n_5 ;
  wire \sp_reg[27]_i_3_n_6 ;
  wire \sp_reg[27]_i_3_n_7 ;
  wire \sp_reg[28]_0 ;
  wire \sp_reg[29]_0 ;
  wire \sp_reg[2]_0 ;
  wire \sp_reg[30]_0 ;
  wire \sp_reg[31]_0 ;
  wire [31:0]\sp_reg[31]_1 ;
  wire \sp_reg[31]_i_4_n_1 ;
  wire \sp_reg[31]_i_4_n_2 ;
  wire \sp_reg[31]_i_4_n_3 ;
  wire \sp_reg[31]_i_4_n_4 ;
  wire \sp_reg[31]_i_4_n_5 ;
  wire \sp_reg[31]_i_4_n_6 ;
  wire \sp_reg[31]_i_4_n_7 ;
  wire \sp_reg[3]_0 ;
  wire \sp_reg[4]_0 ;
  wire \sp_reg[5]_0 ;
  wire \sp_reg[6]_0 ;
  wire \sp_reg[7]_0 ;
  wire \sp_reg[7]_i_3_n_0 ;
  wire \sp_reg[7]_i_3_n_1 ;
  wire \sp_reg[7]_i_3_n_2 ;
  wire \sp_reg[7]_i_3_n_3 ;
  wire \sp_reg[7]_i_3_n_4 ;
  wire \sp_reg[7]_i_3_n_5 ;
  wire \sp_reg[7]_i_3_n_6 ;
  wire \sp_reg[7]_i_3_n_7 ;
  wire \sp_reg[8]_0 ;
  wire \sp_reg[9]_0 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[12]_INST_0_i_15 
       (.CI(\badr[8]_INST_0_i_15_n_0 ),
        .CO({\badr[12]_INST_0_i_15_n_0 ,\badr[12]_INST_0_i_15_n_1 ,\badr[12]_INST_0_i_15_n_2 ,\badr[12]_INST_0_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[11:8]),
        .O(sp_dec_0[11:8]),
        .S({\badr[12]_INST_0_i_22_n_0 ,\badr[12]_INST_0_i_23_n_0 ,\badr[12]_INST_0_i_24_n_0 ,\badr[12]_INST_0_i_25_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_22 
       (.I0(sp[11]),
        .I1(sp[12]),
        .O(\badr[12]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_23 
       (.I0(sp[10]),
        .I1(sp[11]),
        .O(\badr[12]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_24 
       (.I0(sp[9]),
        .I1(sp[10]),
        .O(\badr[12]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[12]_INST_0_i_25 
       (.I0(sp[8]),
        .I1(sp[9]),
        .O(\badr[12]_INST_0_i_25_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[16]_INST_0_i_12 
       (.CI(\badr[12]_INST_0_i_15_n_0 ),
        .CO({\badr[16]_INST_0_i_12_n_0 ,\badr[16]_INST_0_i_12_n_1 ,\badr[16]_INST_0_i_12_n_2 ,\badr[16]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[15:12]),
        .O(sp_dec_0[15:12]),
        .S({\badr[16]_INST_0_i_13_n_0 ,\badr[16]_INST_0_i_14_n_0 ,\badr[16]_INST_0_i_15_n_0 ,\badr[16]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_13 
       (.I0(sp[15]),
        .I1(sp[16]),
        .O(\badr[16]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_14 
       (.I0(sp[14]),
        .I1(sp[15]),
        .O(\badr[16]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_15 
       (.I0(sp[13]),
        .I1(sp[14]),
        .O(\badr[16]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[16]_INST_0_i_16 
       (.I0(sp[12]),
        .I1(sp[13]),
        .O(\badr[16]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[16]_INST_0_i_7 
       (.I0(sp[16]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[15]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[0]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[17]_INST_0_i_7 
       (.I0(sp[17]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[16]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[1]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[18]_INST_0_i_7 
       (.I0(sp[18]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[17]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[2]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[19]_INST_0_i_7 
       (.I0(sp[19]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[18]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[3]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[20]_INST_0_i_12 
       (.CI(\badr[16]_INST_0_i_12_n_0 ),
        .CO({\badr[20]_INST_0_i_12_n_0 ,\badr[20]_INST_0_i_12_n_1 ,\badr[20]_INST_0_i_12_n_2 ,\badr[20]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[19:16]),
        .O(sp_dec_0[19:16]),
        .S({\badr[20]_INST_0_i_13_n_0 ,\badr[20]_INST_0_i_14_n_0 ,\badr[20]_INST_0_i_15_n_0 ,\badr[20]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_13 
       (.I0(sp[19]),
        .I1(sp[20]),
        .O(\badr[20]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_14 
       (.I0(sp[18]),
        .I1(sp[19]),
        .O(\badr[20]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_15 
       (.I0(sp[17]),
        .I1(sp[18]),
        .O(\badr[20]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[20]_INST_0_i_16 
       (.I0(sp[16]),
        .I1(sp[17]),
        .O(\badr[20]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[20]_INST_0_i_7 
       (.I0(sp[20]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[19]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[4]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[21]_INST_0_i_7 
       (.I0(sp[21]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[20]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[5]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[22]_INST_0_i_7 
       (.I0(sp[22]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[21]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[6]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[23]_INST_0_i_7 
       (.I0(sp[23]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[22]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[7]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[24]_INST_0_i_12 
       (.CI(\badr[20]_INST_0_i_12_n_0 ),
        .CO({\badr[24]_INST_0_i_12_n_0 ,\badr[24]_INST_0_i_12_n_1 ,\badr[24]_INST_0_i_12_n_2 ,\badr[24]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[23:20]),
        .O(sp_dec_0[23:20]),
        .S({\badr[24]_INST_0_i_13_n_0 ,\badr[24]_INST_0_i_14_n_0 ,\badr[24]_INST_0_i_15_n_0 ,\badr[24]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_13 
       (.I0(sp[23]),
        .I1(sp[24]),
        .O(\badr[24]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_14 
       (.I0(sp[22]),
        .I1(sp[23]),
        .O(\badr[24]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_15 
       (.I0(sp[21]),
        .I1(sp[22]),
        .O(\badr[24]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[24]_INST_0_i_16 
       (.I0(sp[20]),
        .I1(sp[21]),
        .O(\badr[24]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[24]_INST_0_i_7 
       (.I0(sp[24]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[23]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[8]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[25]_INST_0_i_7 
       (.I0(sp[25]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[24]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[9]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[26]_INST_0_i_7 
       (.I0(sp[26]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[25]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[10]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[27]_INST_0_i_7 
       (.I0(sp[27]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[26]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[11]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[28]_INST_0_i_12 
       (.CI(\badr[24]_INST_0_i_12_n_0 ),
        .CO({\badr[28]_INST_0_i_12_n_0 ,\badr[28]_INST_0_i_12_n_1 ,\badr[28]_INST_0_i_12_n_2 ,\badr[28]_INST_0_i_12_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[27:24]),
        .O(sp_dec_0[27:24]),
        .S({\badr[28]_INST_0_i_13_n_0 ,\badr[28]_INST_0_i_14_n_0 ,\badr[28]_INST_0_i_15_n_0 ,\badr[28]_INST_0_i_16_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_13 
       (.I0(sp[27]),
        .I1(sp[28]),
        .O(\badr[28]_INST_0_i_13_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_14 
       (.I0(sp[26]),
        .I1(sp[27]),
        .O(\badr[28]_INST_0_i_14_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_15 
       (.I0(sp[25]),
        .I1(sp[26]),
        .O(\badr[28]_INST_0_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[28]_INST_0_i_16 
       (.I0(sp[24]),
        .I1(sp[25]),
        .O(\badr[28]_INST_0_i_16_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[28]_INST_0_i_7 
       (.I0(sp[28]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[27]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[12]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[29]_INST_0_i_7 
       (.I0(sp[29]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[28]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[13]));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[30]_INST_0_i_7 
       (.I0(sp[30]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[29]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[14]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[31]_INST_0_i_27 
       (.CI(\badr[28]_INST_0_i_12_n_0 ),
        .CO({\badr[31]_INST_0_i_27_n_2 ,\badr[31]_INST_0_i_27_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,sp[29:28]}),
        .O(sp_dec_0[30:28]),
        .S({\<const0> ,\badr[31]_INST_0_i_45_n_0 ,\badr[31]_INST_0_i_46_n_0 ,\badr[31]_INST_0_i_47_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_45 
       (.I0(sp[30]),
        .I1(sp[31]),
        .O(\badr[31]_INST_0_i_45_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_46 
       (.I0(sp[29]),
        .I1(sp[30]),
        .O(\badr[31]_INST_0_i_46_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[31]_INST_0_i_47 
       (.I0(sp[28]),
        .I1(sp[29]),
        .O(\badr[31]_INST_0_i_47_n_0 ));
  LUT4 #(
    .INIT(16'hF888)) 
    \badr[31]_INST_0_i_8 
       (.I0(sp[31]),
        .I1(abus_sel_cr[0]),
        .I2(sp_dec_0[30]),
        .I3(abus_sel_cr[1]),
        .O(abus_sp[15]));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[4]_INST_0_i_15 
       (.CI(\<const0> ),
        .CO({\badr[4]_INST_0_i_15_n_0 ,\badr[4]_INST_0_i_15_n_1 ,\badr[4]_INST_0_i_15_n_2 ,\badr[4]_INST_0_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI({sp[3],\badr[4]_INST_0_i_22_n_0 ,\badr[4]_INST_0_i_23_n_0 ,\<const0> }),
        .O(sp_dec_0[3:0]),
        .S({\badr[4]_INST_0_i_24_n_0 ,\badr[4]_INST_0_i_25_n_0 ,\badr[4]_INST_0_i_26_n_0 ,\badr[4]_INST_0_i_27_n_0 }));
  LUT2 #(
    .INIT(4'h2)) 
    \badr[4]_INST_0_i_22 
       (.I0(sp[2]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'hE)) 
    \badr[4]_INST_0_i_23 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_24 
       (.I0(sp[3]),
        .I1(sp[4]),
        .O(\badr[4]_INST_0_i_24_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_25 
       (.I0(sp[2]),
        .I1(ctl_sp_id4),
        .I2(sp[3]),
        .O(\badr[4]_INST_0_i_25_n_0 ));
  LUT3 #(
    .INIT(8'h2D)) 
    \badr[4]_INST_0_i_26 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .I2(sp[2]),
        .O(\badr[4]_INST_0_i_26_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[4]_INST_0_i_27 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .O(\badr[4]_INST_0_i_27_n_0 ));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \badr[8]_INST_0_i_15 
       (.CI(\badr[4]_INST_0_i_15_n_0 ),
        .CO({\badr[8]_INST_0_i_15_n_0 ,\badr[8]_INST_0_i_15_n_1 ,\badr[8]_INST_0_i_15_n_2 ,\badr[8]_INST_0_i_15_n_3 }),
        .CYINIT(\<const0> ),
        .DI(sp[7:4]),
        .O(sp_dec_0[7:4]),
        .S({\badr[8]_INST_0_i_22_n_0 ,\badr[8]_INST_0_i_23_n_0 ,\badr[8]_INST_0_i_24_n_0 ,\badr[8]_INST_0_i_25_n_0 }));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_22 
       (.I0(sp[7]),
        .I1(sp[8]),
        .O(\badr[8]_INST_0_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_23 
       (.I0(sp[6]),
        .I1(sp[7]),
        .O(\badr[8]_INST_0_i_23_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_24 
       (.I0(sp[5]),
        .I1(sp[6]),
        .O(\badr[8]_INST_0_i_24_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \badr[8]_INST_0_i_25 
       (.I0(sp[4]),
        .I1(sp[5]),
        .O(\badr[8]_INST_0_i_25_n_0 ));
  LUT2 #(
    .INIT(4'h6)) 
    \sp[0]_i_4 
       (.I0(sp[2]),
        .I1(ctl_sp_id4),
        .O(\sp[0]_i_4_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \sp[0]_i_5 
       (.I0(sp[1]),
        .I1(ctl_sp_id4),
        .O(\sp[0]_i_5_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[10]_i_2 
       (.I0(\sp_reg[11]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[9]),
        .I3(ctl_sp_dec),
        .I4(sp[10]),
        .O(\sp_reg[10]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[11]_i_2 
       (.I0(\sp_reg[11]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[10]),
        .I3(ctl_sp_dec),
        .I4(sp[11]),
        .O(\sp_reg[11]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[12]_i_2 
       (.I0(\sp_reg[15]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[11]),
        .I3(ctl_sp_dec),
        .I4(sp[12]),
        .O(\sp_reg[12]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[13]_i_2 
       (.I0(\sp_reg[15]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[12]),
        .I3(ctl_sp_dec),
        .I4(sp[13]),
        .O(\sp_reg[13]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[14]_i_2 
       (.I0(\sp_reg[15]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[13]),
        .I3(ctl_sp_dec),
        .I4(sp[14]),
        .O(\sp_reg[14]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[15]_i_2 
       (.I0(\sp_reg[15]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[14]),
        .I3(ctl_sp_dec),
        .I4(sp[15]),
        .O(\sp_reg[15]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[16]_i_2 
       (.I0(\sp_reg[19]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[15]),
        .I3(ctl_sp_dec),
        .I4(sp[16]),
        .O(\sp_reg[16]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[17]_i_2 
       (.I0(\sp_reg[19]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[16]),
        .I3(ctl_sp_dec),
        .I4(sp[17]),
        .O(\sp_reg[17]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[18]_i_2 
       (.I0(\sp_reg[19]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[17]),
        .I3(ctl_sp_dec),
        .I4(sp[18]),
        .O(\sp_reg[18]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[19]_i_2 
       (.I0(\sp_reg[19]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[18]),
        .I3(ctl_sp_dec),
        .I4(sp[19]),
        .O(\sp_reg[19]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[1]_i_2 
       (.I0(\sp_reg[0]_i_2_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[0]),
        .I3(ctl_sp_dec),
        .I4(sp[1]),
        .O(\sp_reg[1]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[20]_i_2 
       (.I0(\sp_reg[23]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[19]),
        .I3(ctl_sp_dec),
        .I4(sp[20]),
        .O(\sp_reg[20]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[21]_i_2 
       (.I0(\sp_reg[23]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[20]),
        .I3(ctl_sp_dec),
        .I4(sp[21]),
        .O(\sp_reg[21]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[22]_i_2 
       (.I0(\sp_reg[23]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[21]),
        .I3(ctl_sp_dec),
        .I4(sp[22]),
        .O(\sp_reg[22]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[23]_i_2 
       (.I0(\sp_reg[23]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[22]),
        .I3(ctl_sp_dec),
        .I4(sp[23]),
        .O(\sp_reg[23]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[24]_i_2 
       (.I0(\sp_reg[27]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[23]),
        .I3(ctl_sp_dec),
        .I4(sp[24]),
        .O(\sp_reg[24]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[25]_i_2 
       (.I0(\sp_reg[27]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[24]),
        .I3(ctl_sp_dec),
        .I4(sp[25]),
        .O(\sp_reg[25]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[26]_i_2 
       (.I0(\sp_reg[27]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[25]),
        .I3(ctl_sp_dec),
        .I4(sp[26]),
        .O(\sp_reg[26]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[27]_i_2 
       (.I0(\sp_reg[27]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[26]),
        .I3(ctl_sp_dec),
        .I4(sp[27]),
        .O(\sp_reg[27]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[28]_i_2 
       (.I0(\sp_reg[31]_i_4_n_7 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[27]),
        .I3(ctl_sp_dec),
        .I4(sp[28]),
        .O(\sp_reg[28]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[29]_i_2 
       (.I0(\sp_reg[31]_i_4_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[28]),
        .I3(ctl_sp_dec),
        .I4(sp[29]),
        .O(\sp_reg[29]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[2]_i_2 
       (.I0(\sp_reg[0]_i_2_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[1]),
        .I3(ctl_sp_dec),
        .I4(sp[2]),
        .O(\sp_reg[2]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[30]_i_2 
       (.I0(\sp_reg[31]_i_4_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[29]),
        .I3(ctl_sp_dec),
        .I4(sp[30]),
        .O(\sp_reg[30]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[31]_i_3 
       (.I0(\sp_reg[31]_i_4_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[30]),
        .I3(ctl_sp_dec),
        .I4(sp[31]),
        .O(\sp_reg[31]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[3]_i_2 
       (.I0(\sp_reg[0]_i_2_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[2]),
        .I3(ctl_sp_dec),
        .I4(sp[3]),
        .O(\sp_reg[3]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[4]_i_2 
       (.I0(\sp_reg[7]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[3]),
        .I3(ctl_sp_dec),
        .I4(sp[4]),
        .O(\sp_reg[4]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[5]_i_2 
       (.I0(\sp_reg[7]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[4]),
        .I3(ctl_sp_dec),
        .I4(sp[5]),
        .O(\sp_reg[5]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[6]_i_2 
       (.I0(\sp_reg[7]_i_3_n_5 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[5]),
        .I3(ctl_sp_dec),
        .I4(sp[6]),
        .O(\sp_reg[6]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[7]_i_2 
       (.I0(\sp_reg[7]_i_3_n_4 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[6]),
        .I3(ctl_sp_dec),
        .I4(sp[7]),
        .O(\sp_reg[7]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[8]_i_2 
       (.I0(\sp_reg[11]_i_3_n_7 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[7]),
        .I3(ctl_sp_dec),
        .I4(sp[8]),
        .O(\sp_reg[8]_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sp[9]_i_2 
       (.I0(\sp_reg[11]_i_3_n_6 ),
        .I1(ctl_sp_inc),
        .I2(sp_dec_0[8]),
        .I3(ctl_sp_dec),
        .I4(sp[9]),
        .O(\sp_reg[9]_0 ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [0]),
        .Q(sp[0]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[0]_i_2 
       (.CI(\<const0> ),
        .CO({\sp_reg[0]_i_2_n_0 ,\sp_reg[0]_i_2_n_1 ,\sp_reg[0]_i_2_n_2 ,\sp_reg[0]_i_2_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,sp[2:1],\<const0> }),
        .O({\sp_reg[0]_i_2_n_4 ,\sp_reg[0]_i_2_n_5 ,\sp_reg[0]_i_2_n_6 ,O}),
        .S({sp[3],\sp[0]_i_4_n_0 ,\sp[0]_i_5_n_0 ,sp[0]}));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [10]),
        .Q(sp[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [11]),
        .Q(sp[11]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[11]_i_3 
       (.CI(\sp_reg[7]_i_3_n_0 ),
        .CO({\sp_reg[11]_i_3_n_0 ,\sp_reg[11]_i_3_n_1 ,\sp_reg[11]_i_3_n_2 ,\sp_reg[11]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[11]_i_3_n_4 ,\sp_reg[11]_i_3_n_5 ,\sp_reg[11]_i_3_n_6 ,\sp_reg[11]_i_3_n_7 }),
        .S(sp[11:8]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [12]),
        .Q(sp[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [13]),
        .Q(sp[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [14]),
        .Q(sp[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [15]),
        .Q(sp[15]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[15]_i_3 
       (.CI(\sp_reg[11]_i_3_n_0 ),
        .CO({\sp_reg[15]_i_3_n_0 ,\sp_reg[15]_i_3_n_1 ,\sp_reg[15]_i_3_n_2 ,\sp_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[15]_i_3_n_4 ,\sp_reg[15]_i_3_n_5 ,\sp_reg[15]_i_3_n_6 ,\sp_reg[15]_i_3_n_7 }),
        .S(sp[15:12]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[16] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [16]),
        .Q(sp[16]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[17] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [17]),
        .Q(sp[17]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[18] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [18]),
        .Q(sp[18]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[19] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [19]),
        .Q(sp[19]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[19]_i_3 
       (.CI(\sp_reg[15]_i_3_n_0 ),
        .CO({\sp_reg[19]_i_3_n_0 ,\sp_reg[19]_i_3_n_1 ,\sp_reg[19]_i_3_n_2 ,\sp_reg[19]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[19]_i_3_n_4 ,\sp_reg[19]_i_3_n_5 ,\sp_reg[19]_i_3_n_6 ,\sp_reg[19]_i_3_n_7 }),
        .S(sp[19:16]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [1]),
        .Q(sp[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[20] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [20]),
        .Q(sp[20]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[21] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [21]),
        .Q(sp[21]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[22] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [22]),
        .Q(sp[22]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[23] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [23]),
        .Q(sp[23]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[23]_i_3 
       (.CI(\sp_reg[19]_i_3_n_0 ),
        .CO({\sp_reg[23]_i_3_n_0 ,\sp_reg[23]_i_3_n_1 ,\sp_reg[23]_i_3_n_2 ,\sp_reg[23]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[23]_i_3_n_4 ,\sp_reg[23]_i_3_n_5 ,\sp_reg[23]_i_3_n_6 ,\sp_reg[23]_i_3_n_7 }),
        .S(sp[23:20]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[24] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [24]),
        .Q(sp[24]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[25] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [25]),
        .Q(sp[25]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[26] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [26]),
        .Q(sp[26]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[27] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [27]),
        .Q(sp[27]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[27]_i_3 
       (.CI(\sp_reg[23]_i_3_n_0 ),
        .CO({\sp_reg[27]_i_3_n_0 ,\sp_reg[27]_i_3_n_1 ,\sp_reg[27]_i_3_n_2 ,\sp_reg[27]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[27]_i_3_n_4 ,\sp_reg[27]_i_3_n_5 ,\sp_reg[27]_i_3_n_6 ,\sp_reg[27]_i_3_n_7 }),
        .S(sp[27:24]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[28] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [28]),
        .Q(sp[28]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[29] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [29]),
        .Q(sp[29]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [2]),
        .Q(sp[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[30] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [30]),
        .Q(sp[30]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[31] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [31]),
        .Q(sp[31]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[31]_i_4 
       (.CI(\sp_reg[27]_i_3_n_0 ),
        .CO({\sp_reg[31]_i_4_n_1 ,\sp_reg[31]_i_4_n_2 ,\sp_reg[31]_i_4_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[31]_i_4_n_4 ,\sp_reg[31]_i_4_n_5 ,\sp_reg[31]_i_4_n_6 ,\sp_reg[31]_i_4_n_7 }),
        .S(sp[31:28]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [3]),
        .Q(sp[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [4]),
        .Q(sp[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [5]),
        .Q(sp[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [6]),
        .Q(sp[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [7]),
        .Q(sp[7]),
        .R(SR));
  (* ADDER_THRESHOLD = "35" *) 
  CARRY4 \sp_reg[7]_i_3 
       (.CI(\sp_reg[0]_i_2_n_0 ),
        .CO({\sp_reg[7]_i_3_n_0 ,\sp_reg[7]_i_3_n_1 ,\sp_reg[7]_i_3_n_2 ,\sp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\<const0> }),
        .O({\sp_reg[7]_i_3_n_4 ,\sp_reg[7]_i_3_n_5 ,\sp_reg[7]_i_3_n_6 ,\sp_reg[7]_i_3_n_7 }),
        .S(sp[7:4]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [8]),
        .Q(sp[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sp_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sp_reg[31]_1 [9]),
        .Q(sp[9]),
        .R(SR));
endmodule

module niho_rgf_sreg
   (.out({sr[15],sr[14],sr[13],sr[12],sr[11],sr[10],sr[9],sr[8],sr[7],sr[6],sr[5],sr[4],sr[3],sr[2],sr[1],sr[0]}),
    \sr_reg[1]_0 ,
    \sr_reg[1]_1 ,
    \sr_reg[1]_2 ,
    \sr_reg[1]_3 ,
    \sr_reg[8]_0 ,
    p_2_in,
    \sr_reg[8]_1 ,
    O,
    \sr_reg[8]_2 ,
    \sr_reg[8]_3 ,
    \sr_reg[8]_4 ,
    \sr_reg[8]_5 ,
    \sr_reg[8]_6 ,
    \sr_reg[8]_7 ,
    \sr_reg[8]_8 ,
    \sr_reg[8]_9 ,
    \sr_reg[8]_10 ,
    \sr_reg[8]_11 ,
    alu_sr_flag,
    \sr_reg[8]_12 ,
    \sr_reg[8]_13 ,
    \sr_reg[8]_14 ,
    \iv[11]_i_11_0 ,
    \sr_reg[8]_15 ,
    \iv[13]_i_10_0 ,
    \sr_reg[8]_16 ,
    \iv[10]_i_9 ,
    \sr_reg[8]_17 ,
    \sr_reg[8]_18 ,
    \sr_reg[8]_19 ,
    \sr_reg[8]_20 ,
    \sr_reg[8]_21 ,
    \sr_reg[8]_22 ,
    \iv[14]_i_11_0 ,
    \sr_reg[8]_23 ,
    \sr_reg[8]_24 ,
    \sr_reg[8]_25 ,
    \sr_reg[8]_26 ,
    \sr_reg[8]_27 ,
    \sr_reg[8]_28 ,
    \sr_reg[8]_29 ,
    \sr_reg[8]_30 ,
    \iv[4]_i_35_0 ,
    \sr_reg[8]_31 ,
    \sr_reg[8]_32 ,
    \sr_reg[8]_33 ,
    \sr_reg[8]_34 ,
    \sr_reg[8]_35 ,
    \iv[3]_i_41_0 ,
    \sr_reg[8]_36 ,
    \iv[10]_i_41_0 ,
    \sr_reg[8]_37 ,
    \iv[9]_i_46_0 ,
    \sr_reg[8]_38 ,
    \sr_reg[8]_39 ,
    \sr_reg[8]_40 ,
    \sr_reg[8]_41 ,
    \sr_reg[8]_42 ,
    \sr_reg[8]_43 ,
    \sr_reg[8]_44 ,
    \sr_reg[8]_45 ,
    \sr_reg[8]_46 ,
    \sr_reg[8]_47 ,
    \sr_reg[8]_48 ,
    \sr_reg[8]_49 ,
    \sr_reg[8]_50 ,
    \sr_reg[8]_51 ,
    \iv[8]_i_34 ,
    \sr_reg[8]_52 ,
    \sr_reg[8]_53 ,
    \sr_reg[8]_54 ,
    \sr_reg[8]_55 ,
    \sr_reg[8]_56 ,
    \sr_reg[8]_57 ,
    \sr_reg[8]_58 ,
    \sr_reg[8]_59 ,
    \sr_reg[8]_60 ,
    \sr_reg[8]_61 ,
    \sr_reg[8]_62 ,
    \sr_reg[8]_63 ,
    \sr_reg[8]_64 ,
    \sr_reg[8]_65 ,
    \sr_reg[8]_66 ,
    \sr_reg[8]_67 ,
    \sr_reg[8]_68 ,
    \sr_reg[8]_69 ,
    \sr_reg[8]_70 ,
    \sr_reg[8]_71 ,
    \sr_reg[8]_72 ,
    \sr_reg[8]_73 ,
    \sr_reg[8]_74 ,
    \sr_reg[8]_75 ,
    \iv[13]_i_35 ,
    \badr[16]_INST_0_i_1 ,
    \iv[13]_i_50 ,
    \sr_reg[8]_76 ,
    \sr_reg[8]_77 ,
    \sr_reg[8]_78 ,
    \sr_reg[8]_79 ,
    \sr_reg[8]_80 ,
    \iv[10]_i_34 ,
    \iv[10]_i_44_0 ,
    \sr_reg[8]_81 ,
    \sr_reg[8]_82 ,
    \sr_reg[8]_83 ,
    \sr_reg[8]_84 ,
    \sr_reg[8]_85 ,
    \sr_reg[8]_86 ,
    \sr_reg[8]_87 ,
    \sr_reg[8]_88 ,
    \sr_reg[6]_0 ,
    \sr_reg[6]_1 ,
    \badr[18]_INST_0_i_1 ,
    \sr_reg[8]_89 ,
    \sr_reg[8]_90 ,
    \sr_reg[8]_91 ,
    \sr_reg[8]_92 ,
    \sr_reg[8]_93 ,
    \sr_reg[8]_94 ,
    \sr_reg[8]_95 ,
    \iv[0]_i_31_0 ,
    \sr_reg[6]_2 ,
    \sr_reg[8]_96 ,
    \sr_reg[8]_97 ,
    \iv[12]_i_49 ,
    \sr_reg[8]_98 ,
    \sr_reg[8]_99 ,
    \sr_reg[8]_100 ,
    \iv[8]_i_38 ,
    \badr[16]_INST_0_i_1_0 ,
    \sr_reg[8]_101 ,
    \sr_reg[8]_102 ,
    \sr_reg[8]_103 ,
    \sr_reg[8]_104 ,
    \sr_reg[8]_105 ,
    \badr[17]_INST_0_i_1 ,
    \sr_reg[8]_106 ,
    \sr_reg[8]_107 ,
    \iv[14]_i_30_0 ,
    \sr_reg[8]_108 ,
    \sr_reg[8]_109 ,
    \sr_reg[8]_110 ,
    niho_dsp_a,
    \sr_reg[8]_111 ,
    \sr_reg[8]_112 ,
    \sr_reg[8]_113 ,
    \sr_reg[8]_114 ,
    \sr_reg[8]_115 ,
    \sr_reg[8]_116 ,
    \badr[5]_INST_0_i_1 ,
    \sr_reg[8]_117 ,
    \sr_reg[8]_118 ,
    \sr_reg[8]_119 ,
    \badr[1]_INST_0_i_1 ,
    \sr_reg[8]_120 ,
    \badr[0]_INST_0_i_1 ,
    \iv[15]_i_108 ,
    mul_a_i,
    \iv[15]_i_108_0 ,
    \iv[15]_i_108_1 ,
    \iv[15]_i_108_2 ,
    \iv[15]_i_108_3 ,
    \iv[15]_i_108_4 ,
    \iv[15]_i_108_5 ,
    \iv[15]_i_108_6 ,
    \iv[15]_i_108_7 ,
    \iv[15]_i_108_8 ,
    \iv[15]_i_108_9 ,
    \iv[15]_i_108_10 ,
    \iv[15]_i_108_11 ,
    \iv[15]_i_108_12 ,
    \sr_reg[8]_121 ,
    \iv[15]_i_108_13 ,
    mul_rslt0,
    \quo_reg[19] ,
    \rem_reg[21] ,
    \quo_reg[23] ,
    \quo_reg[27] ,
    \rem_reg[28] ,
    \rem_reg[29] ,
    \sr_reg[8]_122 ,
    \sr_reg[8]_123 ,
    \sr_reg[8]_124 ,
    \sr_reg[8]_125 ,
    \sr_reg[8]_126 ,
    \sr_reg[8]_127 ,
    \sr_reg[8]_128 ,
    \sr_reg[8]_129 ,
    \sr_reg[8]_130 ,
    \sr_reg[8]_131 ,
    abus_o,
    fch_irq_req,
    .irq_lev_0_sp_1(irq_lev_0_sn_1),
    \sr_reg[7]_0 ,
    \sr_reg[5]_0 ,
    \sr_reg[7]_1 ,
    \sr_reg[4]_0 ,
    \sr_reg[7]_2 ,
    \sr_reg[4]_1 ,
    \sr_reg[6]_3 ,
    \sr_reg[7]_3 ,
    \sr_reg[8]_132 ,
    S,
    \sr_reg[8]_133 ,
    \sr_reg[8]_134 ,
    \sr_reg[8]_135 ,
    \sr_reg[8]_136 ,
    \sr_reg[8]_137 ,
    \sr_reg[8]_138 ,
    \sr_reg[8]_139 ,
    \sr_reg[8]_140 ,
    \sr_reg[8]_141 ,
    \sr_reg[8]_142 ,
    \sr_reg[8]_143 ,
    \sr_reg[8]_144 ,
    \sr_reg[8]_145 ,
    \sr_reg[1]_4 ,
    \sr_reg[1]_5 ,
    \stat_reg[0] ,
    .irq_lev_1_sp_1(irq_lev_1_sn_1),
    \sr_reg[5]_1 ,
    \sr_reg[0]_0 ,
    E,
    \sr_reg[1]_6 ,
    \sr_reg[1]_7 ,
    \sr_reg[1]_8 ,
    \sr_reg[0]_1 ,
    \sr_reg[0]_2 ,
    \sr_reg[0]_3 ,
    \sr_reg[0]_4 ,
    \sr_reg[0]_5 ,
    \sr_reg[0]_6 ,
    \sr_reg[0]_7 ,
    \sr_reg[0]_8 ,
    \sr_reg[0]_9 ,
    \sr_reg[0]_10 ,
    \sr_reg[0]_11 ,
    \sr_reg[0]_12 ,
    \sr_reg[0]_13 ,
    \sr_reg[0]_14 ,
    \sr_reg[0]_15 ,
    \sr_reg[0]_16 ,
    \sr_reg[0]_17 ,
    \sr_reg[0]_18 ,
    \sr_reg[0]_19 ,
    \sr_reg[0]_20 ,
    \sr_reg[0]_21 ,
    \sr_reg[0]_22 ,
    \sr_reg[0]_23 ,
    \sr_reg[0]_24 ,
    \sr_reg[0]_25 ,
    \sr_reg[0]_26 ,
    \sr_reg[0]_27 ,
    \sr_reg[0]_28 ,
    \sr_reg[0]_29 ,
    \sr_reg[0]_30 ,
    \sr_reg[0]_31 ,
    \sr_reg[0]_32 ,
    \sr_reg[0]_33 ,
    \sr_reg[0]_34 ,
    \sr_reg[0]_35 ,
    \sr_reg[0]_36 ,
    \sr_reg[0]_37 ,
    \sr_reg[0]_38 ,
    \sr_reg[0]_39 ,
    \sr_reg[0]_40 ,
    \sr_reg[0]_41 ,
    \sr_reg[0]_42 ,
    \sr_reg[0]_43 ,
    \sr_reg[0]_44 ,
    \sr_reg[0]_45 ,
    \sr_reg[0]_46 ,
    \sr_reg[0]_47 ,
    \sr_reg[0]_48 ,
    \sr_reg[0]_49 ,
    \sr_reg[0]_50 ,
    \sr_reg[0]_51 ,
    \sr_reg[0]_52 ,
    \sr_reg[0]_53 ,
    \sr_reg[0]_54 ,
    \sr_reg[0]_55 ,
    \sr_reg[0]_56 ,
    \sr_reg[0]_57 ,
    \sr_reg[0]_58 ,
    \sr_reg[0]_59 ,
    \sr_reg[0]_60 ,
    \sr_reg[0]_61 ,
    \sr_reg[0]_62 ,
    \sr_reg[0]_63 ,
    \sr_reg[0]_64 ,
    \sr_reg[0]_65 ,
    \sr_reg[0]_66 ,
    \sr_reg[0]_67 ,
    \sr_reg[0]_68 ,
    \sr_reg[0]_69 ,
    \sr_reg[0]_70 ,
    \sr_reg[0]_71 ,
    \sr_reg[0]_72 ,
    \sr_reg[0]_73 ,
    \sr_reg[0]_74 ,
    \sr_reg[0]_75 ,
    \sr_reg[0]_76 ,
    \sr_reg[0]_77 ,
    \sr_reg[0]_78 ,
    \sr_reg[0]_79 ,
    \sr_reg[0]_80 ,
    \sr_reg[0]_81 ,
    \sr_reg[0]_82 ,
    \sr_reg[0]_83 ,
    \sr_reg[0]_84 ,
    \sr_reg[0]_85 ,
    \sr_reg[0]_86 ,
    \sr_reg[0]_87 ,
    \sr_reg[0]_88 ,
    \sr_reg[0]_89 ,
    \sr_reg[0]_90 ,
    \sr_reg[0]_91 ,
    \sr_reg[0]_92 ,
    \sr_reg[0]_93 ,
    \sr_reg[0]_94 ,
    \sr_reg[0]_95 ,
    \sr_reg[0]_96 ,
    \sr_reg[8]_146 ,
    \sr_reg[8]_147 ,
    \sr_reg[8]_148 ,
    \sr_reg[8]_149 ,
    \sr_reg[8]_150 ,
    \sr_reg[8]_151 ,
    \sr_reg[8]_152 ,
    \sr_reg[8]_153 ,
    \sr_reg[8]_154 ,
    \sr_reg[8]_155 ,
    \sr_reg[8]_156 ,
    \sr_reg[8]_157 ,
    \sr_reg[8]_158 ,
    \sr_reg[8]_159 ,
    \sr_reg[8]_160 ,
    \sr_reg[8]_161 ,
    \sr_reg[8]_162 ,
    \sr_reg[8]_163 ,
    \sr_reg[8]_164 ,
    \sr_reg[8]_165 ,
    \sr_reg[8]_166 ,
    \sr_reg[8]_167 ,
    \sr_reg[8]_168 ,
    \sr_reg[8]_169 ,
    \sr_reg[8]_170 ,
    \sr_reg[8]_171 ,
    \sr_reg[8]_172 ,
    \sr_reg[8]_173 ,
    \sr_reg[8]_174 ,
    \sr_reg[8]_175 ,
    \sr_reg[8]_176 ,
    \sr_reg[8]_177 ,
    \sr_reg[8]_178 ,
    \sr_reg[8]_179 ,
    \sr_reg[8]_180 ,
    \sr_reg[8]_181 ,
    \sr_reg[8]_182 ,
    \sr_reg[8]_183 ,
    \sr_reg[8]_184 ,
    \sr_reg[8]_185 ,
    \sr_reg[8]_186 ,
    \sr_reg[8]_187 ,
    \sr_reg[8]_188 ,
    \sr_reg[8]_189 ,
    \sr_reg[8]_190 ,
    \sr_reg[8]_191 ,
    \sr_reg[8]_192 ,
    \sr_reg[8]_193 ,
    \sr_reg[8]_194 ,
    \sr_reg[8]_195 ,
    \sr_reg[8]_196 ,
    \sr_reg[8]_197 ,
    \sr_reg[8]_198 ,
    \sr_reg[8]_199 ,
    \sr_reg[8]_200 ,
    \sr_reg[8]_201 ,
    \sr_reg[8]_202 ,
    \sr_reg[8]_203 ,
    \sr_reg[8]_204 ,
    \sr_reg[8]_205 ,
    \sr_reg[8]_206 ,
    \sr_reg[8]_207 ,
    \sr_reg[8]_208 ,
    \sr_reg[8]_209 ,
    \sr_reg[8]_210 ,
    \sr_reg[8]_211 ,
    \sr_reg[8]_212 ,
    \sr_reg[8]_213 ,
    \sr_reg[8]_214 ,
    \sr_reg[8]_215 ,
    \sr_reg[8]_216 ,
    \sr_reg[8]_217 ,
    \sr_reg[8]_218 ,
    \sr_reg[8]_219 ,
    \sr_reg[8]_220 ,
    \badr[6]_INST_0_i_1 ,
    \sr_reg[8]_221 ,
    \badr[4]_INST_0_i_1 ,
    \sr[6]_i_13 ,
    \sr_reg[8]_222 ,
    \sr_reg[8]_223 ,
    \badr[2]_INST_0_i_1 ,
    niho_dsp_b,
    \sr_reg[8]_224 ,
    \sr_reg[8]_225 ,
    \sr_reg[8]_226 ,
    \sr_reg[8]_227 ,
    rst_n,
    \sr_reg[15]_0 ,
    cbus_sel_0,
    \sr_reg[5]_2 ,
    \sr_reg[5]_3 ,
    \sr_reg[6]_4 ,
    \tr_reg[31] ,
    \tr_reg[31]_0 ,
    \sr[4]_i_19 ,
    \sr[4]_i_19_0 ,
    \sr[4]_i_19_1 ,
    \iv[6]_i_3 ,
    \niho_dsp_b[5] ,
    \sr[4]_i_38 ,
    \sr[4]_i_38_0 ,
    \sr[4]_i_91 ,
    \tr[23]_i_3 ,
    \tr[28]_i_3 ,
    \sr_reg[6]_5 ,
    \sr[5]_i_3 ,
    \sr[5]_i_3_0 ,
    \sr[5]_i_3_1 ,
    \sr[5]_i_3_2 ,
    \sr[5]_i_3_3 ,
    \sr[5]_i_3_4 ,
    \sr[5]_i_3_5 ,
    \mul_a_reg[32] ,
    \sr[4]_i_42_0 ,
    \sr[4]_i_42_1 ,
    \sr[4]_i_43 ,
    \iv[11]_i_4_0 ,
    \iv[13]_i_4_0 ,
    \iv[13]_i_4_1 ,
    \iv[0]_i_3 ,
    \iv[0]_i_3_0 ,
    \iv[0]_i_3_1 ,
    \sr[4]_i_17 ,
    \sr[4]_i_34 ,
    \iv[5]_i_3 ,
    \iv[4]_i_3 ,
    \sr[4]_i_32 ,
    \sr[4]_i_39 ,
    \iv[14]_i_2 ,
    \sr[4]_i_40 ,
    \sr[4]_i_37 ,
    \iv[6]_i_8 ,
    \iv[9]_i_4 ,
    \iv[8]_i_4 ,
    \iv[10]_i_4 ,
    \iv[3]_i_8 ,
    \iv[2]_i_8 ,
    \iv[1]_i_8 ,
    \iv[7]_i_8 ,
    \tr[16]_i_2 ,
    \tr[16]_i_2_0 ,
    \iv[15]_i_8 ,
    bbus_0,
    \sr[6]_i_4_0 ,
    \sr[6]_i_4_1 ,
    \sr[6]_i_4_2 ,
    \sr[6]_i_11_0 ,
    \sr[6]_i_11_1 ,
    \iv[0]_i_21 ,
    \iv[15]_i_8_0 ,
    \iv[15]_i_8_1 ,
    \iv[15]_i_8_2 ,
    \sr[4]_i_42_2 ,
    \sr[4]_i_42_3 ,
    \sr[4]_i_91_0 ,
    \iv[10]_i_6 ,
    \sr[4]_i_74 ,
    \sr[4]_i_66 ,
    \tr[27]_i_9 ,
    \sr[4]_i_73 ,
    \sr[4]_i_69_0 ,
    \sr[4]_i_103 ,
    \sr[4]_i_86 ,
    \sr[4]_i_94_0 ,
    \sr[4]_i_87_0 ,
    \sr[4]_i_90_0 ,
    \iv[6]_i_10 ,
    \tr[21]_i_9 ,
    \iv[9]_i_28 ,
    \iv[4]_i_27_0 ,
    \tr[28]_i_8_0 ,
    \tr[21]_i_8 ,
    \mul_a_reg[30] ,
    .niho_dsp_b_0_sp_1(niho_dsp_b_0_sn_1),
    \tr[26]_i_6 ,
    \iv[10]_i_29_0 ,
    \iv[14]_i_13 ,
    \iv[9]_i_28_0 ,
    \iv[5]_i_15 ,
    \iv[15]_i_58 ,
    \tr[23]_i_6 ,
    \tr[23]_i_6_0 ,
    \tr[19]_i_6 ,
    \iv[8]_i_27 ,
    \iv[12]_i_25 ,
    \tr[20]_i_8 ,
    \tr[24]_i_9 ,
    \mul_a_reg[29] ,
    \sr[6]_i_38_0 ,
    \sr[6]_i_10 ,
    \sr[4]_i_139_0 ,
    \mul_a_reg[22] ,
    \mul_a_reg[21] ,
    \mul_a_reg[20] ,
    \mul_a_reg[19] ,
    \iv[15]_i_96 ,
    \iv[15]_i_96_0 ,
    \iv[15]_i_96_1 ,
    \iv[15]_i_96_2 ,
    \iv[15]_i_96_3 ,
    \iv[15]_i_96_4 ,
    \iv[15]_i_96_5 ,
    \iv[15]_i_96_6 ,
    \iv[15]_i_96_7 ,
    \iv[15]_i_96_8 ,
    \iv[13]_i_45_0 ,
    \iv[13]_i_45_1 ,
    \iv[10]_i_44_1 ,
    \iv[10]_i_44_2 ,
    \mul_a_reg[28] ,
    \mul_a_reg[27] ,
    \mul_a_reg[26] ,
    \mul_a_reg[25] ,
    \mul_a_reg[24] ,
    \mul_a_reg[23] ,
    \mul_a_reg[18] ,
    \mul_a_reg[17] ,
    \mul_a_reg[16] ,
    mul_rslt,
    mul_a,
    \niho_dsp_b[5]_0 ,
    .niho_dsp_a_15_sp_1(niho_dsp_a_15_sn_1),
    \remden_reg[26] ,
    DI,
    \remden_reg[29] ,
    \niho_dsp_a[11] ,
    \remden_reg[25] ,
    \remden_reg[24] ,
    \niho_dsp_a[7] ,
    \remden_reg[23] ,
    \remden_reg[22] ,
    \remden_reg[21] ,
    \iv[5]_i_7 ,
    \remden_reg[20] ,
    \niho_dsp_a[3] ,
    \remden_reg[18] ,
    \remden_reg[17] ,
    \remden_reg[16] ,
    \tr[23]_i_5 ,
    Q,
    \tr[19]_i_2 ,
    \tr[29]_i_2 ,
    \tr[19]_i_2_0 ,
    \sr[4]_i_3 ,
    \sr[4]_i_3_0 ,
    CO,
    \abus_o[16] ,
    irq,
    irq_lev,
    \badr[31]_INST_0_i_69 ,
    \stat_reg[1] ,
    \stat[0]_i_6 ,
    \pc_reg[3]_i_2 ,
    \sr[4]_i_42_4 ,
    \sr[4]_i_42_5 ,
    \sr[4]_i_42_6 ,
    \sr[4]_i_41 ,
    \sr[4]_i_41_0 ,
    \sr[4]_i_47 ,
    \sr[4]_i_47_0 ,
    \sr[4]_i_46 ,
    \sr[4]_i_46_0 ,
    \sr[4]_i_35 ,
    \sr[4]_i_35_0 ,
    \sr[4]_i_33 ,
    \sr[4]_i_33_0 ,
    \sr[4]_i_31 ,
    \sr[4]_i_31_0 ,
    \sr[4]_i_39_0 ,
    \sr[4]_i_39_1 ,
    \sr[4]_i_40_0 ,
    \sr[4]_i_40_1 ,
    \sr[4]_i_37_0 ,
    \sr[4]_i_37_1 ,
    \grn_reg[0] ,
    \grn_reg[0]_0 ,
    bbus_sel_0,
    \bdatw[31]_INST_0_i_4 ,
    \bdatw[31]_INST_0_i_4_0 ,
    \i_/badr[31]_INST_0_i_5 ,
    \i_/badr[31]_INST_0_i_5_0 ,
    \bdatw[31]_INST_0_i_4_1 ,
    \bdatw[31]_INST_0_i_4_2 ,
    \i_/badr[31]_INST_0_i_4 ,
    \i_/badr[31]_INST_0_i_4_0 ,
    \i_/badr[31]_INST_0_i_7 ,
    \i_/badr[31]_INST_0_i_7_0 ,
    \i_/badr[31]_INST_0_i_6 ,
    \i_/badr[31]_INST_0_i_6_0 ,
    abus_sel_0,
    \tr[30]_i_10 ,
    \tr[21]_i_9_0 ,
    \tr[21]_i_9_1 ,
    \tr[26]_i_7 ,
    \tr[26]_i_7_0 ,
    \tr[25]_i_9 ,
    \tr[19]_i_7 ,
    \tr[28]_i_9 ,
    \tr[23]_i_7 ,
    \tr[27]_i_7 ,
    \tr[18]_i_9 ,
    \tr[22]_i_9 ,
    \remden_reg[19] ,
    \sr[5]_i_2_0 ,
    \mul_a_reg[32]_0 ,
    \sr[6]_i_4_3 ,
    \tr_reg[31]_i_13_0 ,
    \remden_reg[30] ,
    \tr_reg[31]_i_13_1 ,
    \tr_reg[31]_i_13_2 ,
    \remden_reg[28] ,
    \tr_reg[31]_i_32_0 ,
    \remden_reg[27] ,
    \tr_reg[31]_i_32_1 ,
    \remden_reg[26]_0 ,
    \tr_reg[31]_i_32_2 ,
    \tr_reg[31]_i_32_3 ,
    \tr_reg[23]_i_11_0 ,
    \tr_reg[23]_i_11_1 ,
    \tr_reg[23]_i_11_2 ,
    \tr_reg[23]_i_11_3 ,
    \sr_reg[6]_i_6_0 ,
    \sr_reg[6]_i_6_1 ,
    \sr_reg[6]_i_6_2 ,
    \niho_dsp_b[0]_0 ,
    \niho_dsp_b[5]_1 ,
    \iv[11]_i_10_0 ,
    \iv[12]_i_9 ,
    \tr[20]_i_9 ,
    clk,
    D,
    SR,
    \sr_reg[11]_0 ,
    \sr_reg[10]_0 ,
    \sr_reg[8]_228 ,
    \sr_reg[7]_4 ,
    \sr_reg[6]_6 ,
    \sr_reg[5]_4 ,
    \sr_reg[4]_2 ,
    \sr_reg[3]_0 ,
    \sr_reg[2]_0 ,
    \sr_reg[1]_9 ,
    \sr_reg[0]_97 );
  output [0:0]\sr_reg[1]_0 ;
  output [0:0]\sr_reg[1]_1 ;
  output [0:0]\sr_reg[1]_2 ;
  output [0:0]\sr_reg[1]_3 ;
  output \sr_reg[8]_0 ;
  output [0:0]p_2_in;
  output \sr_reg[8]_1 ;
  output [0:0]O;
  output \sr_reg[8]_2 ;
  output \sr_reg[8]_3 ;
  output \sr_reg[8]_4 ;
  output \sr_reg[8]_5 ;
  output \sr_reg[8]_6 ;
  output \sr_reg[8]_7 ;
  output \sr_reg[8]_8 ;
  output \sr_reg[8]_9 ;
  output \sr_reg[8]_10 ;
  output \sr_reg[8]_11 ;
  output [0:0]alu_sr_flag;
  output \sr_reg[8]_12 ;
  output \sr_reg[8]_13 ;
  output \sr_reg[8]_14 ;
  output \iv[11]_i_11_0 ;
  output \sr_reg[8]_15 ;
  output \iv[13]_i_10_0 ;
  output \sr_reg[8]_16 ;
  output \iv[10]_i_9 ;
  output \sr_reg[8]_17 ;
  output \sr_reg[8]_18 ;
  output \sr_reg[8]_19 ;
  output \sr_reg[8]_20 ;
  output \sr_reg[8]_21 ;
  output \sr_reg[8]_22 ;
  output \iv[14]_i_11_0 ;
  output \sr_reg[8]_23 ;
  output \sr_reg[8]_24 ;
  output \sr_reg[8]_25 ;
  output \sr_reg[8]_26 ;
  output \sr_reg[8]_27 ;
  output \sr_reg[8]_28 ;
  output \sr_reg[8]_29 ;
  output \sr_reg[8]_30 ;
  output \iv[4]_i_35_0 ;
  output \sr_reg[8]_31 ;
  output \sr_reg[8]_32 ;
  output \sr_reg[8]_33 ;
  output \sr_reg[8]_34 ;
  output \sr_reg[8]_35 ;
  output \iv[3]_i_41_0 ;
  output \sr_reg[8]_36 ;
  output \iv[10]_i_41_0 ;
  output \sr_reg[8]_37 ;
  output \iv[9]_i_46_0 ;
  output \sr_reg[8]_38 ;
  output \sr_reg[8]_39 ;
  output \sr_reg[8]_40 ;
  output \sr_reg[8]_41 ;
  output \sr_reg[8]_42 ;
  output \sr_reg[8]_43 ;
  output \sr_reg[8]_44 ;
  output \sr_reg[8]_45 ;
  output \sr_reg[8]_46 ;
  output \sr_reg[8]_47 ;
  output \sr_reg[8]_48 ;
  output \sr_reg[8]_49 ;
  output \sr_reg[8]_50 ;
  output \sr_reg[8]_51 ;
  output \iv[8]_i_34 ;
  output \sr_reg[8]_52 ;
  output \sr_reg[8]_53 ;
  output \sr_reg[8]_54 ;
  output \sr_reg[8]_55 ;
  output \sr_reg[8]_56 ;
  output \sr_reg[8]_57 ;
  output \sr_reg[8]_58 ;
  output \sr_reg[8]_59 ;
  output \sr_reg[8]_60 ;
  output \sr_reg[8]_61 ;
  output \sr_reg[8]_62 ;
  output \sr_reg[8]_63 ;
  output \sr_reg[8]_64 ;
  output \sr_reg[8]_65 ;
  output \sr_reg[8]_66 ;
  output \sr_reg[8]_67 ;
  output \sr_reg[8]_68 ;
  output \sr_reg[8]_69 ;
  output \sr_reg[8]_70 ;
  output \sr_reg[8]_71 ;
  output \sr_reg[8]_72 ;
  output \sr_reg[8]_73 ;
  output \sr_reg[8]_74 ;
  output \sr_reg[8]_75 ;
  output \iv[13]_i_35 ;
  output \badr[16]_INST_0_i_1 ;
  output \iv[13]_i_50 ;
  output \sr_reg[8]_76 ;
  output \sr_reg[8]_77 ;
  output \sr_reg[8]_78 ;
  output \sr_reg[8]_79 ;
  output \sr_reg[8]_80 ;
  output \iv[10]_i_34 ;
  output \iv[10]_i_44_0 ;
  output \sr_reg[8]_81 ;
  output \sr_reg[8]_82 ;
  output \sr_reg[8]_83 ;
  output \sr_reg[8]_84 ;
  output \sr_reg[8]_85 ;
  output \sr_reg[8]_86 ;
  output \sr_reg[8]_87 ;
  output \sr_reg[8]_88 ;
  output \sr_reg[6]_0 ;
  output \sr_reg[6]_1 ;
  output \badr[18]_INST_0_i_1 ;
  output \sr_reg[8]_89 ;
  output \sr_reg[8]_90 ;
  output \sr_reg[8]_91 ;
  output \sr_reg[8]_92 ;
  output \sr_reg[8]_93 ;
  output \sr_reg[8]_94 ;
  output \sr_reg[8]_95 ;
  output \iv[0]_i_31_0 ;
  output \sr_reg[6]_2 ;
  output \sr_reg[8]_96 ;
  output \sr_reg[8]_97 ;
  output \iv[12]_i_49 ;
  output \sr_reg[8]_98 ;
  output \sr_reg[8]_99 ;
  output \sr_reg[8]_100 ;
  output \iv[8]_i_38 ;
  output \badr[16]_INST_0_i_1_0 ;
  output \sr_reg[8]_101 ;
  output \sr_reg[8]_102 ;
  output \sr_reg[8]_103 ;
  output \sr_reg[8]_104 ;
  output \sr_reg[8]_105 ;
  output \badr[17]_INST_0_i_1 ;
  output \sr_reg[8]_106 ;
  output \sr_reg[8]_107 ;
  output \iv[14]_i_30_0 ;
  output \sr_reg[8]_108 ;
  output \sr_reg[8]_109 ;
  output \sr_reg[8]_110 ;
  output [15:0]niho_dsp_a;
  output \sr_reg[8]_111 ;
  output \sr_reg[8]_112 ;
  output \sr_reg[8]_113 ;
  output \sr_reg[8]_114 ;
  output \sr_reg[8]_115 ;
  output \sr_reg[8]_116 ;
  output \badr[5]_INST_0_i_1 ;
  output \sr_reg[8]_117 ;
  output \sr_reg[8]_118 ;
  output \sr_reg[8]_119 ;
  output \badr[1]_INST_0_i_1 ;
  output \sr_reg[8]_120 ;
  output \badr[0]_INST_0_i_1 ;
  output \iv[15]_i_108 ;
  output [13:0]mul_a_i;
  output \iv[15]_i_108_0 ;
  output \iv[15]_i_108_1 ;
  output \iv[15]_i_108_2 ;
  output \iv[15]_i_108_3 ;
  output \iv[15]_i_108_4 ;
  output \iv[15]_i_108_5 ;
  output \iv[15]_i_108_6 ;
  output \iv[15]_i_108_7 ;
  output \iv[15]_i_108_8 ;
  output \iv[15]_i_108_9 ;
  output \iv[15]_i_108_10 ;
  output \iv[15]_i_108_11 ;
  output \iv[15]_i_108_12 ;
  output \sr_reg[8]_121 ;
  output \iv[15]_i_108_13 ;
  output mul_rslt0;
  output \quo_reg[19] ;
  output \rem_reg[21] ;
  output \quo_reg[23] ;
  output \quo_reg[27] ;
  output \rem_reg[28] ;
  output \rem_reg[29] ;
  output \sr_reg[8]_122 ;
  output \sr_reg[8]_123 ;
  output \sr_reg[8]_124 ;
  output \sr_reg[8]_125 ;
  output \sr_reg[8]_126 ;
  output \sr_reg[8]_127 ;
  output \sr_reg[8]_128 ;
  output \sr_reg[8]_129 ;
  output \sr_reg[8]_130 ;
  output \sr_reg[8]_131 ;
  output [15:0]abus_o;
  output fch_irq_req;
  output \sr_reg[7]_0 ;
  output \sr_reg[5]_0 ;
  output \sr_reg[7]_1 ;
  output \sr_reg[4]_0 ;
  output \sr_reg[7]_2 ;
  output \sr_reg[4]_1 ;
  output \sr_reg[6]_3 ;
  output \sr_reg[7]_3 ;
  output \sr_reg[8]_132 ;
  output [0:0]S;
  output \sr_reg[8]_133 ;
  output \sr_reg[8]_134 ;
  output \sr_reg[8]_135 ;
  output \sr_reg[8]_136 ;
  output \sr_reg[8]_137 ;
  output \sr_reg[8]_138 ;
  output \sr_reg[8]_139 ;
  output \sr_reg[8]_140 ;
  output \sr_reg[8]_141 ;
  output \sr_reg[8]_142 ;
  output \sr_reg[8]_143 ;
  output \sr_reg[8]_144 ;
  output \sr_reg[8]_145 ;
  output \sr_reg[1]_4 ;
  output \sr_reg[1]_5 ;
  output \stat_reg[0] ;
  output \sr_reg[5]_1 ;
  output \sr_reg[0]_0 ;
  output [0:0]E;
  output [0:0]\sr_reg[1]_6 ;
  output [0:0]\sr_reg[1]_7 ;
  output [0:0]\sr_reg[1]_8 ;
  output \sr_reg[0]_1 ;
  output \sr_reg[0]_2 ;
  output \sr_reg[0]_3 ;
  output \sr_reg[0]_4 ;
  output \sr_reg[0]_5 ;
  output \sr_reg[0]_6 ;
  output \sr_reg[0]_7 ;
  output \sr_reg[0]_8 ;
  output \sr_reg[0]_9 ;
  output \sr_reg[0]_10 ;
  output \sr_reg[0]_11 ;
  output \sr_reg[0]_12 ;
  output \sr_reg[0]_13 ;
  output \sr_reg[0]_14 ;
  output \sr_reg[0]_15 ;
  output \sr_reg[0]_16 ;
  output \sr_reg[0]_17 ;
  output \sr_reg[0]_18 ;
  output \sr_reg[0]_19 ;
  output \sr_reg[0]_20 ;
  output \sr_reg[0]_21 ;
  output \sr_reg[0]_22 ;
  output \sr_reg[0]_23 ;
  output \sr_reg[0]_24 ;
  output \sr_reg[0]_25 ;
  output \sr_reg[0]_26 ;
  output \sr_reg[0]_27 ;
  output \sr_reg[0]_28 ;
  output \sr_reg[0]_29 ;
  output \sr_reg[0]_30 ;
  output \sr_reg[0]_31 ;
  output \sr_reg[0]_32 ;
  output \sr_reg[0]_33 ;
  output \sr_reg[0]_34 ;
  output \sr_reg[0]_35 ;
  output \sr_reg[0]_36 ;
  output \sr_reg[0]_37 ;
  output \sr_reg[0]_38 ;
  output \sr_reg[0]_39 ;
  output \sr_reg[0]_40 ;
  output \sr_reg[0]_41 ;
  output \sr_reg[0]_42 ;
  output \sr_reg[0]_43 ;
  output \sr_reg[0]_44 ;
  output \sr_reg[0]_45 ;
  output \sr_reg[0]_46 ;
  output \sr_reg[0]_47 ;
  output \sr_reg[0]_48 ;
  output \sr_reg[0]_49 ;
  output \sr_reg[0]_50 ;
  output \sr_reg[0]_51 ;
  output \sr_reg[0]_52 ;
  output \sr_reg[0]_53 ;
  output \sr_reg[0]_54 ;
  output \sr_reg[0]_55 ;
  output \sr_reg[0]_56 ;
  output \sr_reg[0]_57 ;
  output \sr_reg[0]_58 ;
  output \sr_reg[0]_59 ;
  output \sr_reg[0]_60 ;
  output \sr_reg[0]_61 ;
  output \sr_reg[0]_62 ;
  output \sr_reg[0]_63 ;
  output \sr_reg[0]_64 ;
  output \sr_reg[0]_65 ;
  output \sr_reg[0]_66 ;
  output \sr_reg[0]_67 ;
  output \sr_reg[0]_68 ;
  output \sr_reg[0]_69 ;
  output \sr_reg[0]_70 ;
  output \sr_reg[0]_71 ;
  output \sr_reg[0]_72 ;
  output \sr_reg[0]_73 ;
  output \sr_reg[0]_74 ;
  output \sr_reg[0]_75 ;
  output \sr_reg[0]_76 ;
  output \sr_reg[0]_77 ;
  output \sr_reg[0]_78 ;
  output \sr_reg[0]_79 ;
  output \sr_reg[0]_80 ;
  output \sr_reg[0]_81 ;
  output \sr_reg[0]_82 ;
  output \sr_reg[0]_83 ;
  output \sr_reg[0]_84 ;
  output \sr_reg[0]_85 ;
  output \sr_reg[0]_86 ;
  output \sr_reg[0]_87 ;
  output \sr_reg[0]_88 ;
  output \sr_reg[0]_89 ;
  output \sr_reg[0]_90 ;
  output \sr_reg[0]_91 ;
  output \sr_reg[0]_92 ;
  output \sr_reg[0]_93 ;
  output \sr_reg[0]_94 ;
  output \sr_reg[0]_95 ;
  output \sr_reg[0]_96 ;
  output \sr_reg[8]_146 ;
  output \sr_reg[8]_147 ;
  output \sr_reg[8]_148 ;
  output \sr_reg[8]_149 ;
  output \sr_reg[8]_150 ;
  output \sr_reg[8]_151 ;
  output \sr_reg[8]_152 ;
  output \sr_reg[8]_153 ;
  output \sr_reg[8]_154 ;
  output \sr_reg[8]_155 ;
  output \sr_reg[8]_156 ;
  output \sr_reg[8]_157 ;
  output \sr_reg[8]_158 ;
  output \sr_reg[8]_159 ;
  output \sr_reg[8]_160 ;
  output \sr_reg[8]_161 ;
  output \sr_reg[8]_162 ;
  output \sr_reg[8]_163 ;
  output \sr_reg[8]_164 ;
  output \sr_reg[8]_165 ;
  output \sr_reg[8]_166 ;
  output \sr_reg[8]_167 ;
  output \sr_reg[8]_168 ;
  output \sr_reg[8]_169 ;
  output \sr_reg[8]_170 ;
  output \sr_reg[8]_171 ;
  output \sr_reg[8]_172 ;
  output \sr_reg[8]_173 ;
  output \sr_reg[8]_174 ;
  output \sr_reg[8]_175 ;
  output \sr_reg[8]_176 ;
  output \sr_reg[8]_177 ;
  output \sr_reg[8]_178 ;
  output \sr_reg[8]_179 ;
  output \sr_reg[8]_180 ;
  output \sr_reg[8]_181 ;
  output \sr_reg[8]_182 ;
  output \sr_reg[8]_183 ;
  output \sr_reg[8]_184 ;
  output \sr_reg[8]_185 ;
  output \sr_reg[8]_186 ;
  output \sr_reg[8]_187 ;
  output \sr_reg[8]_188 ;
  output \sr_reg[8]_189 ;
  output \sr_reg[8]_190 ;
  output \sr_reg[8]_191 ;
  output \sr_reg[8]_192 ;
  output \sr_reg[8]_193 ;
  output \sr_reg[8]_194 ;
  output \sr_reg[8]_195 ;
  output \sr_reg[8]_196 ;
  output \sr_reg[8]_197 ;
  output \sr_reg[8]_198 ;
  output \sr_reg[8]_199 ;
  output \sr_reg[8]_200 ;
  output \sr_reg[8]_201 ;
  output \sr_reg[8]_202 ;
  output \sr_reg[8]_203 ;
  output \sr_reg[8]_204 ;
  output \sr_reg[8]_205 ;
  output \sr_reg[8]_206 ;
  output \sr_reg[8]_207 ;
  output \sr_reg[8]_208 ;
  output \sr_reg[8]_209 ;
  output \sr_reg[8]_210 ;
  output \sr_reg[8]_211 ;
  output \sr_reg[8]_212 ;
  output \sr_reg[8]_213 ;
  output \sr_reg[8]_214 ;
  output \sr_reg[8]_215 ;
  output \sr_reg[8]_216 ;
  output \sr_reg[8]_217 ;
  output \sr_reg[8]_218 ;
  output [1:0]\sr_reg[8]_219 ;
  output \sr_reg[8]_220 ;
  output \badr[6]_INST_0_i_1 ;
  output \sr_reg[8]_221 ;
  output \badr[4]_INST_0_i_1 ;
  output \sr[6]_i_13 ;
  output \sr_reg[8]_222 ;
  output \sr_reg[8]_223 ;
  output \badr[2]_INST_0_i_1 ;
  output [1:0]niho_dsp_b;
  output \sr_reg[8]_224 ;
  output \sr_reg[8]_225 ;
  output \sr_reg[8]_226 ;
  output \sr_reg[8]_227 ;
  input rst_n;
  input \sr_reg[15]_0 ;
  input [0:0]cbus_sel_0;
  input \sr_reg[5]_2 ;
  input [0:0]\sr_reg[5]_3 ;
  input \sr_reg[6]_4 ;
  input \tr_reg[31] ;
  input \tr_reg[31]_0 ;
  input \sr[4]_i_19 ;
  input \sr[4]_i_19_0 ;
  input \sr[4]_i_19_1 ;
  input \iv[6]_i_3 ;
  input \niho_dsp_b[5] ;
  input \sr[4]_i_38 ;
  input \sr[4]_i_38_0 ;
  input \sr[4]_i_91 ;
  input \tr[23]_i_3 ;
  input \tr[28]_i_3 ;
  input \sr_reg[6]_5 ;
  input \sr[5]_i_3 ;
  input \sr[5]_i_3_0 ;
  input \sr[5]_i_3_1 ;
  input \sr[5]_i_3_2 ;
  input \sr[5]_i_3_3 ;
  input \sr[5]_i_3_4 ;
  input \sr[5]_i_3_5 ;
  input \mul_a_reg[32] ;
  input \sr[4]_i_42_0 ;
  input \sr[4]_i_42_1 ;
  input \sr[4]_i_43 ;
  input \iv[11]_i_4_0 ;
  input \iv[13]_i_4_0 ;
  input \iv[13]_i_4_1 ;
  input \iv[0]_i_3 ;
  input \iv[0]_i_3_0 ;
  input \iv[0]_i_3_1 ;
  input \sr[4]_i_17 ;
  input \sr[4]_i_34 ;
  input \iv[5]_i_3 ;
  input \iv[4]_i_3 ;
  input \sr[4]_i_32 ;
  input \sr[4]_i_39 ;
  input \iv[14]_i_2 ;
  input \sr[4]_i_40 ;
  input \sr[4]_i_37 ;
  input \iv[6]_i_8 ;
  input \iv[9]_i_4 ;
  input \iv[8]_i_4 ;
  input \iv[10]_i_4 ;
  input \iv[3]_i_8 ;
  input \iv[2]_i_8 ;
  input \iv[1]_i_8 ;
  input \iv[7]_i_8 ;
  input \tr[16]_i_2 ;
  input \tr[16]_i_2_0 ;
  input \iv[15]_i_8 ;
  input [2:0]bbus_0;
  input \sr[6]_i_4_0 ;
  input \sr[6]_i_4_1 ;
  input \sr[6]_i_4_2 ;
  input \sr[6]_i_11_0 ;
  input \sr[6]_i_11_1 ;
  input \iv[0]_i_21 ;
  input \iv[15]_i_8_0 ;
  input \iv[15]_i_8_1 ;
  input \iv[15]_i_8_2 ;
  input \sr[4]_i_42_2 ;
  input \sr[4]_i_42_3 ;
  input \sr[4]_i_91_0 ;
  input \iv[10]_i_6 ;
  input \sr[4]_i_74 ;
  input \sr[4]_i_66 ;
  input \tr[27]_i_9 ;
  input \sr[4]_i_73 ;
  input \sr[4]_i_69_0 ;
  input \sr[4]_i_103 ;
  input \sr[4]_i_86 ;
  input \sr[4]_i_94_0 ;
  input \sr[4]_i_87_0 ;
  input \sr[4]_i_90_0 ;
  input \iv[6]_i_10 ;
  input \tr[21]_i_9 ;
  input \iv[9]_i_28 ;
  input \iv[4]_i_27_0 ;
  input \tr[28]_i_8_0 ;
  input \tr[21]_i_8 ;
  input \mul_a_reg[30] ;
  input \tr[26]_i_6 ;
  input \iv[10]_i_29_0 ;
  input \iv[14]_i_13 ;
  input \iv[9]_i_28_0 ;
  input \iv[5]_i_15 ;
  input \iv[15]_i_58 ;
  input \tr[23]_i_6 ;
  input \tr[23]_i_6_0 ;
  input \tr[19]_i_6 ;
  input \iv[8]_i_27 ;
  input \iv[12]_i_25 ;
  input \tr[20]_i_8 ;
  input \tr[24]_i_9 ;
  input \mul_a_reg[29] ;
  input \sr[6]_i_38_0 ;
  input \sr[6]_i_10 ;
  input \sr[4]_i_139_0 ;
  input \mul_a_reg[22] ;
  input \mul_a_reg[21] ;
  input \mul_a_reg[20] ;
  input \mul_a_reg[19] ;
  input \iv[15]_i_96 ;
  input \iv[15]_i_96_0 ;
  input \iv[15]_i_96_1 ;
  input \iv[15]_i_96_2 ;
  input \iv[15]_i_96_3 ;
  input \iv[15]_i_96_4 ;
  input \iv[15]_i_96_5 ;
  input \iv[15]_i_96_6 ;
  input \iv[15]_i_96_7 ;
  input \iv[15]_i_96_8 ;
  input \iv[13]_i_45_0 ;
  input \iv[13]_i_45_1 ;
  input \iv[10]_i_44_1 ;
  input \iv[10]_i_44_2 ;
  input \mul_a_reg[28] ;
  input \mul_a_reg[27] ;
  input \mul_a_reg[26] ;
  input \mul_a_reg[25] ;
  input \mul_a_reg[24] ;
  input \mul_a_reg[23] ;
  input \mul_a_reg[18] ;
  input \mul_a_reg[17] ;
  input \mul_a_reg[16] ;
  input mul_rslt;
  input [15:0]mul_a;
  input \niho_dsp_b[5]_0 ;
  input \remden_reg[26] ;
  input [3:0]DI;
  input \remden_reg[29] ;
  input [3:0]\niho_dsp_a[11] ;
  input \remden_reg[25] ;
  input \remden_reg[24] ;
  input [3:0]\niho_dsp_a[7] ;
  input \remden_reg[23] ;
  input \remden_reg[22] ;
  input \remden_reg[21] ;
  input \iv[5]_i_7 ;
  input \remden_reg[20] ;
  input [3:0]\niho_dsp_a[3] ;
  input \remden_reg[18] ;
  input \remden_reg[17] ;
  input \remden_reg[16] ;
  input \tr[23]_i_5 ;
  input [5:0]Q;
  input \tr[19]_i_2 ;
  input [5:0]\tr[29]_i_2 ;
  input \tr[19]_i_2_0 ;
  input \sr[4]_i_3 ;
  input \sr[4]_i_3_0 ;
  input [0:0]CO;
  input \abus_o[16] ;
  input irq;
  input [1:0]irq_lev;
  input [5:0]\badr[31]_INST_0_i_69 ;
  input \stat_reg[1] ;
  input [1:0]\stat[0]_i_6 ;
  input [0:0]\pc_reg[3]_i_2 ;
  input \sr[4]_i_42_4 ;
  input \sr[4]_i_42_5 ;
  input \sr[4]_i_42_6 ;
  input \sr[4]_i_41 ;
  input \sr[4]_i_41_0 ;
  input \sr[4]_i_47 ;
  input \sr[4]_i_47_0 ;
  input \sr[4]_i_46 ;
  input \sr[4]_i_46_0 ;
  input \sr[4]_i_35 ;
  input \sr[4]_i_35_0 ;
  input \sr[4]_i_33 ;
  input \sr[4]_i_33_0 ;
  input \sr[4]_i_31 ;
  input \sr[4]_i_31_0 ;
  input \sr[4]_i_39_0 ;
  input \sr[4]_i_39_1 ;
  input \sr[4]_i_40_0 ;
  input \sr[4]_i_40_1 ;
  input \sr[4]_i_37_0 ;
  input \sr[4]_i_37_1 ;
  input \grn_reg[0] ;
  input \grn_reg[0]_0 ;
  input [7:0]bbus_sel_0;
  input [15:0]\bdatw[31]_INST_0_i_4 ;
  input [15:0]\bdatw[31]_INST_0_i_4_0 ;
  input [15:0]\i_/badr[31]_INST_0_i_5 ;
  input [15:0]\i_/badr[31]_INST_0_i_5_0 ;
  input [15:0]\bdatw[31]_INST_0_i_4_1 ;
  input [15:0]\bdatw[31]_INST_0_i_4_2 ;
  input [15:0]\i_/badr[31]_INST_0_i_4 ;
  input [15:0]\i_/badr[31]_INST_0_i_4_0 ;
  input [15:0]\i_/badr[31]_INST_0_i_7 ;
  input [15:0]\i_/badr[31]_INST_0_i_7_0 ;
  input [15:0]\i_/badr[31]_INST_0_i_6 ;
  input [15:0]\i_/badr[31]_INST_0_i_6_0 ;
  input [3:0]abus_sel_0;
  input \tr[30]_i_10 ;
  input \tr[21]_i_9_0 ;
  input \tr[21]_i_9_1 ;
  input \tr[26]_i_7 ;
  input \tr[26]_i_7_0 ;
  input \tr[25]_i_9 ;
  input \tr[19]_i_7 ;
  input \tr[28]_i_9 ;
  input \tr[23]_i_7 ;
  input \tr[27]_i_7 ;
  input \tr[18]_i_9 ;
  input \tr[22]_i_9 ;
  input \remden_reg[19] ;
  input \sr[5]_i_2_0 ;
  input \mul_a_reg[32]_0 ;
  input \sr[6]_i_4_3 ;
  input \tr_reg[31]_i_13_0 ;
  input \remden_reg[30] ;
  input \tr_reg[31]_i_13_1 ;
  input \tr_reg[31]_i_13_2 ;
  input \remden_reg[28] ;
  input \tr_reg[31]_i_32_0 ;
  input \remden_reg[27] ;
  input \tr_reg[31]_i_32_1 ;
  input \remden_reg[26]_0 ;
  input \tr_reg[31]_i_32_2 ;
  input \tr_reg[31]_i_32_3 ;
  input \tr_reg[23]_i_11_0 ;
  input \tr_reg[23]_i_11_1 ;
  input \tr_reg[23]_i_11_2 ;
  input \tr_reg[23]_i_11_3 ;
  input \sr_reg[6]_i_6_0 ;
  input \sr_reg[6]_i_6_1 ;
  input \sr_reg[6]_i_6_2 ;
  input \niho_dsp_b[0]_0 ;
  input \niho_dsp_b[5]_1 ;
  input \iv[11]_i_10_0 ;
  input \iv[12]_i_9 ;
  input \tr[20]_i_9 ;
  input clk;
  input [1:0]D;
  input [0:0]SR;
  input \sr_reg[11]_0 ;
  input \sr_reg[10]_0 ;
  input \sr_reg[8]_228 ;
  input \sr_reg[7]_4 ;
  input \sr_reg[6]_6 ;
  input \sr_reg[5]_4 ;
  input \sr_reg[4]_2 ;
  input \sr_reg[3]_0 ;
  input \sr_reg[2]_0 ;
  input \sr_reg[1]_9 ;
  input \sr_reg[0]_97 ;
     output [15:0]sr;
  output irq_lev_0_sn_1;
  output irq_lev_1_sn_1;
  input niho_dsp_b_0_sn_1;
  input niho_dsp_a_15_sn_1;

  wire \<const0> ;
  wire \<const1> ;
  wire [0:0]CO;
  wire [1:0]D;
  wire [3:0]DI;
  wire [0:0]E;
  wire [0:0]O;
  wire [5:0]Q;
  wire [0:0]S;
  wire [0:0]SR;
  wire [15:0]abus_o;
  wire \abus_o[16] ;
  wire [3:0]abus_sel_0;
  wire [34:18]\alu/art/add/tout ;
  wire [16:16]\alu/asr0 ;
  wire [0:0]alu_sr_flag;
  wire \badr[0]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1 ;
  wire \badr[16]_INST_0_i_1_0 ;
  wire \badr[17]_INST_0_i_1 ;
  wire \badr[18]_INST_0_i_1 ;
  wire \badr[1]_INST_0_i_1 ;
  wire \badr[2]_INST_0_i_1 ;
  wire [5:0]\badr[31]_INST_0_i_69 ;
  wire \badr[4]_INST_0_i_1 ;
  wire \badr[5]_INST_0_i_1 ;
  wire \badr[6]_INST_0_i_1 ;
  wire [2:0]bbus_0;
  wire [7:0]bbus_sel_0;
  wire [15:0]\bdatw[31]_INST_0_i_4 ;
  wire [15:0]\bdatw[31]_INST_0_i_4_0 ;
  wire [15:0]\bdatw[31]_INST_0_i_4_1 ;
  wire [15:0]\bdatw[31]_INST_0_i_4_2 ;
  wire [0:0]cbus_sel_0;
  wire clk;
  wire ctl_fetch_inferred_i_43_n_0;
  wire fch_irq_req;
  wire \grn_reg[0] ;
  wire \grn_reg[0]_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_4 ;
  wire [15:0]\i_/badr[31]_INST_0_i_4_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_5 ;
  wire [15:0]\i_/badr[31]_INST_0_i_5_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_6 ;
  wire [15:0]\i_/badr[31]_INST_0_i_6_0 ;
  wire [15:0]\i_/badr[31]_INST_0_i_7 ;
  wire [15:0]\i_/badr[31]_INST_0_i_7_0 ;
  wire irq;
  wire [1:0]irq_lev;
  wire irq_lev_0_sn_1;
  wire irq_lev_1_sn_1;
  wire \iv[0]_i_21 ;
  wire \iv[0]_i_3 ;
  wire \iv[0]_i_31_0 ;
  wire \iv[0]_i_33_n_0 ;
  wire \iv[0]_i_34_n_0 ;
  wire \iv[0]_i_35_n_0 ;
  wire \iv[0]_i_36_n_0 ;
  wire \iv[0]_i_37_n_0 ;
  wire \iv[0]_i_3_0 ;
  wire \iv[0]_i_3_1 ;
  wire \iv[10]_i_23_n_0 ;
  wire \iv[10]_i_29_0 ;
  wire \iv[10]_i_34 ;
  wire \iv[10]_i_4 ;
  wire \iv[10]_i_41_0 ;
  wire \iv[10]_i_41_n_0 ;
  wire \iv[10]_i_44_0 ;
  wire \iv[10]_i_44_1 ;
  wire \iv[10]_i_44_2 ;
  wire \iv[10]_i_44_n_0 ;
  wire \iv[10]_i_6 ;
  wire \iv[10]_i_9 ;
  wire \iv[11]_i_10_0 ;
  wire \iv[11]_i_10_n_0 ;
  wire \iv[11]_i_11_0 ;
  wire \iv[11]_i_11_n_0 ;
  wire \iv[11]_i_23_n_0 ;
  wire \iv[11]_i_24_n_0 ;
  wire \iv[11]_i_42_n_0 ;
  wire \iv[11]_i_47_n_0 ;
  wire \iv[11]_i_4_0 ;
  wire \iv[12]_i_23_n_0 ;
  wire \iv[12]_i_25 ;
  wire \iv[12]_i_38_n_0 ;
  wire \iv[12]_i_39_n_0 ;
  wire \iv[12]_i_40_n_0 ;
  wire \iv[12]_i_41_n_0 ;
  wire \iv[12]_i_42_n_0 ;
  wire \iv[12]_i_43_n_0 ;
  wire \iv[12]_i_47_n_0 ;
  wire \iv[12]_i_48_n_0 ;
  wire \iv[12]_i_49 ;
  wire \iv[12]_i_51_n_0 ;
  wire \iv[12]_i_9 ;
  wire \iv[13]_i_10_0 ;
  wire \iv[13]_i_10_n_0 ;
  wire \iv[13]_i_22_n_0 ;
  wire \iv[13]_i_35 ;
  wire \iv[13]_i_40_n_0 ;
  wire \iv[13]_i_42_n_0 ;
  wire \iv[13]_i_43_n_0 ;
  wire \iv[13]_i_45_0 ;
  wire \iv[13]_i_45_1 ;
  wire \iv[13]_i_48_n_0 ;
  wire \iv[13]_i_49_n_0 ;
  wire \iv[13]_i_4_0 ;
  wire \iv[13]_i_4_1 ;
  wire \iv[13]_i_50 ;
  wire \iv[13]_i_51_n_0 ;
  wire \iv[13]_i_52_n_0 ;
  wire \iv[13]_i_53_n_0 ;
  wire \iv[13]_i_9_n_0 ;
  wire \iv[14]_i_11_0 ;
  wire \iv[14]_i_11_n_0 ;
  wire \iv[14]_i_13 ;
  wire \iv[14]_i_2 ;
  wire \iv[14]_i_27_n_0 ;
  wire \iv[14]_i_30_0 ;
  wire \iv[14]_i_50_n_0 ;
  wire \iv[14]_i_52_n_0 ;
  wire \iv[14]_i_55_n_0 ;
  wire \iv[14]_i_56_n_0 ;
  wire \iv[14]_i_65_n_0 ;
  wire \iv[14]_i_66_n_0 ;
  wire \iv[14]_i_67_n_0 ;
  wire \iv[14]_i_68_n_0 ;
  wire \iv[14]_i_69_n_0 ;
  wire \iv[14]_i_70_n_0 ;
  wire \iv[15]_i_108 ;
  wire \iv[15]_i_108_0 ;
  wire \iv[15]_i_108_1 ;
  wire \iv[15]_i_108_10 ;
  wire \iv[15]_i_108_11 ;
  wire \iv[15]_i_108_12 ;
  wire \iv[15]_i_108_13 ;
  wire \iv[15]_i_108_2 ;
  wire \iv[15]_i_108_3 ;
  wire \iv[15]_i_108_4 ;
  wire \iv[15]_i_108_5 ;
  wire \iv[15]_i_108_6 ;
  wire \iv[15]_i_108_7 ;
  wire \iv[15]_i_108_8 ;
  wire \iv[15]_i_108_9 ;
  wire \iv[15]_i_127_n_0 ;
  wire \iv[15]_i_128_n_0 ;
  wire \iv[15]_i_131_n_0 ;
  wire \iv[15]_i_132_n_0 ;
  wire \iv[15]_i_133_n_0 ;
  wire \iv[15]_i_134_n_0 ;
  wire \iv[15]_i_136_n_0 ;
  wire \iv[15]_i_138_n_0 ;
  wire \iv[15]_i_141_n_0 ;
  wire \iv[15]_i_142_n_0 ;
  wire \iv[15]_i_143_n_0 ;
  wire \iv[15]_i_144_n_0 ;
  wire \iv[15]_i_145_n_0 ;
  wire \iv[15]_i_146_n_0 ;
  wire \iv[15]_i_147_n_0 ;
  wire \iv[15]_i_163_n_0 ;
  wire \iv[15]_i_164_n_0 ;
  wire \iv[15]_i_165_n_0 ;
  wire \iv[15]_i_166_n_0 ;
  wire \iv[15]_i_168_n_0 ;
  wire \iv[15]_i_169_n_0 ;
  wire \iv[15]_i_170_n_0 ;
  wire \iv[15]_i_51_n_0 ;
  wire \iv[15]_i_54_n_0 ;
  wire \iv[15]_i_58 ;
  wire \iv[15]_i_62_n_0 ;
  wire \iv[15]_i_8 ;
  wire \iv[15]_i_8_0 ;
  wire \iv[15]_i_8_1 ;
  wire \iv[15]_i_8_2 ;
  wire \iv[15]_i_95_n_0 ;
  wire \iv[15]_i_96 ;
  wire \iv[15]_i_96_0 ;
  wire \iv[15]_i_96_1 ;
  wire \iv[15]_i_96_2 ;
  wire \iv[15]_i_96_3 ;
  wire \iv[15]_i_96_4 ;
  wire \iv[15]_i_96_5 ;
  wire \iv[15]_i_96_6 ;
  wire \iv[15]_i_96_7 ;
  wire \iv[15]_i_96_8 ;
  wire \iv[1]_i_8 ;
  wire \iv[2]_i_8 ;
  wire \iv[3]_i_41_0 ;
  wire \iv[3]_i_41_n_0 ;
  wire \iv[3]_i_42_n_0 ;
  wire \iv[3]_i_8 ;
  wire \iv[4]_i_27_0 ;
  wire \iv[4]_i_3 ;
  wire \iv[4]_i_35_0 ;
  wire \iv[4]_i_35_n_0 ;
  wire \iv[4]_i_36_n_0 ;
  wire \iv[5]_i_15 ;
  wire \iv[5]_i_3 ;
  wire \iv[5]_i_7 ;
  wire \iv[6]_i_10 ;
  wire \iv[6]_i_28_n_0 ;
  wire \iv[6]_i_3 ;
  wire \iv[6]_i_8 ;
  wire \iv[7]_i_36_n_0 ;
  wire \iv[7]_i_47_n_0 ;
  wire \iv[7]_i_48_n_0 ;
  wire \iv[7]_i_8 ;
  wire \iv[8]_i_27 ;
  wire \iv[8]_i_34 ;
  wire \iv[8]_i_38 ;
  wire \iv[8]_i_4 ;
  wire \iv[9]_i_28 ;
  wire \iv[9]_i_28_0 ;
  wire \iv[9]_i_4 ;
  wire \iv[9]_i_46_0 ;
  wire \iv[9]_i_46_n_0 ;
  wire [15:0]mul_a;
  wire [13:0]mul_a_i;
  wire \mul_a_reg[16] ;
  wire \mul_a_reg[17] ;
  wire \mul_a_reg[18] ;
  wire \mul_a_reg[19] ;
  wire \mul_a_reg[20] ;
  wire \mul_a_reg[21] ;
  wire \mul_a_reg[22] ;
  wire \mul_a_reg[23] ;
  wire \mul_a_reg[24] ;
  wire \mul_a_reg[25] ;
  wire \mul_a_reg[26] ;
  wire \mul_a_reg[27] ;
  wire \mul_a_reg[28] ;
  wire \mul_a_reg[29] ;
  wire \mul_a_reg[30] ;
  wire \mul_a_reg[32] ;
  wire \mul_a_reg[32]_0 ;
  wire mul_rslt;
  wire mul_rslt0;
  wire [15:0]niho_dsp_a;
  wire [3:0]\niho_dsp_a[11] ;
  wire [3:0]\niho_dsp_a[3] ;
  wire [3:0]\niho_dsp_a[7] ;
  wire niho_dsp_a_15_sn_1;
  wire [1:0]niho_dsp_b;
  wire \niho_dsp_b[0]_0 ;
  wire \niho_dsp_b[5] ;
  wire \niho_dsp_b[5]_0 ;
  wire \niho_dsp_b[5]_1 ;
  wire niho_dsp_b_0_sn_1;
  wire [15:9]p_0_in__0;
  wire [0:0]p_2_in;
  wire [0:0]\pc_reg[3]_i_2 ;
  wire \quo_reg[19] ;
  wire \quo_reg[23] ;
  wire \quo_reg[27] ;
  wire \rem_reg[21] ;
  wire \rem_reg[28] ;
  wire \rem_reg[29] ;
  wire \remden_reg[16] ;
  wire \remden_reg[17] ;
  wire \remden_reg[18] ;
  wire \remden_reg[19] ;
  wire \remden_reg[20] ;
  wire \remden_reg[21] ;
  wire \remden_reg[22] ;
  wire \remden_reg[23] ;
  wire \remden_reg[24] ;
  wire \remden_reg[25] ;
  wire \remden_reg[26] ;
  wire \remden_reg[26]_0 ;
  wire \remden_reg[27] ;
  wire \remden_reg[28] ;
  wire \remden_reg[29] ;
  wire \remden_reg[30] ;
  wire rst_n;
  (* DONT_TOUCH *) wire [15:0]sr;
  wire \sr[4]_i_103 ;
  wire \sr[4]_i_111_n_0 ;
  wire \sr[4]_i_112_n_0 ;
  wire \sr[4]_i_119_n_0 ;
  wire \sr[4]_i_121_n_0 ;
  wire \sr[4]_i_128_n_0 ;
  wire \sr[4]_i_130_n_0 ;
  wire \sr[4]_i_139_0 ;
  wire \sr[4]_i_141_n_0 ;
  wire \sr[4]_i_143_n_0 ;
  wire \sr[4]_i_145_n_0 ;
  wire \sr[4]_i_150_n_0 ;
  wire \sr[4]_i_152_n_0 ;
  wire \sr[4]_i_163_n_0 ;
  wire \sr[4]_i_164_n_0 ;
  wire \sr[4]_i_169_n_0 ;
  wire \sr[4]_i_17 ;
  wire \sr[4]_i_170_n_0 ;
  wire \sr[4]_i_19 ;
  wire \sr[4]_i_19_0 ;
  wire \sr[4]_i_19_1 ;
  wire \sr[4]_i_28_n_0 ;
  wire \sr[4]_i_3 ;
  wire \sr[4]_i_31 ;
  wire \sr[4]_i_31_0 ;
  wire \sr[4]_i_32 ;
  wire \sr[4]_i_33 ;
  wire \sr[4]_i_33_0 ;
  wire \sr[4]_i_34 ;
  wire \sr[4]_i_35 ;
  wire \sr[4]_i_35_0 ;
  wire \sr[4]_i_37 ;
  wire \sr[4]_i_37_0 ;
  wire \sr[4]_i_37_1 ;
  wire \sr[4]_i_38 ;
  wire \sr[4]_i_38_0 ;
  wire \sr[4]_i_39 ;
  wire \sr[4]_i_39_0 ;
  wire \sr[4]_i_39_1 ;
  wire \sr[4]_i_3_0 ;
  wire \sr[4]_i_40 ;
  wire \sr[4]_i_40_0 ;
  wire \sr[4]_i_40_1 ;
  wire \sr[4]_i_41 ;
  wire \sr[4]_i_41_0 ;
  wire \sr[4]_i_42_0 ;
  wire \sr[4]_i_42_1 ;
  wire \sr[4]_i_42_2 ;
  wire \sr[4]_i_42_3 ;
  wire \sr[4]_i_42_4 ;
  wire \sr[4]_i_42_5 ;
  wire \sr[4]_i_42_6 ;
  wire \sr[4]_i_43 ;
  wire \sr[4]_i_46 ;
  wire \sr[4]_i_46_0 ;
  wire \sr[4]_i_47 ;
  wire \sr[4]_i_47_0 ;
  wire \sr[4]_i_48_n_0 ;
  wire \sr[4]_i_49_n_0 ;
  wire \sr[4]_i_66 ;
  wire \sr[4]_i_69_0 ;
  wire \sr[4]_i_73 ;
  wire \sr[4]_i_74 ;
  wire \sr[4]_i_86 ;
  wire \sr[4]_i_87_0 ;
  wire \sr[4]_i_87_n_0 ;
  wire \sr[4]_i_88_n_0 ;
  wire \sr[4]_i_90_0 ;
  wire \sr[4]_i_90_n_0 ;
  wire \sr[4]_i_91 ;
  wire \sr[4]_i_91_0 ;
  wire \sr[4]_i_94_0 ;
  wire \sr[5]_i_2_0 ;
  wire \sr[5]_i_3 ;
  wire \sr[5]_i_3_0 ;
  wire \sr[5]_i_3_1 ;
  wire \sr[5]_i_3_2 ;
  wire \sr[5]_i_3_3 ;
  wire \sr[5]_i_3_4 ;
  wire \sr[5]_i_3_5 ;
  wire \sr[5]_i_7_n_0 ;
  wire \sr[6]_i_10 ;
  wire \sr[6]_i_11_0 ;
  wire \sr[6]_i_11_1 ;
  wire \sr[6]_i_11_n_0 ;
  wire \sr[6]_i_13 ;
  wire \sr[6]_i_15_n_0 ;
  wire \sr[6]_i_16_n_0 ;
  wire \sr[6]_i_17_n_0 ;
  wire \sr[6]_i_18_n_0 ;
  wire \sr[6]_i_19_n_0 ;
  wire \sr[6]_i_20_n_0 ;
  wire \sr[6]_i_21_n_0 ;
  wire \sr[6]_i_22_n_0 ;
  wire \sr[6]_i_23_n_0 ;
  wire \sr[6]_i_24_n_0 ;
  wire \sr[6]_i_29_n_0 ;
  wire \sr[6]_i_33_n_0 ;
  wire \sr[6]_i_38_0 ;
  wire \sr[6]_i_41_n_0 ;
  wire \sr[6]_i_4_0 ;
  wire \sr[6]_i_4_1 ;
  wire \sr[6]_i_4_2 ;
  wire \sr[6]_i_4_3 ;
  wire \sr[6]_i_9_n_0 ;
  wire \sr[7]_i_26_n_0 ;
  wire \sr[7]_i_30_n_0 ;
  wire \sr[7]_i_45_n_0 ;
  wire \sr[7]_i_46_n_0 ;
  wire \sr[7]_i_47_n_0 ;
  wire \sr[7]_i_48_n_0 ;
  wire \sr[7]_i_50_n_0 ;
  wire \sr[7]_i_51_n_0 ;
  wire \sr[7]_i_52_n_0 ;
  wire \sr[7]_i_9_n_0 ;
  wire \sr_reg[0]_0 ;
  wire \sr_reg[0]_1 ;
  wire \sr_reg[0]_10 ;
  wire \sr_reg[0]_11 ;
  wire \sr_reg[0]_12 ;
  wire \sr_reg[0]_13 ;
  wire \sr_reg[0]_14 ;
  wire \sr_reg[0]_15 ;
  wire \sr_reg[0]_16 ;
  wire \sr_reg[0]_17 ;
  wire \sr_reg[0]_18 ;
  wire \sr_reg[0]_19 ;
  wire \sr_reg[0]_2 ;
  wire \sr_reg[0]_20 ;
  wire \sr_reg[0]_21 ;
  wire \sr_reg[0]_22 ;
  wire \sr_reg[0]_23 ;
  wire \sr_reg[0]_24 ;
  wire \sr_reg[0]_25 ;
  wire \sr_reg[0]_26 ;
  wire \sr_reg[0]_27 ;
  wire \sr_reg[0]_28 ;
  wire \sr_reg[0]_29 ;
  wire \sr_reg[0]_3 ;
  wire \sr_reg[0]_30 ;
  wire \sr_reg[0]_31 ;
  wire \sr_reg[0]_32 ;
  wire \sr_reg[0]_33 ;
  wire \sr_reg[0]_34 ;
  wire \sr_reg[0]_35 ;
  wire \sr_reg[0]_36 ;
  wire \sr_reg[0]_37 ;
  wire \sr_reg[0]_38 ;
  wire \sr_reg[0]_39 ;
  wire \sr_reg[0]_4 ;
  wire \sr_reg[0]_40 ;
  wire \sr_reg[0]_41 ;
  wire \sr_reg[0]_42 ;
  wire \sr_reg[0]_43 ;
  wire \sr_reg[0]_44 ;
  wire \sr_reg[0]_45 ;
  wire \sr_reg[0]_46 ;
  wire \sr_reg[0]_47 ;
  wire \sr_reg[0]_48 ;
  wire \sr_reg[0]_49 ;
  wire \sr_reg[0]_5 ;
  wire \sr_reg[0]_50 ;
  wire \sr_reg[0]_51 ;
  wire \sr_reg[0]_52 ;
  wire \sr_reg[0]_53 ;
  wire \sr_reg[0]_54 ;
  wire \sr_reg[0]_55 ;
  wire \sr_reg[0]_56 ;
  wire \sr_reg[0]_57 ;
  wire \sr_reg[0]_58 ;
  wire \sr_reg[0]_59 ;
  wire \sr_reg[0]_6 ;
  wire \sr_reg[0]_60 ;
  wire \sr_reg[0]_61 ;
  wire \sr_reg[0]_62 ;
  wire \sr_reg[0]_63 ;
  wire \sr_reg[0]_64 ;
  wire \sr_reg[0]_65 ;
  wire \sr_reg[0]_66 ;
  wire \sr_reg[0]_67 ;
  wire \sr_reg[0]_68 ;
  wire \sr_reg[0]_69 ;
  wire \sr_reg[0]_7 ;
  wire \sr_reg[0]_70 ;
  wire \sr_reg[0]_71 ;
  wire \sr_reg[0]_72 ;
  wire \sr_reg[0]_73 ;
  wire \sr_reg[0]_74 ;
  wire \sr_reg[0]_75 ;
  wire \sr_reg[0]_76 ;
  wire \sr_reg[0]_77 ;
  wire \sr_reg[0]_78 ;
  wire \sr_reg[0]_79 ;
  wire \sr_reg[0]_8 ;
  wire \sr_reg[0]_80 ;
  wire \sr_reg[0]_81 ;
  wire \sr_reg[0]_82 ;
  wire \sr_reg[0]_83 ;
  wire \sr_reg[0]_84 ;
  wire \sr_reg[0]_85 ;
  wire \sr_reg[0]_86 ;
  wire \sr_reg[0]_87 ;
  wire \sr_reg[0]_88 ;
  wire \sr_reg[0]_89 ;
  wire \sr_reg[0]_9 ;
  wire \sr_reg[0]_90 ;
  wire \sr_reg[0]_91 ;
  wire \sr_reg[0]_92 ;
  wire \sr_reg[0]_93 ;
  wire \sr_reg[0]_94 ;
  wire \sr_reg[0]_95 ;
  wire \sr_reg[0]_96 ;
  wire \sr_reg[0]_97 ;
  wire \sr_reg[10]_0 ;
  wire \sr_reg[11]_0 ;
  wire \sr_reg[15]_0 ;
  wire [0:0]\sr_reg[1]_0 ;
  wire [0:0]\sr_reg[1]_1 ;
  wire [0:0]\sr_reg[1]_2 ;
  wire [0:0]\sr_reg[1]_3 ;
  wire \sr_reg[1]_4 ;
  wire \sr_reg[1]_5 ;
  wire [0:0]\sr_reg[1]_6 ;
  wire [0:0]\sr_reg[1]_7 ;
  wire [0:0]\sr_reg[1]_8 ;
  wire \sr_reg[1]_9 ;
  wire \sr_reg[2]_0 ;
  wire \sr_reg[3]_0 ;
  wire \sr_reg[4]_0 ;
  wire \sr_reg[4]_1 ;
  wire \sr_reg[4]_2 ;
  wire \sr_reg[5]_0 ;
  wire \sr_reg[5]_1 ;
  wire \sr_reg[5]_2 ;
  wire [0:0]\sr_reg[5]_3 ;
  wire \sr_reg[5]_4 ;
  wire \sr_reg[6]_0 ;
  wire \sr_reg[6]_1 ;
  wire \sr_reg[6]_2 ;
  wire \sr_reg[6]_3 ;
  wire \sr_reg[6]_4 ;
  wire \sr_reg[6]_5 ;
  wire \sr_reg[6]_6 ;
  wire \sr_reg[6]_i_6_0 ;
  wire \sr_reg[6]_i_6_1 ;
  wire \sr_reg[6]_i_6_2 ;
  wire \sr_reg[6]_i_6_n_0 ;
  wire \sr_reg[6]_i_6_n_1 ;
  wire \sr_reg[6]_i_6_n_2 ;
  wire \sr_reg[6]_i_6_n_3 ;
  wire \sr_reg[6]_i_6_n_4 ;
  wire \sr_reg[6]_i_6_n_5 ;
  wire \sr_reg[6]_i_6_n_7 ;
  wire \sr_reg[7]_0 ;
  wire \sr_reg[7]_1 ;
  wire \sr_reg[7]_2 ;
  wire \sr_reg[7]_3 ;
  wire \sr_reg[7]_4 ;
  wire \sr_reg[8]_0 ;
  wire \sr_reg[8]_1 ;
  wire \sr_reg[8]_10 ;
  wire \sr_reg[8]_100 ;
  wire \sr_reg[8]_101 ;
  wire \sr_reg[8]_102 ;
  wire \sr_reg[8]_103 ;
  wire \sr_reg[8]_104 ;
  wire \sr_reg[8]_105 ;
  wire \sr_reg[8]_106 ;
  wire \sr_reg[8]_107 ;
  wire \sr_reg[8]_108 ;
  wire \sr_reg[8]_109 ;
  wire \sr_reg[8]_11 ;
  wire \sr_reg[8]_110 ;
  wire \sr_reg[8]_111 ;
  wire \sr_reg[8]_112 ;
  wire \sr_reg[8]_113 ;
  wire \sr_reg[8]_114 ;
  wire \sr_reg[8]_115 ;
  wire \sr_reg[8]_116 ;
  wire \sr_reg[8]_117 ;
  wire \sr_reg[8]_118 ;
  wire \sr_reg[8]_119 ;
  wire \sr_reg[8]_12 ;
  wire \sr_reg[8]_120 ;
  wire \sr_reg[8]_121 ;
  wire \sr_reg[8]_122 ;
  wire \sr_reg[8]_123 ;
  wire \sr_reg[8]_124 ;
  wire \sr_reg[8]_125 ;
  wire \sr_reg[8]_126 ;
  wire \sr_reg[8]_127 ;
  wire \sr_reg[8]_128 ;
  wire \sr_reg[8]_129 ;
  wire \sr_reg[8]_13 ;
  wire \sr_reg[8]_130 ;
  wire \sr_reg[8]_131 ;
  wire \sr_reg[8]_132 ;
  wire \sr_reg[8]_133 ;
  wire \sr_reg[8]_134 ;
  wire \sr_reg[8]_135 ;
  wire \sr_reg[8]_136 ;
  wire \sr_reg[8]_137 ;
  wire \sr_reg[8]_138 ;
  wire \sr_reg[8]_139 ;
  wire \sr_reg[8]_14 ;
  wire \sr_reg[8]_140 ;
  wire \sr_reg[8]_141 ;
  wire \sr_reg[8]_142 ;
  wire \sr_reg[8]_143 ;
  wire \sr_reg[8]_144 ;
  wire \sr_reg[8]_145 ;
  wire \sr_reg[8]_146 ;
  wire \sr_reg[8]_147 ;
  wire \sr_reg[8]_148 ;
  wire \sr_reg[8]_149 ;
  wire \sr_reg[8]_15 ;
  wire \sr_reg[8]_150 ;
  wire \sr_reg[8]_151 ;
  wire \sr_reg[8]_152 ;
  wire \sr_reg[8]_153 ;
  wire \sr_reg[8]_154 ;
  wire \sr_reg[8]_155 ;
  wire \sr_reg[8]_156 ;
  wire \sr_reg[8]_157 ;
  wire \sr_reg[8]_158 ;
  wire \sr_reg[8]_159 ;
  wire \sr_reg[8]_16 ;
  wire \sr_reg[8]_160 ;
  wire \sr_reg[8]_161 ;
  wire \sr_reg[8]_162 ;
  wire \sr_reg[8]_163 ;
  wire \sr_reg[8]_164 ;
  wire \sr_reg[8]_165 ;
  wire \sr_reg[8]_166 ;
  wire \sr_reg[8]_167 ;
  wire \sr_reg[8]_168 ;
  wire \sr_reg[8]_169 ;
  wire \sr_reg[8]_17 ;
  wire \sr_reg[8]_170 ;
  wire \sr_reg[8]_171 ;
  wire \sr_reg[8]_172 ;
  wire \sr_reg[8]_173 ;
  wire \sr_reg[8]_174 ;
  wire \sr_reg[8]_175 ;
  wire \sr_reg[8]_176 ;
  wire \sr_reg[8]_177 ;
  wire \sr_reg[8]_178 ;
  wire \sr_reg[8]_179 ;
  wire \sr_reg[8]_18 ;
  wire \sr_reg[8]_180 ;
  wire \sr_reg[8]_181 ;
  wire \sr_reg[8]_182 ;
  wire \sr_reg[8]_183 ;
  wire \sr_reg[8]_184 ;
  wire \sr_reg[8]_185 ;
  wire \sr_reg[8]_186 ;
  wire \sr_reg[8]_187 ;
  wire \sr_reg[8]_188 ;
  wire \sr_reg[8]_189 ;
  wire \sr_reg[8]_19 ;
  wire \sr_reg[8]_190 ;
  wire \sr_reg[8]_191 ;
  wire \sr_reg[8]_192 ;
  wire \sr_reg[8]_193 ;
  wire \sr_reg[8]_194 ;
  wire \sr_reg[8]_195 ;
  wire \sr_reg[8]_196 ;
  wire \sr_reg[8]_197 ;
  wire \sr_reg[8]_198 ;
  wire \sr_reg[8]_199 ;
  wire \sr_reg[8]_2 ;
  wire \sr_reg[8]_20 ;
  wire \sr_reg[8]_200 ;
  wire \sr_reg[8]_201 ;
  wire \sr_reg[8]_202 ;
  wire \sr_reg[8]_203 ;
  wire \sr_reg[8]_204 ;
  wire \sr_reg[8]_205 ;
  wire \sr_reg[8]_206 ;
  wire \sr_reg[8]_207 ;
  wire \sr_reg[8]_208 ;
  wire \sr_reg[8]_209 ;
  wire \sr_reg[8]_21 ;
  wire \sr_reg[8]_210 ;
  wire \sr_reg[8]_211 ;
  wire \sr_reg[8]_212 ;
  wire \sr_reg[8]_213 ;
  wire \sr_reg[8]_214 ;
  wire \sr_reg[8]_215 ;
  wire \sr_reg[8]_216 ;
  wire \sr_reg[8]_217 ;
  wire \sr_reg[8]_218 ;
  wire [1:0]\sr_reg[8]_219 ;
  wire \sr_reg[8]_22 ;
  wire \sr_reg[8]_220 ;
  wire \sr_reg[8]_221 ;
  wire \sr_reg[8]_222 ;
  wire \sr_reg[8]_223 ;
  wire \sr_reg[8]_224 ;
  wire \sr_reg[8]_225 ;
  wire \sr_reg[8]_226 ;
  wire \sr_reg[8]_227 ;
  wire \sr_reg[8]_228 ;
  wire \sr_reg[8]_23 ;
  wire \sr_reg[8]_24 ;
  wire \sr_reg[8]_25 ;
  wire \sr_reg[8]_26 ;
  wire \sr_reg[8]_27 ;
  wire \sr_reg[8]_28 ;
  wire \sr_reg[8]_29 ;
  wire \sr_reg[8]_3 ;
  wire \sr_reg[8]_30 ;
  wire \sr_reg[8]_31 ;
  wire \sr_reg[8]_32 ;
  wire \sr_reg[8]_33 ;
  wire \sr_reg[8]_34 ;
  wire \sr_reg[8]_35 ;
  wire \sr_reg[8]_36 ;
  wire \sr_reg[8]_37 ;
  wire \sr_reg[8]_38 ;
  wire \sr_reg[8]_39 ;
  wire \sr_reg[8]_4 ;
  wire \sr_reg[8]_40 ;
  wire \sr_reg[8]_41 ;
  wire \sr_reg[8]_42 ;
  wire \sr_reg[8]_43 ;
  wire \sr_reg[8]_44 ;
  wire \sr_reg[8]_45 ;
  wire \sr_reg[8]_46 ;
  wire \sr_reg[8]_47 ;
  wire \sr_reg[8]_48 ;
  wire \sr_reg[8]_49 ;
  wire \sr_reg[8]_5 ;
  wire \sr_reg[8]_50 ;
  wire \sr_reg[8]_51 ;
  wire \sr_reg[8]_52 ;
  wire \sr_reg[8]_53 ;
  wire \sr_reg[8]_54 ;
  wire \sr_reg[8]_55 ;
  wire \sr_reg[8]_56 ;
  wire \sr_reg[8]_57 ;
  wire \sr_reg[8]_58 ;
  wire \sr_reg[8]_59 ;
  wire \sr_reg[8]_6 ;
  wire \sr_reg[8]_60 ;
  wire \sr_reg[8]_61 ;
  wire \sr_reg[8]_62 ;
  wire \sr_reg[8]_63 ;
  wire \sr_reg[8]_64 ;
  wire \sr_reg[8]_65 ;
  wire \sr_reg[8]_66 ;
  wire \sr_reg[8]_67 ;
  wire \sr_reg[8]_68 ;
  wire \sr_reg[8]_69 ;
  wire \sr_reg[8]_7 ;
  wire \sr_reg[8]_70 ;
  wire \sr_reg[8]_71 ;
  wire \sr_reg[8]_72 ;
  wire \sr_reg[8]_73 ;
  wire \sr_reg[8]_74 ;
  wire \sr_reg[8]_75 ;
  wire \sr_reg[8]_76 ;
  wire \sr_reg[8]_77 ;
  wire \sr_reg[8]_78 ;
  wire \sr_reg[8]_79 ;
  wire \sr_reg[8]_8 ;
  wire \sr_reg[8]_80 ;
  wire \sr_reg[8]_81 ;
  wire \sr_reg[8]_82 ;
  wire \sr_reg[8]_83 ;
  wire \sr_reg[8]_84 ;
  wire \sr_reg[8]_85 ;
  wire \sr_reg[8]_86 ;
  wire \sr_reg[8]_87 ;
  wire \sr_reg[8]_88 ;
  wire \sr_reg[8]_89 ;
  wire \sr_reg[8]_9 ;
  wire \sr_reg[8]_90 ;
  wire \sr_reg[8]_91 ;
  wire \sr_reg[8]_92 ;
  wire \sr_reg[8]_93 ;
  wire \sr_reg[8]_94 ;
  wire \sr_reg[8]_95 ;
  wire \sr_reg[8]_96 ;
  wire \sr_reg[8]_97 ;
  wire \sr_reg[8]_98 ;
  wire \sr_reg[8]_99 ;
  wire [1:0]\stat[0]_i_6 ;
  wire \stat[2]_i_10_n_0 ;
  wire \stat_reg[0] ;
  wire \stat_reg[1] ;
  wire \tr[16]_i_11_n_0 ;
  wire \tr[16]_i_2 ;
  wire \tr[16]_i_25_n_0 ;
  wire \tr[16]_i_2_0 ;
  wire \tr[18]_i_9 ;
  wire \tr[19]_i_2 ;
  wire \tr[19]_i_2_0 ;
  wire \tr[19]_i_6 ;
  wire \tr[19]_i_7 ;
  wire \tr[20]_i_8 ;
  wire \tr[20]_i_9 ;
  wire \tr[21]_i_8 ;
  wire \tr[21]_i_9 ;
  wire \tr[21]_i_9_0 ;
  wire \tr[21]_i_9_1 ;
  wire \tr[22]_i_9 ;
  wire \tr[23]_i_16_n_0 ;
  wire \tr[23]_i_17_n_0 ;
  wire \tr[23]_i_18_n_0 ;
  wire \tr[23]_i_19_n_0 ;
  wire \tr[23]_i_20_n_0 ;
  wire \tr[23]_i_21_n_0 ;
  wire \tr[23]_i_22_n_0 ;
  wire \tr[23]_i_23_n_0 ;
  wire \tr[23]_i_3 ;
  wire \tr[23]_i_5 ;
  wire \tr[23]_i_6 ;
  wire \tr[23]_i_6_0 ;
  wire \tr[23]_i_7 ;
  wire \tr[24]_i_9 ;
  wire \tr[25]_i_9 ;
  wire \tr[26]_i_6 ;
  wire \tr[26]_i_7 ;
  wire \tr[26]_i_7_0 ;
  wire \tr[27]_i_18_n_0 ;
  wire \tr[27]_i_7 ;
  wire \tr[27]_i_9 ;
  wire \tr[28]_i_3 ;
  wire \tr[28]_i_8_0 ;
  wire \tr[28]_i_9 ;
  wire \tr[29]_i_10_n_0 ;
  wire [5:0]\tr[29]_i_2 ;
  wire \tr[30]_i_10 ;
  wire \tr[31]_i_33_n_0 ;
  wire \tr[31]_i_34_n_0 ;
  wire \tr[31]_i_35_n_0 ;
  wire \tr[31]_i_36_n_0 ;
  wire \tr[31]_i_37_n_0 ;
  wire \tr[31]_i_38_n_0 ;
  wire \tr[31]_i_39_n_0 ;
  wire \tr[31]_i_40_n_0 ;
  wire \tr[31]_i_62_n_0 ;
  wire \tr[31]_i_63_n_0 ;
  wire \tr[31]_i_64_n_0 ;
  wire \tr[31]_i_65_n_0 ;
  wire \tr[31]_i_66_n_0 ;
  wire \tr[31]_i_67_n_0 ;
  wire \tr[31]_i_68_n_0 ;
  wire \tr[31]_i_69_n_0 ;
  wire \tr_reg[23]_i_11_0 ;
  wire \tr_reg[23]_i_11_1 ;
  wire \tr_reg[23]_i_11_2 ;
  wire \tr_reg[23]_i_11_3 ;
  wire \tr_reg[23]_i_11_n_0 ;
  wire \tr_reg[23]_i_11_n_1 ;
  wire \tr_reg[23]_i_11_n_2 ;
  wire \tr_reg[23]_i_11_n_3 ;
  wire \tr_reg[23]_i_11_n_4 ;
  wire \tr_reg[23]_i_11_n_5 ;
  wire \tr_reg[23]_i_11_n_6 ;
  wire \tr_reg[23]_i_11_n_7 ;
  wire \tr_reg[31] ;
  wire \tr_reg[31]_0 ;
  wire \tr_reg[31]_i_13_0 ;
  wire \tr_reg[31]_i_13_1 ;
  wire \tr_reg[31]_i_13_2 ;
  wire \tr_reg[31]_i_13_n_0 ;
  wire \tr_reg[31]_i_13_n_1 ;
  wire \tr_reg[31]_i_13_n_2 ;
  wire \tr_reg[31]_i_13_n_3 ;
  wire \tr_reg[31]_i_13_n_5 ;
  wire \tr_reg[31]_i_13_n_6 ;
  wire \tr_reg[31]_i_13_n_7 ;
  wire \tr_reg[31]_i_32_0 ;
  wire \tr_reg[31]_i_32_1 ;
  wire \tr_reg[31]_i_32_2 ;
  wire \tr_reg[31]_i_32_3 ;
  wire \tr_reg[31]_i_32_n_0 ;
  wire \tr_reg[31]_i_32_n_1 ;
  wire \tr_reg[31]_i_32_n_2 ;
  wire \tr_reg[31]_i_32_n_3 ;
  wire \tr_reg[31]_i_32_n_4 ;
  wire \tr_reg[31]_i_32_n_5 ;
  wire \tr_reg[31]_i_32_n_6 ;
  wire \tr_reg[31]_i_32_n_7 ;

  GND GND
       (.G(\<const0> ));
  VCC VCC
       (.P(\<const1> ));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[16]_INST_0 
       (.I0(\mul_a_reg[16] ),
        .I1(\abus_o[16] ),
        .O(abus_o[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[17]_INST_0 
       (.I0(\mul_a_reg[17] ),
        .I1(\abus_o[16] ),
        .O(abus_o[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[18]_INST_0 
       (.I0(\mul_a_reg[18] ),
        .I1(\abus_o[16] ),
        .O(abus_o[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[19]_INST_0 
       (.I0(\mul_a_reg[19] ),
        .I1(\abus_o[16] ),
        .O(abus_o[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[20]_INST_0 
       (.I0(\mul_a_reg[20] ),
        .I1(\abus_o[16] ),
        .O(abus_o[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[21]_INST_0 
       (.I0(\mul_a_reg[21] ),
        .I1(\abus_o[16] ),
        .O(abus_o[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[22]_INST_0 
       (.I0(\mul_a_reg[22] ),
        .I1(\abus_o[16] ),
        .O(abus_o[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[23]_INST_0 
       (.I0(\mul_a_reg[23] ),
        .I1(\abus_o[16] ),
        .O(abus_o[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[24]_INST_0 
       (.I0(\mul_a_reg[24] ),
        .I1(\abus_o[16] ),
        .O(abus_o[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[25]_INST_0 
       (.I0(\mul_a_reg[25] ),
        .I1(\abus_o[16] ),
        .O(abus_o[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[26]_INST_0 
       (.I0(\mul_a_reg[26] ),
        .I1(\abus_o[16] ),
        .O(abus_o[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[27]_INST_0 
       (.I0(\mul_a_reg[27] ),
        .I1(\abus_o[16] ),
        .O(abus_o[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[28]_INST_0 
       (.I0(\mul_a_reg[28] ),
        .I1(\abus_o[16] ),
        .O(abus_o[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[29]_INST_0 
       (.I0(\mul_a_reg[29] ),
        .I1(\abus_o[16] ),
        .O(abus_o[13]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[30]_INST_0 
       (.I0(\mul_a_reg[30] ),
        .I1(\abus_o[16] ),
        .O(abus_o[14]));
  LUT2 #(
    .INIT(4'h8)) 
    \abus_o[31]_INST_0 
       (.I0(\mul_a_reg[32] ),
        .I1(\abus_o[16] ),
        .O(abus_o[15]));
  LUT3 #(
    .INIT(8'h02)) 
    \badr[15]_INST_0_i_44 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(sr[8]),
        .O(\sr_reg[1]_5 ));
  LUT3 #(
    .INIT(8'h08)) 
    \badr[15]_INST_0_i_45 
       (.I0(sr[1]),
        .I1(sr[0]),
        .I2(sr[8]),
        .O(\sr_reg[1]_4 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \badr[15]_INST_0_i_46 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(sr[1]),
        .O(\sr_reg[0]_0 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[16]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [0]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [0]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_194 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[16]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [0]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [0]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_178 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[16]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [0]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [0]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_162 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[16]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [0]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [0]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_146 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[17]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [1]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [1]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_195 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[17]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [1]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [1]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_179 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[17]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [1]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [1]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_163 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[17]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [1]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [1]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_147 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[18]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [2]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [2]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_196 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[18]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [2]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [2]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_180 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[18]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [2]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [2]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_164 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[18]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [2]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [2]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_148 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[19]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [3]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [3]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_197 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[19]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [3]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [3]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_181 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[19]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [3]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [3]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_165 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[19]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [3]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [3]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_149 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[20]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [4]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [4]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_198 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[20]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [4]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [4]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_182 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[20]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [4]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [4]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_166 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[20]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [4]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [4]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_150 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[21]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [5]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [5]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_199 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[21]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [5]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [5]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_183 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[21]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [5]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [5]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_167 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[21]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [5]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [5]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_151 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[22]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [6]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [6]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_200 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[22]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [6]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [6]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_184 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[22]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [6]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [6]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_168 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[22]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [6]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [6]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_152 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[23]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [7]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [7]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_201 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[23]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [7]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [7]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_185 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[23]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [7]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [7]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_169 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[23]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [7]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [7]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_153 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[24]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [8]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [8]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_202 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[24]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [8]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [8]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_186 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[24]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [8]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [8]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_170 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[24]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [8]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [8]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_154 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[25]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [9]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [9]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_203 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[25]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [9]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [9]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_187 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[25]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [9]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [9]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_171 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[25]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [9]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [9]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_155 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[26]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [10]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [10]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_204 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[26]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [10]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [10]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_188 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[26]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [10]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [10]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_172 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[26]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [10]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [10]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_156 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[27]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [11]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [11]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_205 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[27]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [11]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [11]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_189 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[27]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [11]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [11]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_173 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[27]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [11]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [11]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_157 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[28]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [12]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [12]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_206 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[28]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [12]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [12]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_190 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[28]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [12]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [12]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_174 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[28]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [12]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [12]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_158 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[29]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [13]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [13]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_207 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[29]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [13]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [13]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_191 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[29]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [13]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [13]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_175 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[29]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [13]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [13]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_159 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[30]_INST_0_i_10 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [14]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [14]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_208 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[30]_INST_0_i_11 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [14]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [14]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_192 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[30]_INST_0_i_8 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [14]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [14]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_176 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[30]_INST_0_i_9 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [14]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [14]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_160 ));
  LUT6 #(
    .INIT(64'h000000007B4BBB8B)) 
    \badr[31]_INST_0_i_112 
       (.I0(sr[5]),
        .I1(\badr[31]_INST_0_i_69 [4]),
        .I2(\badr[31]_INST_0_i_69 [2]),
        .I3(sr[4]),
        .I4(sr[7]),
        .I5(\badr[31]_INST_0_i_69 [5]),
        .O(\sr_reg[5]_0 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[31]_INST_0_i_16 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_4 [15]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_4_0 [15]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_177 ));
  LUT6 #(
    .INIT(64'h2222200020002000)) 
    \badr[31]_INST_0_i_19 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_5 [15]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_5_0 [15]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_161 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[31]_INST_0_i_22 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_6 [15]),
        .I3(abus_sel_0[3]),
        .I4(\i_/badr[31]_INST_0_i_6_0 [15]),
        .I5(abus_sel_0[2]),
        .O(\sr_reg[8]_209 ));
  LUT6 #(
    .INIT(64'h8888800080008000)) 
    \badr[31]_INST_0_i_25 
       (.I0(sr[8]),
        .I1(sr[0]),
        .I2(\i_/badr[31]_INST_0_i_7 [15]),
        .I3(abus_sel_0[1]),
        .I4(\i_/badr[31]_INST_0_i_7_0 [15]),
        .I5(abus_sel_0[0]),
        .O(\sr_reg[8]_193 ));
  LUT5 #(
    .INIT(32'hBB2BFFFF)) 
    \bcmd[1]_INST_0_i_14 
       (.I0(irq_lev[1]),
        .I1(sr[3]),
        .I2(sr[2]),
        .I3(irq_lev[0]),
        .I4(irq),
        .O(irq_lev_1_sn_1));
  LUT5 #(
    .INIT(32'h5FCFA0CF)) 
    \bdatw[15]_INST_0_i_15 
       (.I0(sr[7]),
        .I1(sr[4]),
        .I2(\badr[31]_INST_0_i_69 [2]),
        .I3(\badr[31]_INST_0_i_69 [4]),
        .I4(sr[5]),
        .O(\sr_reg[7]_1 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [0]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [0]),
        .O(\sr_reg[0]_80 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[16]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [0]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [0]),
        .O(\sr_reg[0]_96 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [0]),
        .I5(\bdatw[31]_INST_0_i_4_0 [0]),
        .O(\sr_reg[0]_16 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [0]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [0]),
        .O(\sr_reg[0]_32 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [0]),
        .I5(\bdatw[31]_INST_0_i_4_2 [0]),
        .O(\sr_reg[0]_48 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[16]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [0]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [0]),
        .O(\sr_reg[0]_64 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [1]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [1]),
        .O(\sr_reg[0]_79 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[17]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [1]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [1]),
        .O(\sr_reg[0]_95 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [1]),
        .I5(\bdatw[31]_INST_0_i_4_0 [1]),
        .O(\sr_reg[0]_15 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [1]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [1]),
        .O(\sr_reg[0]_31 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [1]),
        .I5(\bdatw[31]_INST_0_i_4_2 [1]),
        .O(\sr_reg[0]_47 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[17]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [1]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [1]),
        .O(\sr_reg[0]_63 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [2]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [2]),
        .O(\sr_reg[0]_78 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[18]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [2]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [2]),
        .O(\sr_reg[0]_94 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [2]),
        .I5(\bdatw[31]_INST_0_i_4_0 [2]),
        .O(\sr_reg[0]_14 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [2]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [2]),
        .O(\sr_reg[0]_30 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [2]),
        .I5(\bdatw[31]_INST_0_i_4_2 [2]),
        .O(\sr_reg[0]_46 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[18]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [2]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [2]),
        .O(\sr_reg[0]_62 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [3]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [3]),
        .O(\sr_reg[0]_77 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[19]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [3]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [3]),
        .O(\sr_reg[0]_93 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [3]),
        .I5(\bdatw[31]_INST_0_i_4_0 [3]),
        .O(\sr_reg[0]_13 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [3]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [3]),
        .O(\sr_reg[0]_29 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [3]),
        .I5(\bdatw[31]_INST_0_i_4_2 [3]),
        .O(\sr_reg[0]_45 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[19]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [3]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [3]),
        .O(\sr_reg[0]_61 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [4]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [4]),
        .O(\sr_reg[0]_76 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[20]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [4]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [4]),
        .O(\sr_reg[0]_92 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [4]),
        .I5(\bdatw[31]_INST_0_i_4_0 [4]),
        .O(\sr_reg[0]_12 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [4]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [4]),
        .O(\sr_reg[0]_28 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [4]),
        .I5(\bdatw[31]_INST_0_i_4_2 [4]),
        .O(\sr_reg[0]_44 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[20]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [4]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [4]),
        .O(\sr_reg[0]_60 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [5]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [5]),
        .O(\sr_reg[0]_75 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[21]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [5]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [5]),
        .O(\sr_reg[0]_91 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [5]),
        .I5(\bdatw[31]_INST_0_i_4_0 [5]),
        .O(\sr_reg[0]_11 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [5]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [5]),
        .O(\sr_reg[0]_27 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [5]),
        .I5(\bdatw[31]_INST_0_i_4_2 [5]),
        .O(\sr_reg[0]_43 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[21]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [5]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [5]),
        .O(\sr_reg[0]_59 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [6]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [6]),
        .O(\sr_reg[0]_74 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[22]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [6]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [6]),
        .O(\sr_reg[0]_90 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [6]),
        .I5(\bdatw[31]_INST_0_i_4_0 [6]),
        .O(\sr_reg[0]_10 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [6]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [6]),
        .O(\sr_reg[0]_26 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [6]),
        .I5(\bdatw[31]_INST_0_i_4_2 [6]),
        .O(\sr_reg[0]_42 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[22]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [6]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [6]),
        .O(\sr_reg[0]_58 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [7]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [7]),
        .O(\sr_reg[0]_73 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[23]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [7]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [7]),
        .O(\sr_reg[0]_89 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [7]),
        .I5(\bdatw[31]_INST_0_i_4_0 [7]),
        .O(\sr_reg[0]_9 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [7]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [7]),
        .O(\sr_reg[0]_25 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [7]),
        .I5(\bdatw[31]_INST_0_i_4_2 [7]),
        .O(\sr_reg[0]_41 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[23]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [7]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [7]),
        .O(\sr_reg[0]_57 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [8]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [8]),
        .O(\sr_reg[0]_72 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[24]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [8]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [8]),
        .O(\sr_reg[0]_88 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [8]),
        .I5(\bdatw[31]_INST_0_i_4_0 [8]),
        .O(\sr_reg[0]_8 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [8]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [8]),
        .O(\sr_reg[0]_24 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [8]),
        .I5(\bdatw[31]_INST_0_i_4_2 [8]),
        .O(\sr_reg[0]_40 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[24]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [8]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [8]),
        .O(\sr_reg[0]_56 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [9]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [9]),
        .O(\sr_reg[0]_71 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[25]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [9]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [9]),
        .O(\sr_reg[0]_87 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [9]),
        .I5(\bdatw[31]_INST_0_i_4_0 [9]),
        .O(\sr_reg[0]_7 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [9]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [9]),
        .O(\sr_reg[0]_23 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [9]),
        .I5(\bdatw[31]_INST_0_i_4_2 [9]),
        .O(\sr_reg[0]_39 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[25]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [9]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [9]),
        .O(\sr_reg[0]_55 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [10]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [10]),
        .O(\sr_reg[0]_70 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[26]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [10]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [10]),
        .O(\sr_reg[0]_86 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [10]),
        .I5(\bdatw[31]_INST_0_i_4_0 [10]),
        .O(\sr_reg[0]_6 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [10]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [10]),
        .O(\sr_reg[0]_22 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [10]),
        .I5(\bdatw[31]_INST_0_i_4_2 [10]),
        .O(\sr_reg[0]_38 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[26]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [10]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [10]),
        .O(\sr_reg[0]_54 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [11]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [11]),
        .O(\sr_reg[0]_69 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[27]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [11]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [11]),
        .O(\sr_reg[0]_85 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [11]),
        .I5(\bdatw[31]_INST_0_i_4_0 [11]),
        .O(\sr_reg[0]_5 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [11]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [11]),
        .O(\sr_reg[0]_21 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [11]),
        .I5(\bdatw[31]_INST_0_i_4_2 [11]),
        .O(\sr_reg[0]_37 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[27]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [11]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [11]),
        .O(\sr_reg[0]_53 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [12]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [12]),
        .O(\sr_reg[0]_68 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[28]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [12]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [12]),
        .O(\sr_reg[0]_84 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [12]),
        .I5(\bdatw[31]_INST_0_i_4_0 [12]),
        .O(\sr_reg[0]_4 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [12]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [12]),
        .O(\sr_reg[0]_20 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [12]),
        .I5(\bdatw[31]_INST_0_i_4_2 [12]),
        .O(\sr_reg[0]_36 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[28]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [12]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [12]),
        .O(\sr_reg[0]_52 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [13]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [13]),
        .O(\sr_reg[0]_67 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[29]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [13]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [13]),
        .O(\sr_reg[0]_83 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [13]),
        .I5(\bdatw[31]_INST_0_i_4_0 [13]),
        .O(\sr_reg[0]_3 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [13]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [13]),
        .O(\sr_reg[0]_19 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [13]),
        .I5(\bdatw[31]_INST_0_i_4_2 [13]),
        .O(\sr_reg[0]_35 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[29]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [13]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [13]),
        .O(\sr_reg[0]_51 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [14]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [14]),
        .O(\sr_reg[0]_66 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[30]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [14]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [14]),
        .O(\sr_reg[0]_82 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_4 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [14]),
        .I5(\bdatw[31]_INST_0_i_4_0 [14]),
        .O(\sr_reg[0]_2 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_5 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [14]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [14]),
        .O(\sr_reg[0]_18 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_6 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [14]),
        .I5(\bdatw[31]_INST_0_i_4_2 [14]),
        .O(\sr_reg[0]_34 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[30]_INST_0_i_7 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [14]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [14]),
        .O(\sr_reg[0]_50 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_10 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_5 [15]),
        .I5(\i_/badr[31]_INST_0_i_5_0 [15]),
        .O(\sr_reg[0]_17 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_11 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[7]),
        .I3(bbus_sel_0[0]),
        .I4(\bdatw[31]_INST_0_i_4_1 [15]),
        .I5(\bdatw[31]_INST_0_i_4_2 [15]),
        .O(\sr_reg[0]_33 ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_12 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_4 [15]),
        .I5(\i_/badr[31]_INST_0_i_4_0 [15]),
        .O(\sr_reg[0]_49 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_42 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[1]),
        .I3(bbus_sel_0[2]),
        .I4(\i_/badr[31]_INST_0_i_7 [15]),
        .I5(\i_/badr[31]_INST_0_i_7_0 [15]),
        .O(\sr_reg[0]_65 ));
  LUT6 #(
    .INIT(64'h8880808088000000)) 
    \bdatw[31]_INST_0_i_45 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[5]),
        .I3(bbus_sel_0[6]),
        .I4(\i_/badr[31]_INST_0_i_6 [15]),
        .I5(\i_/badr[31]_INST_0_i_6_0 [15]),
        .O(\sr_reg[0]_81 ));
  LUT6 #(
    .INIT(64'h0400000044440400)) 
    \bdatw[31]_INST_0_i_61 
       (.I0(\stat[0]_i_6 [0]),
        .I1(irq),
        .I2(irq_lev[0]),
        .I3(sr[2]),
        .I4(sr[3]),
        .I5(irq_lev[1]),
        .O(\stat_reg[0] ));
  LUT6 #(
    .INIT(64'h4440404044000000)) 
    \bdatw[31]_INST_0_i_9 
       (.I0(sr[0]),
        .I1(sr[8]),
        .I2(bbus_sel_0[3]),
        .I3(bbus_sel_0[4]),
        .I4(\bdatw[31]_INST_0_i_4 [15]),
        .I5(\bdatw[31]_INST_0_i_4_0 [15]),
        .O(\sr_reg[0]_1 ));
  LUT6 #(
    .INIT(64'h00300F3F50305030)) 
    ctl_fetch_inferred_i_25
       (.I0(ctl_fetch_inferred_i_43_n_0),
        .I1(sr[4]),
        .I2(\badr[31]_INST_0_i_69 [2]),
        .I3(\badr[31]_INST_0_i_69 [4]),
        .I4(sr[6]),
        .I5(\badr[31]_INST_0_i_69 [3]),
        .O(\sr_reg[4]_0 ));
  LUT3 #(
    .INIT(8'h60)) 
    ctl_fetch_inferred_i_30
       (.I0(sr[5]),
        .I1(sr[7]),
        .I2(\badr[31]_INST_0_i_69 [4]),
        .O(\sr_reg[5]_1 ));
  LUT3 #(
    .INIT(8'h31)) 
    ctl_fetch_inferred_i_40
       (.I0(sr[8]),
        .I1(\badr[31]_INST_0_i_69 [0]),
        .I2(\stat[0]_i_6 [0]),
        .O(\sr_reg[8]_132 ));
  LUT2 #(
    .INIT(4'h6)) 
    ctl_fetch_inferred_i_43
       (.I0(sr[7]),
        .I1(sr[5]),
        .O(ctl_fetch_inferred_i_43_n_0));
  LUT4 #(
    .INIT(16'hBF0B)) 
    ctl_fetch_inferred_i_52
       (.I0(irq_lev[0]),
        .I1(sr[2]),
        .I2(sr[3]),
        .I3(irq_lev[1]),
        .O(irq_lev_0_sn_1));
  LUT5 #(
    .INIT(32'h2000AA20)) 
    fch_irq_req_fl_i_1
       (.I0(irq),
        .I1(irq_lev[0]),
        .I2(sr[2]),
        .I3(sr[3]),
        .I4(irq_lev[1]),
        .O(fch_irq_req));
  LUT4 #(
    .INIT(16'h0D00)) 
    \grn[15]_i_1 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(cbus_sel_0),
        .O(\sr_reg[1]_0 ));
  LUT4 #(
    .INIT(16'hE000)) 
    \grn[15]_i_1__0 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(cbus_sel_0),
        .O(\sr_reg[1]_1 ));
  LUT4 #(
    .INIT(16'h0E00)) 
    \grn[15]_i_1__1 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(cbus_sel_0),
        .O(\sr_reg[1]_2 ));
  LUT5 #(
    .INIT(32'h00001101)) 
    \grn[15]_i_1__10 
       (.I0(\grn_reg[0] ),
        .I1(\grn_reg[0]_0 ),
        .I2(sr[1]),
        .I3(sr[8]),
        .I4(sr[0]),
        .O(\sr_reg[1]_8 ));
  LUT4 #(
    .INIT(16'hD000)) 
    \grn[15]_i_1__2 
       (.I0(sr[1]),
        .I1(sr[8]),
        .I2(sr[0]),
        .I3(cbus_sel_0),
        .O(\sr_reg[1]_3 ));
  LUT5 #(
    .INIT(32'h11010000)) 
    \grn[15]_i_1__7 
       (.I0(\grn_reg[0] ),
        .I1(\grn_reg[0]_0 ),
        .I2(sr[1]),
        .I3(sr[8]),
        .I4(sr[0]),
        .O(E));
  LUT5 #(
    .INIT(32'h00001110)) 
    \grn[15]_i_1__8 
       (.I0(\grn_reg[0] ),
        .I1(\grn_reg[0]_0 ),
        .I2(sr[1]),
        .I3(sr[8]),
        .I4(sr[0]),
        .O(\sr_reg[1]_6 ));
  LUT5 #(
    .INIT(32'h11100000)) 
    \grn[15]_i_1__9 
       (.I0(\grn_reg[0] ),
        .I1(\grn_reg[0]_0 ),
        .I2(sr[1]),
        .I3(sr[8]),
        .I4(sr[0]),
        .O(\sr_reg[1]_7 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[0]_i_11 
       (.I0(\mul_a_reg[24] ),
        .I1(\iv[5]_i_7 ),
        .I2(\niho_dsp_a[3] [0]),
        .O(\badr[0]_INST_0_i_1 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \iv[0]_i_24 
       (.I0(\sr[4]_i_91 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\sr_reg[8]_45 ),
        .I3(\iv[0]_i_21 ),
        .I4(\sr_reg[8]_46 ),
        .O(\sr_reg[8]_44 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_25 
       (.I0(\iv[0]_i_33_n_0 ),
        .I1(\iv[0]_i_34_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[4]_i_36_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\sr_reg[8]_82 ),
        .O(\sr_reg[8]_71 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_26 
       (.I0(\iv[12]_i_39_n_0 ),
        .I1(\iv[12]_i_40_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[0]_i_35_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[0]_i_36_n_0 ),
        .O(\sr_reg[8]_70 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[0]_i_29 
       (.I0(\iv[12]_i_48_n_0 ),
        .I1(\sr_reg[8]_100 ),
        .I2(\iv[0]_i_21 ),
        .I3(\sr_reg[8]_97 ),
        .I4(\iv[9]_i_28 ),
        .I5(\iv[12]_i_47_n_0 ),
        .O(\sr_reg[8]_99 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[0]_i_31 
       (.I0(\iv[0]_i_37_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[12]_i_41_n_0 ),
        .O(\sr_reg[8]_45 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[0]_i_32 
       (.I0(\iv[12]_i_42_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr[7]_i_48_n_0 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\iv[8]_i_27 ),
        .O(\sr_reg[8]_46 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_33 
       (.I0(sr[8]),
        .I1(\mul_a_reg[22] ),
        .I2(\mul_a_reg[23] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[0]_i_33_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_34 
       (.I0(sr[8]),
        .I1(\mul_a_reg[20] ),
        .I2(\mul_a_reg[21] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[0]_i_34_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_35 
       (.I0(sr[8]),
        .I1(\mul_a_reg[26] ),
        .I2(\mul_a_reg[27] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[0]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[0]_i_36 
       (.I0(sr[8]),
        .I1(\mul_a_reg[24] ),
        .I2(\mul_a_reg[25] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[0]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[0]_i_37 
       (.I0(\sr[7]_i_50_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\sr[7]_i_51_n_0 ),
        .O(\iv[0]_i_37_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \iv[0]_i_8 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_42_0 ),
        .I2(\iv[0]_i_3 ),
        .I3(\sr_reg[8]_14 ),
        .I4(\iv[0]_i_3_0 ),
        .I5(\iv[0]_i_3_1 ),
        .O(\sr_reg[8]_16 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[10]_i_10 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[10]_i_4 ),
        .I2(\iv[13]_i_4_0 ),
        .I3(\iv[10]_i_23_n_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_17 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[10]_i_13 
       (.I0(\sr_reg[8]_59 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\iv[10]_i_6 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_60 ),
        .I5(\sr[4]_i_91 ),
        .O(\sr_reg[8]_58 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_23 
       (.I0(\iv[10]_i_41_n_0 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr_reg[8]_40 ),
        .O(\iv[10]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[10]_i_25 
       (.I0(\sr[7]_i_30_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr[7]_i_26_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[27]_i_7 ),
        .O(\sr_reg[8]_216 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \iv[10]_i_26 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[8]_77 ),
        .O(\sr_reg[8]_59 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_28 
       (.I0(\iv[14]_i_56_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[14]_i_52_n_0 ),
        .O(\sr_reg[8]_60 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[10]_i_29 
       (.I0(\iv[10]_i_44_n_0 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\tr[26]_i_6 ),
        .O(\iv[10]_i_34 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[10]_i_40 
       (.I0(\iv[0]_i_34_n_0 ),
        .I1(\iv[4]_i_36_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[0]_i_36_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[0]_i_33_n_0 ),
        .O(\sr_reg[8]_81 ));
  LUT6 #(
    .INIT(64'hFA0AFCFCFA0A0C0C)) 
    \iv[10]_i_41 
       (.I0(\iv[12]_i_40_n_0 ),
        .I1(\iv[0]_i_35_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[12]_i_39_n_0 ),
        .O(\iv[10]_i_41_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \iv[10]_i_44 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[10]_i_29_0 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\iv[12]_i_51_n_0 ),
        .O(\iv[10]_i_44_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[11]_i_10 
       (.I0(\sr[5]_i_3_0 ),
        .I1(\mul_a_reg[32] ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[11]_i_23_n_0 ),
        .I4(\iv[11]_i_4_0 ),
        .I5(\sr[5]_i_3_5 ),
        .O(\iv[11]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[11]_i_11 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[11]_i_23_n_0 ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[11]_i_24_n_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\iv[11]_i_11_n_0 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[11]_i_13 
       (.I0(\sr_reg[8]_56 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\sr[4]_i_91_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_57 ),
        .I5(\sr[4]_i_91 ),
        .O(\sr_reg[8]_55 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[11]_i_23 
       (.I0(\iv[9]_i_28 ),
        .I1(\iv[11]_i_10_0 ),
        .I2(\sr_reg[8]_107 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\iv[11]_i_42_n_0 ),
        .O(\iv[11]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \iv[11]_i_24 
       (.I0(\iv[9]_i_28 ),
        .I1(\iv[15]_i_131_n_0 ),
        .I2(\tr[28]_i_8_0 ),
        .I3(\iv[15]_i_132_n_0 ),
        .I4(\sr[6]_i_11_0 ),
        .I5(\sr_reg[8]_40 ),
        .O(\iv[11]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \iv[11]_i_25 
       (.I0(\iv[15]_i_136_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[15]_i_138_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[28]_i_9 ),
        .O(\sr_reg[8]_215 ));
  LUT5 #(
    .INIT(32'hFBFFFB00)) 
    \iv[11]_i_27 
       (.I0(bbus_0[0]),
        .I1(\mul_a_reg[32] ),
        .I2(niho_dsp_b_0_sn_1),
        .I3(\iv[9]_i_28 ),
        .I4(\sr_reg[8]_94 ),
        .O(\sr_reg[8]_56 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_29 
       (.I0(\iv[11]_i_47_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[8]_93 ),
        .O(\sr_reg[8]_57 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[11]_i_4 
       (.I0(\sr[4]_i_19_1 ),
        .I1(\iv[11]_i_10_n_0 ),
        .I2(\iv[11]_i_11_n_0 ),
        .O(\iv[11]_i_11_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[11]_i_41 
       (.I0(\sr_reg[8]_90 ),
        .I1(\tr[28]_i_8_0 ),
        .I2(\sr_reg[8]_91 ),
        .O(\sr_reg[8]_107 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[11]_i_42 
       (.I0(\iv[15]_i_133_n_0 ),
        .I1(\iv[15]_i_134_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[15]_i_127_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[15]_i_128_n_0 ),
        .O(\iv[11]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[11]_i_45 
       (.I0(\iv[15]_i_141_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[13]_i_51_n_0 ),
        .O(\sr_reg[8]_94 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[11]_i_46 
       (.I0(\mul_a_reg[17] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[18] ),
        .O(\badr[18]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[11]_i_47 
       (.I0(\iv[13]_i_52_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[13]_i_53_n_0 ),
        .O(\iv[11]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[12]_i_10 
       (.I0(\sr_reg[8]_14 ),
        .I1(\sr_reg[8]_33 ),
        .I2(\iv[13]_i_4_0 ),
        .I3(\iv[12]_i_23_n_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_32 ));
  LUT5 #(
    .INIT(32'hB1FFB100)) 
    \iv[12]_i_21 
       (.I0(\iv[9]_i_28 ),
        .I1(\iv[12]_i_9 ),
        .I2(\sr_reg[8]_101 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\iv[12]_i_38_n_0 ),
        .O(\sr_reg[8]_33 ));
  LUT6 #(
    .INIT(64'hFFB8FFFF00B80000)) 
    \iv[12]_i_23 
       (.I0(\iv[12]_i_39_n_0 ),
        .I1(\tr[28]_i_8_0 ),
        .I2(\iv[12]_i_40_n_0 ),
        .I3(\iv[9]_i_28 ),
        .I4(\sr[6]_i_11_0 ),
        .I5(\sr_reg[8]_40 ),
        .O(\iv[12]_i_23_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[12]_i_24 
       (.I0(\iv[12]_i_41_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[12]_i_42_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\iv[12]_i_43_n_0 ),
        .O(\sr_reg[8]_227 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[12]_i_28 
       (.I0(\iv[12]_i_47_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[12]_i_48_n_0 ),
        .O(\sr_reg[8]_98 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[12]_i_38 
       (.I0(\iv[0]_i_35_n_0 ),
        .I1(\iv[0]_i_36_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[0]_i_33_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[0]_i_34_n_0 ),
        .O(\iv[12]_i_38_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[12]_i_39 
       (.I0(sr[8]),
        .I1(\mul_a_reg[30] ),
        .I2(\mul_a_reg[32] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[12]_i_39_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[12]_i_40 
       (.I0(sr[8]),
        .I1(\mul_a_reg[28] ),
        .I2(\mul_a_reg[29] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[12]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_41 
       (.I0(\sr[7]_i_52_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\sr[7]_i_45_n_0 ),
        .O(\iv[12]_i_41_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_42 
       (.I0(\sr[7]_i_46_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\sr[7]_i_47_n_0 ),
        .O(\iv[12]_i_42_n_0 ));
  LUT5 #(
    .INIT(32'hE2EEE222)) 
    \iv[12]_i_43 
       (.I0(\iv[0]_i_37_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[4]_i_27_0 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\badr[16]_INST_0_i_1 ),
        .O(\iv[12]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'h30303F305F505F50)) 
    \iv[12]_i_44 
       (.I0(\mul_a_reg[32] ),
        .I1(\mul_a_reg[30] ),
        .I2(\tr[28]_i_8_0 ),
        .I3(\iv[12]_i_25 ),
        .I4(sr[6]),
        .I5(niho_dsp_b_0_sn_1),
        .O(\sr_reg[6]_2 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_45 
       (.I0(\iv[12]_i_51_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[14]_i_67_n_0 ),
        .O(\sr_reg[8]_97 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_46 
       (.I0(\iv[14]_i_66_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\badr[16]_INST_0_i_1_0 ),
        .O(\sr_reg[8]_100 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_47 
       (.I0(\iv[14]_i_68_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[14]_i_69_n_0 ),
        .O(\iv[12]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[12]_i_48 
       (.I0(\iv[14]_i_70_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[14]_i_65_n_0 ),
        .O(\iv[12]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[12]_i_51 
       (.I0(\mul_a_reg[32] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[30] ),
        .O(\iv[12]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[13]_i_10 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[13]_i_22_n_0 ),
        .I2(\iv[13]_i_4_0 ),
        .I3(\sr_reg[8]_34 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\iv[13]_i_10_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_22 
       (.I0(\sr_reg[8]_89 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\iv[13]_i_40_n_0 ),
        .O(\iv[13]_i_22_n_0 ));
  LUT5 #(
    .INIT(32'hCDC8CCCC)) 
    \iv[13]_i_24 
       (.I0(\tr[23]_i_6_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\tr[28]_i_8_0 ),
        .I3(\iv[15]_i_131_n_0 ),
        .I4(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_34 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \iv[13]_i_26 
       (.I0(\iv[13]_i_42_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[30]_i_10 ),
        .O(\sr_reg[8]_210 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[13]_i_30 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[13]_i_49_n_0 ),
        .O(\sr_reg[8]_76 ));
  LUT3 #(
    .INIT(8'h8A)) 
    \iv[13]_i_4 
       (.I0(\sr[4]_i_19_1 ),
        .I1(\iv[13]_i_9_n_0 ),
        .I2(\iv[13]_i_10_n_0 ),
        .O(\iv[13]_i_10_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[13]_i_40 
       (.I0(\iv[15]_i_132_n_0 ),
        .I1(\iv[15]_i_133_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[15]_i_134_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[15]_i_127_n_0 ),
        .O(\iv[13]_i_40_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_42 
       (.I0(\iv[15]_i_166_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_163_n_0 ),
        .O(\iv[13]_i_42_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_43 
       (.I0(\iv[15]_i_170_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_165_n_0 ),
        .O(\iv[13]_i_43_n_0 ));
  LUT6 #(
    .INIT(64'hDDDDFFFFDDD1000C)) 
    \iv[13]_i_45 
       (.I0(\mul_a_reg[32] ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_141_n_0 ),
        .O(\sr_reg[8]_84 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_47 
       (.I0(\iv[7]_i_48_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\badr[18]_INST_0_i_1 ),
        .O(\sr_reg[8]_86 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_48 
       (.I0(\iv[13]_i_51_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[13]_i_52_n_0 ),
        .O(\iv[13]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[13]_i_49 
       (.I0(\iv[13]_i_53_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[7]_i_47_n_0 ),
        .O(\iv[13]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[13]_i_51 
       (.I0(\mul_a_reg[27] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[28] ),
        .O(\iv[13]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[13]_i_52 
       (.I0(\mul_a_reg[25] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[26] ),
        .O(\iv[13]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[13]_i_53 
       (.I0(\mul_a_reg[23] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[24] ),
        .O(\iv[13]_i_53_n_0 ));
  LUT6 #(
    .INIT(64'h8A80FFFF8A808A80)) 
    \iv[13]_i_9 
       (.I0(\sr[5]_i_3_0 ),
        .I1(\mul_a_reg[32] ),
        .I2(\iv[13]_i_4_0 ),
        .I3(\iv[13]_i_22_n_0 ),
        .I4(\iv[13]_i_4_1 ),
        .I5(\sr[5]_i_3_5 ),
        .O(\iv[13]_i_9_n_0 ));
  LUT4 #(
    .INIT(16'h57F7)) 
    \iv[14]_i_11 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[14]_i_27_n_0 ),
        .I2(\sr[4]_i_42_0 ),
        .I3(\mul_a_reg[32] ),
        .O(\iv[14]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_27 
       (.I0(\sr_reg[8]_62 ),
        .I1(\tr[23]_i_3 ),
        .I2(\sr_reg[8]_63 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\iv[14]_i_50_n_0 ),
        .O(\iv[14]_i_27_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[14]_i_29 
       (.I0(\iv[14]_i_52_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\badr[16]_INST_0_i_1_0 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\iv[14]_i_13 ),
        .O(\sr_reg[8]_74 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[14]_i_30 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[14]_i_56_n_0 ),
        .O(\sr_reg[8]_108 ));
  LUT5 #(
    .INIT(32'h8A88AAAA)) 
    \iv[14]_i_4 
       (.I0(\sr[4]_i_19_1 ),
        .I1(\iv[15]_i_54_n_0 ),
        .I2(\iv[14]_i_2 ),
        .I3(\sr[5]_i_3_5 ),
        .I4(\iv[14]_i_11_n_0 ),
        .O(\iv[14]_i_11_0 ));
  LUT6 #(
    .INIT(64'hAFAFA0A0C0CFC0CF)) 
    \iv[14]_i_49 
       (.I0(\iv[0]_i_34_n_0 ),
        .I1(\iv[4]_i_36_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[14]_i_13 ),
        .I4(\sr_reg[8]_82 ),
        .I5(\tr[28]_i_8_0 ),
        .O(\sr_reg[8]_63 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[14]_i_50 
       (.I0(\iv[12]_i_40_n_0 ),
        .I1(\iv[0]_i_35_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[0]_i_36_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[0]_i_33_n_0 ),
        .O(\iv[14]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'hA9A9AAFFFFFFAAFF)) 
    \iv[14]_i_51 
       (.I0(bbus_0[0]),
        .I1(\sr_reg[8]_79 ),
        .I2(\sr_reg[8]_80 ),
        .I3(\mul_a_reg[30] ),
        .I4(niho_dsp_b_0_sn_1),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_77 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[14]_i_52 
       (.I0(\iv[14]_i_65_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[14]_i_66_n_0 ),
        .O(\iv[14]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[14]_i_53 
       (.I0(\mul_a_reg[17] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[16] ),
        .O(\badr[16]_INST_0_i_1_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[14]_i_55 
       (.I0(\iv[14]_i_67_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[14]_i_68_n_0 ),
        .O(\iv[14]_i_55_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[14]_i_56 
       (.I0(\iv[14]_i_69_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[14]_i_70_n_0 ),
        .O(\iv[14]_i_56_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_65 
       (.I0(\mul_a_reg[20] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[21] ),
        .O(\iv[14]_i_65_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_66 
       (.I0(\mul_a_reg[18] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[19] ),
        .O(\iv[14]_i_66_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[14]_i_67 
       (.I0(\mul_a_reg[29] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[28] ),
        .O(\iv[14]_i_67_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_68 
       (.I0(\mul_a_reg[26] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[27] ),
        .O(\iv[14]_i_68_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[14]_i_69 
       (.I0(\mul_a_reg[25] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[24] ),
        .O(\iv[14]_i_69_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[14]_i_70 
       (.I0(\mul_a_reg[22] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[23] ),
        .O(\iv[14]_i_70_n_0 ));
  LUT6 #(
    .INIT(64'h5F50CFCF5F50C0C0)) 
    \iv[15]_i_101 
       (.I0(\iv[15]_i_141_n_0 ),
        .I1(\iv[15]_i_142_n_0 ),
        .I2(\tr[23]_i_6_0 ),
        .I3(\iv[15]_i_143_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[15]_i_144_n_0 ),
        .O(\sr_reg[8]_51 ));
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \iv[15]_i_102 
       (.I0(\iv[15]_i_145_n_0 ),
        .I1(\iv[15]_i_146_n_0 ),
        .I2(\tr[23]_i_6_0 ),
        .I3(\iv[15]_i_147_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[15]_i_58 ),
        .O(\sr_reg[8]_50 ));
  LUT2 #(
    .INIT(4'h2)) 
    \iv[15]_i_105 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_139_0 ),
        .O(\iv[8]_i_34 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_127 
       (.I0(sr[8]),
        .I1(\mul_a_reg[21] ),
        .I2(\mul_a_reg[22] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[15]_i_127_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_128 
       (.I0(sr[8]),
        .I1(\mul_a_reg[19] ),
        .I2(\mul_a_reg[20] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[15]_i_128_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_129 
       (.I0(sr[8]),
        .I1(\mul_a_reg[17] ),
        .I2(\mul_a_reg[18] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\sr_reg[8]_90 ));
  LUT4 #(
    .INIT(16'hDF80)) 
    \iv[15]_i_130 
       (.I0(sr[8]),
        .I1(\mul_a_reg[16] ),
        .I2(niho_dsp_b_0_sn_1),
        .I3(DI[3]),
        .O(\sr_reg[8]_91 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_131 
       (.I0(sr[8]),
        .I1(\mul_a_reg[29] ),
        .I2(\mul_a_reg[30] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[15]_i_131_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_132 
       (.I0(sr[8]),
        .I1(\mul_a_reg[27] ),
        .I2(\mul_a_reg[28] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[15]_i_132_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_133 
       (.I0(sr[8]),
        .I1(\mul_a_reg[25] ),
        .I2(\mul_a_reg[26] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[15]_i_133_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[15]_i_134 
       (.I0(sr[8]),
        .I1(\mul_a_reg[23] ),
        .I2(\mul_a_reg[24] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[15]_i_134_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_135 
       (.I0(\iv[15]_i_163_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_164_n_0 ),
        .O(\sr_reg[8]_104 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_136 
       (.I0(\iv[15]_i_165_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_166_n_0 ),
        .O(\iv[15]_i_136_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_137 
       (.I0(\badr[17]_INST_0_i_1 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_168_n_0 ),
        .O(\sr_reg[8]_105 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[15]_i_138 
       (.I0(\iv[15]_i_169_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_170_n_0 ),
        .O(\iv[15]_i_138_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_141 
       (.I0(\mul_a_reg[29] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[30] ),
        .O(\iv[15]_i_141_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_142 
       (.I0(\mul_a_reg[28] ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\mul_a_reg[27] ),
        .O(\iv[15]_i_142_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_143 
       (.I0(\mul_a_reg[26] ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\mul_a_reg[25] ),
        .O(\iv[15]_i_143_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_144 
       (.I0(\mul_a_reg[24] ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\mul_a_reg[23] ),
        .O(\iv[15]_i_144_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_145 
       (.I0(\mul_a_reg[22] ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\mul_a_reg[21] ),
        .O(\iv[15]_i_145_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_146 
       (.I0(\mul_a_reg[20] ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\mul_a_reg[19] ),
        .O(\iv[15]_i_146_n_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[15]_i_147 
       (.I0(\mul_a_reg[18] ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\mul_a_reg[17] ),
        .O(\iv[15]_i_147_n_0 ));
  LUT6 #(
    .INIT(64'h3333333333333335)) 
    \iv[15]_i_156 
       (.I0(\mul_a_reg[32] ),
        .I1(sr[6]),
        .I2(\iv[13]_i_45_0 ),
        .I3(\iv[13]_i_45_1 ),
        .I4(\iv[10]_i_44_1 ),
        .I5(\iv[10]_i_44_2 ),
        .O(\sr_reg[6]_1 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[15]_i_163 
       (.I0(\mul_a_reg[29] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[30] ),
        .O(\iv[15]_i_163_n_0 ));
  LUT6 #(
    .INIT(64'h5555555455555557)) 
    \iv[15]_i_164 
       (.I0(\mul_a_reg[32] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(sr[6]),
        .O(\iv[15]_i_164_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_165 
       (.I0(\mul_a_reg[26] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[25] ),
        .O(\iv[15]_i_165_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_166 
       (.I0(\mul_a_reg[28] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[27] ),
        .O(\iv[15]_i_166_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_167 
       (.I0(\mul_a_reg[18] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[17] ),
        .O(\badr[17]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_168 
       (.I0(\mul_a_reg[20] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[19] ),
        .O(\iv[15]_i_168_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_169 
       (.I0(\mul_a_reg[22] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[21] ),
        .O(\iv[15]_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[15]_i_170 
       (.I0(\mul_a_reg[24] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[23] ),
        .O(\iv[15]_i_170_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \iv[15]_i_21 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_42_0 ),
        .I2(\iv[15]_i_51_n_0 ),
        .I3(\sr_reg[8]_14 ),
        .I4(\iv[15]_i_8 ),
        .I5(\iv[15]_i_54_n_0 ),
        .O(\sr_reg[8]_41 ));
  LUT6 #(
    .INIT(64'hBBBBBBBBBBBBABAA)) 
    \iv[15]_i_23 
       (.I0(sr[8]),
        .I1(\iv[15]_i_8_0 ),
        .I2(\sr[4]_i_38_0 ),
        .I3(\iv[15]_i_62_n_0 ),
        .I4(\iv[15]_i_8_1 ),
        .I5(\iv[15]_i_8_2 ),
        .O(\sr_reg[8]_47 ));
  LUT5 #(
    .INIT(32'hFFB800B8)) 
    \iv[15]_i_51 
       (.I0(\sr_reg[8]_49 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\iv[15]_i_95_n_0 ),
        .I3(\tr[23]_i_3 ),
        .I4(\sr_reg[8]_40 ),
        .O(\iv[15]_i_51_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \iv[15]_i_52 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5] ),
        .O(\sr_reg[8]_14 ));
  LUT6 #(
    .INIT(64'h8A8A8A8080808A80)) 
    \iv[15]_i_54 
       (.I0(\sr[5]_i_3_0 ),
        .I1(\mul_a_reg[32] ),
        .I2(\tr[23]_i_3 ),
        .I3(\iv[15]_i_95_n_0 ),
        .I4(\sr[6]_i_11_0 ),
        .I5(\sr_reg[8]_49 ),
        .O(\iv[15]_i_54_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \iv[15]_i_56 
       (.I0(sr[8]),
        .I1(\iv[15]_i_96 ),
        .I2(\iv[15]_i_96_0 ),
        .I3(\iv[15]_i_96_1 ),
        .I4(\iv[15]_i_96_2 ),
        .I5(\iv[15]_i_96_3 ),
        .O(\sr_reg[8]_79 ));
  LUT6 #(
    .INIT(64'hFFFF00FF47474747)) 
    \iv[15]_i_62 
       (.I0(\sr_reg[8]_50 ),
        .I1(\iv[0]_i_21 ),
        .I2(\sr_reg[8]_51 ),
        .I3(\iv[8]_i_34 ),
        .I4(bbus_0[1]),
        .I5(\tr[23]_i_3 ),
        .O(\iv[15]_i_62_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_94 
       (.I0(\iv[15]_i_127_n_0 ),
        .I1(\iv[15]_i_128_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\sr_reg[8]_90 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\sr_reg[8]_91 ),
        .O(\sr_reg[8]_49 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[15]_i_95 
       (.I0(\iv[15]_i_131_n_0 ),
        .I1(\iv[15]_i_132_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[15]_i_133_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[15]_i_134_n_0 ),
        .O(\iv[15]_i_95_n_0 ));
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \iv[15]_i_97 
       (.I0(\sr_reg[8]_104 ),
        .I1(\iv[15]_i_136_n_0 ),
        .I2(\iv[0]_i_21 ),
        .I3(\sr_reg[8]_105 ),
        .I4(\iv[9]_i_28 ),
        .I5(\iv[15]_i_138_n_0 ),
        .O(\sr_reg[8]_103 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[1]_i_11 
       (.I0(\mul_a_reg[25] ),
        .I1(\iv[5]_i_7 ),
        .I2(\niho_dsp_a[3] [1]),
        .O(\badr[1]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[1]_i_15 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[1]_i_8 ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[9]_i_46_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_37 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[1]_i_24 
       (.I0(\sr_reg[8]_69 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\iv[9]_i_46_n_0 ),
        .O(\iv[9]_i_46_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \iv[1]_i_26 
       (.I0(\sr_reg[8]_88 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\sr_reg[8]_87 ),
        .I4(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_212 ));
  LUT6 #(
    .INIT(64'h55335533000FFF0F)) 
    \iv[1]_i_27 
       (.I0(\iv[13]_i_49_n_0 ),
        .I1(\sr_reg[8]_86 ),
        .I2(\iv[13]_i_48_n_0 ),
        .I3(\iv[9]_i_28 ),
        .I4(\sr_reg[8]_84 ),
        .I5(\iv[0]_i_21 ),
        .O(\sr_reg[8]_85 ));
  LUT5 #(
    .INIT(32'hFF00E2E2)) 
    \iv[1]_i_28 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[6]_0 ),
        .I3(\sr_reg[8]_66 ),
        .I4(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_135 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[2]_i_11 
       (.I0(\mul_a_reg[26] ),
        .I1(\iv[5]_i_7 ),
        .I2(\niho_dsp_a[3] [2]),
        .O(\badr[2]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[2]_i_15 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[2]_i_8 ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[10]_i_41_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_36 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[2]_i_23 
       (.I0(\sr_reg[8]_81 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\iv[10]_i_41_n_0 ),
        .O(\iv[10]_i_41_0 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \iv[2]_i_24 
       (.I0(\sr[7]_i_30_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr[7]_i_26_n_0 ),
        .I3(\tr[18]_i_9 ),
        .I4(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_217 ));
  LUT6 #(
    .INIT(64'h55335533000FFF0F)) 
    \iv[2]_i_27 
       (.I0(\iv[14]_i_56_n_0 ),
        .I1(\iv[14]_i_52_n_0 ),
        .I2(\iv[14]_i_55_n_0 ),
        .I3(\iv[9]_i_28 ),
        .I4(\sr_reg[8]_77 ),
        .I5(\iv[0]_i_21 ),
        .O(\sr_reg[8]_78 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[2]_i_28 
       (.I0(\sr_reg[8]_60 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\iv[10]_i_44_n_0 ),
        .O(\iv[10]_i_44_0 ));
  LUT3 #(
    .INIT(8'h53)) 
    \iv[3]_i_12 
       (.I0(\mul_a_reg[27] ),
        .I1(\niho_dsp_a[3] [3]),
        .I2(\iv[5]_i_7 ),
        .O(\sr[6]_i_13 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[3]_i_16 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[3]_i_8 ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[3]_i_41_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_35 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[3]_i_29 
       (.I0(\iv[11]_i_42_n_0 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\iv[3]_i_41_n_0 ),
        .O(\iv[3]_i_41_0 ));
  LUT5 #(
    .INIT(32'hFF00E2E2)) 
    \iv[3]_i_31 
       (.I0(\iv[15]_i_136_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[15]_i_138_n_0 ),
        .I3(\tr[19]_i_7 ),
        .I4(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_214 ));
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \iv[3]_i_32 
       (.I0(\iv[11]_i_47_n_0 ),
        .I1(\sr_reg[8]_93 ),
        .I2(\iv[3]_i_42_n_0 ),
        .I3(\iv[9]_i_28 ),
        .I4(\sr_reg[8]_94 ),
        .I5(\iv[0]_i_21 ),
        .O(\sr_reg[8]_92 ));
  LUT5 #(
    .INIT(32'hCFCAC5C0)) 
    \iv[3]_i_33 
       (.I0(\iv[9]_i_28 ),
        .I1(\sr_reg[8]_57 ),
        .I2(\sr[6]_i_11_0 ),
        .I3(\sr_reg[8]_94 ),
        .I4(\tr[19]_i_6 ),
        .O(\sr_reg[8]_138 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[3]_i_41 
       (.I0(\sr_reg[8]_40 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[15]_i_131_n_0 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\iv[15]_i_132_n_0 ),
        .O(\iv[3]_i_41_n_0 ));
  LUT3 #(
    .INIT(8'hFB)) 
    \iv[3]_i_42 
       (.I0(bbus_0[0]),
        .I1(\mul_a_reg[32] ),
        .I2(niho_dsp_b_0_sn_1),
        .O(\iv[3]_i_42_n_0 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[4]_i_11 
       (.I0(\mul_a_reg[28] ),
        .I1(\iv[5]_i_7 ),
        .I2(\niho_dsp_a[7] [0]),
        .O(\badr[4]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[4]_i_14 
       (.I0(\sr_reg[8]_14 ),
        .I1(\sr[4]_i_32 ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[4]_i_35_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_21 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_22 
       (.I0(\iv[12]_i_38_n_0 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\iv[4]_i_35_n_0 ),
        .O(\iv[4]_i_35_0 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_26 
       (.I0(\iv[4]_i_36_n_0 ),
        .I1(\tr[28]_i_8_0 ),
        .I2(\sr_reg[8]_82 ),
        .O(\sr_reg[8]_101 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_27 
       (.I0(\iv[12]_i_43_n_0 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\tr[21]_i_9 ),
        .O(\iv[13]_i_35 ));
  LUT6 #(
    .INIT(64'hFFCC3300B8B8B8B8)) 
    \iv[4]_i_29 
       (.I0(\iv[12]_i_41_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[12]_i_42_n_0 ),
        .I3(\tr[20]_i_9 ),
        .I4(\sr_reg[6]_2 ),
        .I5(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_226 ));
  LUT5 #(
    .INIT(32'h5353000F)) 
    \iv[4]_i_30 
       (.I0(\iv[12]_i_47_n_0 ),
        .I1(\iv[12]_i_48_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\sr_reg[8]_97 ),
        .I4(\iv[0]_i_21 ),
        .O(\sr_reg[8]_96 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[4]_i_31 
       (.I0(\sr_reg[8]_98 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\tr[20]_i_8 ),
        .O(\iv[12]_i_49 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[4]_i_35 
       (.I0(\sr_reg[8]_40 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[12]_i_39_n_0 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\iv[12]_i_40_n_0 ),
        .O(\iv[4]_i_35_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[4]_i_36 
       (.I0(sr[8]),
        .I1(\mul_a_reg[18] ),
        .I2(\mul_a_reg[19] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\iv[4]_i_36_n_0 ));
  LUT5 #(
    .INIT(32'hFFFFA088)) 
    \iv[4]_i_37 
       (.I0(sr[8]),
        .I1(\mul_a_reg[16] ),
        .I2(\mul_a_reg[17] ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(niho_dsp_a_15_sn_1),
        .O(\sr_reg[8]_82 ));
  LUT6 #(
    .INIT(64'h0002220222222222)) 
    \iv[4]_i_8 
       (.I0(\sr_reg[8]_21 ),
        .I1(\iv[4]_i_3 ),
        .I2(\sr[4]_i_32 ),
        .I3(\sr[4]_i_91 ),
        .I4(\mul_a_reg[32] ),
        .I5(\sr[5]_i_3_0 ),
        .O(\sr_reg[8]_20 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[5]_i_11 
       (.I0(\mul_a_reg[29] ),
        .I1(\iv[5]_i_7 ),
        .I2(\niho_dsp_a[7] [1]),
        .O(\badr[5]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[5]_i_14 
       (.I0(\sr_reg[8]_14 ),
        .I1(\sr[4]_i_34 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr_reg[8]_31 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_19 ));
  LUT6 #(
    .INIT(64'hFFFF0000CDC8CDC8)) 
    \iv[5]_i_22 
       (.I0(\iv[9]_i_28 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\tr[28]_i_8_0 ),
        .I3(\iv[15]_i_131_n_0 ),
        .I4(\iv[13]_i_40_n_0 ),
        .I5(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_31 ));
  LUT6 #(
    .INIT(64'hAFA0C0C0AFA0CFCF)) 
    \iv[5]_i_23 
       (.I0(\iv[15]_i_128_n_0 ),
        .I1(\sr_reg[8]_90 ),
        .I2(\iv[9]_i_28 ),
        .I3(\sr_reg[8]_91 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[5]_i_15 ),
        .O(\sr_reg[8]_89 ));
  LUT6 #(
    .INIT(64'hFF33CC00E2E2E2E2)) 
    \iv[5]_i_26 
       (.I0(\iv[13]_i_42_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\tr[21]_i_9_0 ),
        .I4(\tr[21]_i_9_1 ),
        .I5(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_211 ));
  LUT5 #(
    .INIT(32'h5353000F)) 
    \iv[5]_i_29 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\iv[13]_i_49_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\sr_reg[8]_84 ),
        .I4(\iv[0]_i_21 ),
        .O(\sr_reg[8]_83 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[5]_i_30 
       (.I0(\sr_reg[8]_76 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\tr[21]_i_8 ),
        .O(\iv[13]_i_50 ));
  LUT6 #(
    .INIT(64'h0000000002A2AAAA)) 
    \iv[5]_i_8 
       (.I0(\sr_reg[8]_19 ),
        .I1(\sr[4]_i_34 ),
        .I2(\sr[4]_i_91 ),
        .I3(\mul_a_reg[32] ),
        .I4(\sr[5]_i_3_0 ),
        .I5(\iv[5]_i_3 ),
        .O(\sr_reg[8]_18 ));
  LUT3 #(
    .INIT(8'h47)) 
    \iv[6]_i_11 
       (.I0(\mul_a_reg[30] ),
        .I1(\iv[5]_i_7 ),
        .I2(\niho_dsp_a[7] [2]),
        .O(\badr[6]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[6]_i_16 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[6]_i_8 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr_reg[8]_26 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_25 ));
  LUT6 #(
    .INIT(64'h550000035500FF03)) 
    \iv[6]_i_17 
       (.I0(\sr_reg[8]_6 ),
        .I1(\niho_dsp_b[5] ),
        .I2(\sr[4]_i_38 ),
        .I3(\sr[4]_i_38_0 ),
        .I4(\sr[4]_i_91 ),
        .I5(\sr_reg[8]_7 ),
        .O(\sr_reg[8]_4 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \iv[6]_i_18 
       (.I0(\iv[6]_i_28_n_0 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[6]_i_10 ),
        .I4(\sr[6]_i_11_0 ),
        .I5(\sr_reg[8]_74 ),
        .O(\sr_reg[8]_5 ));
  LUT6 #(
    .INIT(64'hFFFF0000CDC8CDC8)) 
    \iv[6]_i_25 
       (.I0(\iv[9]_i_28 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\tr[28]_i_8_0 ),
        .I3(\iv[12]_i_39_n_0 ),
        .I4(\iv[14]_i_50_n_0 ),
        .I5(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_26 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \iv[6]_i_26 
       (.I0(\sr_reg[8]_110 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr[7]_i_30_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[23]_i_7 ),
        .O(\sr_reg[8]_6 ));
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \iv[6]_i_27 
       (.I0(\sr[7]_i_26_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[8]_109 ),
        .I3(\tr[22]_i_9 ),
        .I4(\sr[6]_i_11_0 ),
        .O(\sr_reg[8]_7 ));
  LUT5 #(
    .INIT(32'h5353000F)) 
    \iv[6]_i_28 
       (.I0(\iv[14]_i_55_n_0 ),
        .I1(\iv[14]_i_56_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\sr_reg[8]_77 ),
        .I4(\sr[6]_i_11_0 ),
        .O(\iv[6]_i_28_n_0 ));
  LUT5 #(
    .INIT(32'hB0B0AAA0)) 
    \iv[6]_i_9 
       (.I0(\sr_reg[8]_4 ),
        .I1(\sr_reg[8]_5 ),
        .I2(\iv[6]_i_3 ),
        .I3(sr[8]),
        .I4(\niho_dsp_b[5] ),
        .O(\sr_reg[8]_3 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[7]_i_17 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[7]_i_8 ),
        .I2(\sr[4]_i_91 ),
        .I3(\iv[7]_i_36_n_0 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_38 ));
  LUT5 #(
    .INIT(32'h00044404)) 
    \iv[7]_i_21 
       (.I0(\sr[4]_i_38_0 ),
        .I1(\sr[4]_i_91 ),
        .I2(\iv[8]_i_34 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_51 ),
        .O(\sr_reg[8]_75 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[7]_i_36 
       (.I0(\iv[15]_i_95_n_0 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr_reg[8]_40 ),
        .O(\iv[7]_i_36_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[7]_i_39 
       (.I0(\sr_reg[8]_94 ),
        .I1(\iv[11]_i_47_n_0 ),
        .I2(\sr[6]_i_11_0 ),
        .I3(\tr[23]_i_6 ),
        .I4(\tr[23]_i_6_0 ),
        .I5(\tr[19]_i_6 ),
        .O(\sr_reg[8]_95 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[7]_i_42 
       (.I0(\iv[7]_i_47_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[7]_i_48_n_0 ),
        .O(\sr_reg[8]_93 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[7]_i_47 
       (.I0(\mul_a_reg[21] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[22] ),
        .O(\iv[7]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \iv[7]_i_48 
       (.I0(\mul_a_reg[19] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[20] ),
        .O(\iv[7]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[8]_i_11 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[8]_i_4 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr_reg[8]_30 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_29 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[8]_i_13 
       (.I0(\sr_reg[8]_54 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\sr[4]_i_74 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_53 ),
        .I5(\tr[23]_i_3 ),
        .O(\sr_reg[8]_61 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_25 
       (.I0(\sr_reg[8]_70 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr_reg[8]_40 ),
        .O(\sr_reg[8]_30 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_28 
       (.I0(\sr_reg[8]_97 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[12]_i_47_n_0 ),
        .O(\sr_reg[8]_54 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_30 
       (.I0(\iv[12]_i_48_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[8]_100 ),
        .O(\sr_reg[8]_53 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[8]_i_31 
       (.I0(\sr_reg[8]_54 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\tr[24]_i_9 ),
        .O(\iv[8]_i_38 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \iv[9]_i_11 
       (.I0(\sr_reg[8]_14 ),
        .I1(\iv[9]_i_4 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr_reg[8]_28 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\sr_reg[8]_27 ));
  LUT6 #(
    .INIT(64'h2233223330333000)) 
    \iv[9]_i_13 
       (.I0(\sr_reg[8]_65 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\sr[4]_i_66 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_66 ),
        .I5(\tr[23]_i_3 ),
        .O(\sr_reg[8]_64 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_26 
       (.I0(\iv[9]_i_46_n_0 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr_reg[8]_40 ),
        .O(\sr_reg[8]_28 ));
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \iv[9]_i_27 
       (.I0(\sr_reg[8]_88 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[13]_i_43_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[26]_i_7 ),
        .I5(\tr[26]_i_7_0 ),
        .O(\sr_reg[8]_213 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \iv[9]_i_29 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[8]_84 ),
        .O(\sr_reg[8]_65 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \iv[9]_i_31 
       (.I0(\iv[13]_i_49_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[8]_86 ),
        .O(\sr_reg[8]_66 ));
  LUT5 #(
    .INIT(32'hE2FFE200)) 
    \iv[9]_i_32 
       (.I0(\iv[13]_i_48_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr_reg[6]_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[25]_i_9 ),
        .O(\sr_reg[8]_145 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_45 
       (.I0(\iv[15]_i_134_n_0 ),
        .I1(\iv[15]_i_127_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[15]_i_128_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\sr_reg[8]_90 ),
        .O(\sr_reg[8]_69 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \iv[9]_i_46 
       (.I0(\sr_reg[8]_40 ),
        .I1(\iv[15]_i_131_n_0 ),
        .I2(\iv[9]_i_28 ),
        .I3(\iv[15]_i_132_n_0 ),
        .I4(\tr[28]_i_8_0 ),
        .I5(\iv[15]_i_133_n_0 ),
        .O(\iv[9]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[9]_i_47 
       (.I0(\iv[15]_i_168_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_169_n_0 ),
        .O(\sr_reg[8]_88 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \iv[9]_i_49 
       (.I0(\iv[13]_i_42_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[15]_i_164_n_0 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\iv[9]_i_28_0 ),
        .O(\sr_reg[8]_87 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \iv[9]_i_50 
       (.I0(\sr_reg[6]_1 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[15]_i_141_n_0 ),
        .O(\sr_reg[6]_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[16]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[16] ),
        .O(\sr_reg[8]_121 ));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[17]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[17] ),
        .O(mul_a_i[0]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[18]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[18] ),
        .O(mul_a_i[1]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[19]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[19] ),
        .O(mul_a_i[2]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[20]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[20] ),
        .O(mul_a_i[3]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[21]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[21] ),
        .O(mul_a_i[4]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[22]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[22] ),
        .O(mul_a_i[5]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[23]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[23] ),
        .O(mul_a_i[6]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[24]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[24] ),
        .O(mul_a_i[7]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[25]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[25] ),
        .O(mul_a_i[8]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[26]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[26] ),
        .O(mul_a_i[9]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[27]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[27] ),
        .O(mul_a_i[10]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[28]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[28] ),
        .O(mul_a_i[11]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[29]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[29] ),
        .O(mul_a_i[12]));
  LUT2 #(
    .INIT(4'h8)) 
    \mul_a[30]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[30] ),
        .O(mul_a_i[13]));
  LUT3 #(
    .INIT(8'h80)) 
    \mul_a[31]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(rst_n),
        .O(\sr_reg[8]_219 [0]));
  LUT4 #(
    .INIT(16'h8000)) 
    \mul_a[32]_i_1 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\mul_a_reg[32]_0 ),
        .I3(rst_n),
        .O(\sr_reg[8]_219 [1]));
  LUT2 #(
    .INIT(4'h2)) 
    mul_rslt_i_1
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .O(mul_rslt0));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[0]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[3] [0]),
        .I3(mul_rslt),
        .I4(mul_a[0]),
        .O(niho_dsp_a[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[10]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[11] [2]),
        .I3(mul_rslt),
        .I4(mul_a[10]),
        .O(niho_dsp_a[10]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[11]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[11] [3]),
        .I3(mul_rslt),
        .I4(mul_a[11]),
        .O(niho_dsp_a[11]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[12]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(DI[0]),
        .I3(mul_rslt),
        .I4(mul_a[12]),
        .O(niho_dsp_a[12]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[13]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(DI[1]),
        .I3(mul_rslt),
        .I4(mul_a[13]),
        .O(niho_dsp_a[13]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[14]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(DI[2]),
        .I3(mul_rslt),
        .I4(mul_a[14]),
        .O(niho_dsp_a[14]));
  LUT5 #(
    .INIT(32'h80FF8080)) 
    \niho_dsp_a[15]_INST_0 
       (.I0(sr[8]),
        .I1(mul_rslt),
        .I2(mul_a[15]),
        .I3(\niho_dsp_b[5]_0 ),
        .I4(niho_dsp_a_15_sn_1),
        .O(niho_dsp_a[15]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[1]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[3] [1]),
        .I3(mul_rslt),
        .I4(mul_a[1]),
        .O(niho_dsp_a[1]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[2]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[3] [2]),
        .I3(mul_rslt),
        .I4(mul_a[2]),
        .O(niho_dsp_a[2]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[3]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[3] [3]),
        .I3(mul_rslt),
        .I4(mul_a[3]),
        .O(niho_dsp_a[3]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[4]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[7] [0]),
        .I3(mul_rslt),
        .I4(mul_a[4]),
        .O(niho_dsp_a[4]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[5]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[7] [1]),
        .I3(mul_rslt),
        .I4(mul_a[5]),
        .O(niho_dsp_a[5]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[6]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[7] [2]),
        .I3(mul_rslt),
        .I4(mul_a[6]),
        .O(niho_dsp_a[6]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[7]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[7] [3]),
        .I3(mul_rslt),
        .I4(mul_a[7]),
        .O(niho_dsp_a[7]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[8]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[11] [0]),
        .I3(mul_rslt),
        .I4(mul_a[8]),
        .O(niho_dsp_a[8]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_a[9]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_a[11] [1]),
        .I3(mul_rslt),
        .I4(mul_a[9]),
        .O(niho_dsp_a[9]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[0]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(niho_dsp_b_0_sn_1),
        .I3(mul_rslt),
        .I4(\niho_dsp_b[0]_0 ),
        .O(niho_dsp_b[0]));
  LUT5 #(
    .INIT(32'hBA101010)) 
    \niho_dsp_b[5]_INST_0 
       (.I0(sr[8]),
        .I1(\niho_dsp_b[5]_0 ),
        .I2(\niho_dsp_b[5] ),
        .I3(mul_rslt),
        .I4(\niho_dsp_b[5]_1 ),
        .O(niho_dsp_b[1]));
  LUT6 #(
    .INIT(64'h5955555599995955)) 
    \pc[3]_i_3 
       (.I0(\pc_reg[3]_i_2 ),
        .I1(irq),
        .I2(irq_lev[0]),
        .I3(sr[2]),
        .I4(sr[3]),
        .I5(irq_lev[1]),
        .O(S));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[16]_i_2 
       (.I0(\mul_a_reg[16] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[3] [0]),
        .I4(\remden_reg[16] ),
        .O(\sr_reg[8]_120 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[17]_i_2 
       (.I0(\mul_a_reg[17] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[3] [1]),
        .I4(\remden_reg[17] ),
        .O(\sr_reg[8]_119 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[18]_i_2 
       (.I0(\mul_a_reg[18] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[3] [2]),
        .I4(\remden_reg[18] ),
        .O(\sr_reg[8]_118 ));
  LUT5 #(
    .INIT(32'h30503F5F)) 
    \remden[19]_i_2 
       (.I0(\niho_dsp_a[3] [3]),
        .I1(\mul_a_reg[19] ),
        .I2(\remden_reg[26] ),
        .I3(sr[8]),
        .I4(\remden_reg[19] ),
        .O(\sr_reg[8]_218 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[20]_i_2 
       (.I0(\mul_a_reg[20] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[7] [0]),
        .I4(\remden_reg[20] ),
        .O(\sr_reg[8]_117 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[21]_i_2 
       (.I0(\mul_a_reg[21] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[7] [1]),
        .I4(\remden_reg[21] ),
        .O(\sr_reg[8]_116 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[22]_i_2 
       (.I0(\mul_a_reg[22] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[7] [2]),
        .I4(\remden_reg[22] ),
        .O(\sr_reg[8]_115 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[23]_i_2 
       (.I0(\mul_a_reg[23] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[7] [3]),
        .I4(\remden_reg[23] ),
        .O(\sr_reg[8]_114 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[24]_i_2 
       (.I0(\mul_a_reg[24] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[11] [0]),
        .I4(\remden_reg[24] ),
        .O(\sr_reg[8]_113 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[25]_i_2 
       (.I0(\mul_a_reg[25] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(\niho_dsp_a[11] [1]),
        .I4(\remden_reg[25] ),
        .O(\sr_reg[8]_112 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[26]_i_2 
       (.I0(\mul_a_reg[26] ),
        .I1(\niho_dsp_a[11] [2]),
        .I2(\remden_reg[26] ),
        .I3(sr[8]),
        .I4(\remden_reg[26]_0 ),
        .O(\sr_reg[8]_223 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[27]_i_2 
       (.I0(\mul_a_reg[27] ),
        .I1(\niho_dsp_a[11] [3]),
        .I2(\remden_reg[26] ),
        .I3(sr[8]),
        .I4(\remden_reg[27] ),
        .O(\sr_reg[8]_222 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[28]_i_2 
       (.I0(\mul_a_reg[28] ),
        .I1(DI[0]),
        .I2(\remden_reg[26] ),
        .I3(sr[8]),
        .I4(\remden_reg[28] ),
        .O(\sr_reg[8]_221 ));
  LUT5 #(
    .INIT(32'hBFB38C80)) 
    \remden[29]_i_2 
       (.I0(\mul_a_reg[29] ),
        .I1(\remden_reg[26] ),
        .I2(sr[8]),
        .I3(DI[1]),
        .I4(\remden_reg[29] ),
        .O(\sr_reg[8]_111 ));
  LUT5 #(
    .INIT(32'h50305F3F)) 
    \remden[30]_i_2 
       (.I0(\mul_a_reg[30] ),
        .I1(DI[2]),
        .I2(\remden_reg[26] ),
        .I3(sr[8]),
        .I4(\remden_reg[30] ),
        .O(\sr_reg[8]_220 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \remden[31]_i_2 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(niho_dsp_a_15_sn_1),
        .O(\sr_reg[8]_40 ));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[14]_i_1 
       (.I0(sr[14]),
        .I1(rst_n),
        .I2(\sr_reg[15]_0 ),
        .O(p_0_in__0[14]));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[15]_i_1 
       (.I0(sr[15]),
        .I1(rst_n),
        .I2(\sr_reg[15]_0 ),
        .O(p_0_in__0[15]));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_105 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_46 ),
        .I2(\sr[4]_i_46_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\sr_reg[8]_138 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_137 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_109 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_47 ),
        .I2(\sr[4]_i_47_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\iv[10]_i_44_0 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_136 ));
  LUT4 #(
    .INIT(16'h0002)) 
    \sr[4]_i_11 
       (.I0(\sr[4]_i_28_n_0 ),
        .I1(\sr_reg[6]_4 ),
        .I2(\sr[4]_i_3 ),
        .I3(\sr[4]_i_3_0 ),
        .O(\sr_reg[8]_122 ));
  LUT5 #(
    .INIT(32'hF0F0F0E0)) 
    \sr[4]_i_111 
       (.I0(\tr_reg[23]_i_11_n_5 ),
        .I1(\tr_reg[31]_i_32_n_6 ),
        .I2(sr[8]),
        .I3(\sr_reg[6]_i_6_n_5 ),
        .I4(\tr_reg[23]_i_11_n_7 ),
        .O(\sr[4]_i_111_n_0 ));
  LUT4 #(
    .INIT(16'hFFFE)) 
    \sr[4]_i_112 
       (.I0(\tr_reg[31]_i_13_n_6 ),
        .I1(\tr_reg[31]_i_32_n_4 ),
        .I2(\tr_reg[23]_i_11_n_4 ),
        .I3(\tr_reg[23]_i_11_n_6 ),
        .O(\sr[4]_i_112_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[4]_i_119 
       (.I0(\iv[9]_i_46_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr[4]_i_69_0 ),
        .I4(\iv[0]_i_21 ),
        .I5(\sr_reg[8]_69 ),
        .O(\sr[4]_i_119_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \sr[4]_i_121 
       (.I0(\sr_reg[8]_69 ),
        .I1(\iv[0]_i_21 ),
        .I2(\sr[4]_i_69_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\mul_a_reg[32] ),
        .I5(\sr[5]_i_3_0 ),
        .O(\sr[4]_i_121_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_123 
       (.I0(sr[8]),
        .I1(\sr[4]_i_73 ),
        .I2(\tr[23]_i_3 ),
        .O(\sr_reg[8]_68 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \sr[4]_i_128 
       (.I0(\sr_reg[8]_70 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr[4]_i_74 ),
        .I4(\iv[0]_i_21 ),
        .I5(\sr_reg[8]_71 ),
        .O(\sr[4]_i_128_n_0 ));
  LUT6 #(
    .INIT(64'hFF2E002E00000000)) 
    \sr[4]_i_130 
       (.I0(\sr_reg[8]_71 ),
        .I1(\iv[0]_i_21 ),
        .I2(\sr[4]_i_74 ),
        .I3(\sr[4]_i_91 ),
        .I4(\mul_a_reg[32] ),
        .I5(\sr[5]_i_3_0 ),
        .O(\sr[4]_i_130_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_137 
       (.I0(sr[8]),
        .I1(\sr[4]_i_86 ),
        .I2(\tr[23]_i_3 ),
        .O(\sr_reg[8]_73 ));
  LUT6 #(
    .INIT(64'h1310131313101010)) 
    \sr[4]_i_139 
       (.I0(\sr[4]_i_163_n_0 ),
        .I1(\sr[4]_i_38_0 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr[4]_i_90_0 ),
        .I4(\sr[6]_i_11_0 ),
        .I5(\sr[4]_i_164_n_0 ),
        .O(\sr_reg[8]_48 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_141 
       (.I0(sr[8]),
        .I1(\sr[4]_i_87_0 ),
        .I2(\sr[4]_i_91 ),
        .O(\sr[4]_i_141_n_0 ));
  LUT6 #(
    .INIT(64'hA0AFCFCFA0AFC0C0)) 
    \sr[4]_i_143 
       (.I0(\iv[15]_i_95_n_0 ),
        .I1(\sr_reg[8]_40 ),
        .I2(\sr[4]_i_91 ),
        .I3(\sr[4]_i_90_0 ),
        .I4(\iv[0]_i_21 ),
        .I5(\sr_reg[8]_49 ),
        .O(\sr[4]_i_143_n_0 ));
  LUT6 #(
    .INIT(64'hFF2E002E00000000)) 
    \sr[4]_i_145 
       (.I0(\sr_reg[8]_49 ),
        .I1(\iv[0]_i_21 ),
        .I2(\sr[4]_i_90_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\mul_a_reg[32] ),
        .I5(\sr[5]_i_3_0 ),
        .O(\sr[4]_i_145_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[4]_i_150 
       (.I0(\iv[11]_i_24_n_0 ),
        .I1(\sr[4]_i_91 ),
        .I2(\sr[4]_i_94_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\iv[11]_i_42_n_0 ),
        .O(\sr[4]_i_150_n_0 ));
  LUT6 #(
    .INIT(64'hFFE200E200000000)) 
    \sr[4]_i_152 
       (.I0(\iv[11]_i_42_n_0 ),
        .I1(\iv[0]_i_21 ),
        .I2(\sr[4]_i_94_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\mul_a_reg[32] ),
        .I5(\sr[5]_i_3_0 ),
        .O(\sr[4]_i_152_n_0 ));
  LUT3 #(
    .INIT(8'hBA)) 
    \sr[4]_i_155 
       (.I0(sr[8]),
        .I1(\sr[4]_i_103 ),
        .I2(\tr[23]_i_3 ),
        .O(\sr_reg[8]_72 ));
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \sr[4]_i_163 
       (.I0(\sr[4]_i_169_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr[4]_i_170_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\mul_a_reg[32] ),
        .I5(\sr[4]_i_139_0 ),
        .O(\sr[4]_i_163_n_0 ));
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \sr[4]_i_164 
       (.I0(\sr_reg[8]_93 ),
        .I1(\iv[9]_i_28 ),
        .I2(\badr[18]_INST_0_i_1 ),
        .I3(\tr[28]_i_8_0 ),
        .I4(\iv[15]_i_58 ),
        .O(\sr[4]_i_164_n_0 ));
  LUT6 #(
    .INIT(64'h55510004555DFFF7)) 
    \sr[4]_i_169 
       (.I0(\iv[15]_i_141_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[13]_i_51_n_0 ),
        .O(\sr[4]_i_169_n_0 ));
  LUT6 #(
    .INIT(64'h55510004555DFFF7)) 
    \sr[4]_i_170 
       (.I0(\iv[13]_i_52_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\iv[13]_i_53_n_0 ),
        .O(\sr[4]_i_170_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFF)) 
    \sr[4]_i_28 
       (.I0(\sr[4]_i_48_n_0 ),
        .I1(\sr_reg[6]_i_6_n_4 ),
        .I2(\tr_reg[31]_i_13_n_7 ),
        .I3(O),
        .I4(\sr[4]_i_49_n_0 ),
        .I5(sr[8]),
        .O(\sr[4]_i_28_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \sr[4]_i_36 
       (.I0(\sr_reg[8]_17 ),
        .I1(\sr[4]_i_17 ),
        .O(\iv[10]_i_9 ));
  LUT6 #(
    .INIT(64'hD5DD0000D5DDD5DD)) 
    \sr[4]_i_42 
       (.I0(\sr[4]_i_19 ),
        .I1(\sr[4]_i_87_n_0 ),
        .I2(\sr[4]_i_88_n_0 ),
        .I3(\sr[4]_i_19_0 ),
        .I4(\sr[4]_i_90_n_0 ),
        .I5(\sr[4]_i_19_1 ),
        .O(\sr_reg[8]_2 ));
  LUT5 #(
    .INIT(32'hFFFFF0E0)) 
    \sr[4]_i_48 
       (.I0(\sr_reg[6]_i_6_n_7 ),
        .I1(\tr_reg[31]_i_32_n_7 ),
        .I2(sr[8]),
        .I3(\tr_reg[31]_i_13_n_5 ),
        .I4(\sr[4]_i_111_n_0 ),
        .O(\sr[4]_i_48_n_0 ));
  LUT4 #(
    .INIT(16'hEEEA)) 
    \sr[4]_i_49 
       (.I0(\sr[4]_i_112_n_0 ),
        .I1(sr[8]),
        .I2(\tr_reg[31]_i_32_n_5 ),
        .I3(\alu/art/add/tout [18]),
        .O(\sr[4]_i_49_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_54 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_31 ),
        .I2(\sr[4]_i_31_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\iv[12]_i_49 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_141 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_59 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_33 ),
        .I2(\sr[4]_i_33_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\iv[13]_i_50 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_140 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_64 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_35 ),
        .I2(\sr[4]_i_35_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\iv[10]_i_34 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_139 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_67 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_37_0 ),
        .I2(\sr[4]_i_37_1 ),
        .I3(\sr[4]_i_91 ),
        .I4(\sr_reg[8]_145 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_144 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_69 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_42_0 ),
        .I2(\sr[4]_i_119_n_0 ),
        .I3(\sr_reg[8]_14 ),
        .I4(\sr[4]_i_37 ),
        .I5(\sr[4]_i_121_n_0 ),
        .O(\sr_reg[8]_24 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_75 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_39_0 ),
        .I2(\sr[4]_i_39_1 ),
        .I3(\sr[4]_i_91 ),
        .I4(\iv[8]_i_38 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_142 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_77 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_42_0 ),
        .I2(\sr[4]_i_128_n_0 ),
        .I3(\sr_reg[8]_14 ),
        .I4(\sr[4]_i_39 ),
        .I5(\sr[4]_i_130_n_0 ),
        .O(\sr_reg[8]_22 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_79 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_40_0 ),
        .I2(\iv[14]_i_30_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\sr[4]_i_40_1 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_143 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_81 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_42_0 ),
        .I2(\iv[14]_i_27_n_0 ),
        .I3(\sr_reg[8]_14 ),
        .I4(\sr[4]_i_40 ),
        .I5(\iv[15]_i_54_n_0 ),
        .O(\sr_reg[8]_23 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_84 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_41 ),
        .I2(\sr[4]_i_41_0 ),
        .I3(\sr[4]_i_91 ),
        .I4(\sr_reg[8]_135 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr_reg[8]_134 ));
  LUT6 #(
    .INIT(64'hFF4FFF4FFF5F5555)) 
    \sr[4]_i_87 
       (.I0(\sr[4]_i_42_2 ),
        .I1(\sr_reg[8]_48 ),
        .I2(\sr[4]_i_42_3 ),
        .I3(\sr[4]_i_141_n_0 ),
        .I4(sr[8]),
        .I5(bbus_0[2]),
        .O(\sr[4]_i_87_n_0 ));
  LUT6 #(
    .INIT(64'h4444444455544454)) 
    \sr[4]_i_88 
       (.I0(\sr_reg[8]_79 ),
        .I1(\sr[4]_i_42_4 ),
        .I2(\sr[4]_i_42_5 ),
        .I3(\sr[4]_i_91 ),
        .I4(\sr_reg[8]_95 ),
        .I5(\sr[4]_i_42_6 ),
        .O(\sr[4]_i_88_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_90 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_42_0 ),
        .I2(\sr[4]_i_143_n_0 ),
        .I3(\sr_reg[8]_14 ),
        .I4(\sr[4]_i_42_1 ),
        .I5(\sr[4]_i_145_n_0 ),
        .O(\sr[4]_i_90_n_0 ));
  LUT6 #(
    .INIT(64'h00000000000047FF)) 
    \sr[4]_i_94 
       (.I0(\mul_a_reg[32] ),
        .I1(\sr[4]_i_42_0 ),
        .I2(\sr[4]_i_150_n_0 ),
        .I3(\sr_reg[8]_14 ),
        .I4(\sr[4]_i_43 ),
        .I5(\sr[4]_i_152_n_0 ),
        .O(\sr_reg[8]_15 ));
  LUT6 #(
    .INIT(64'h00000000FFFF0140)) 
    \sr[5]_i_2 
       (.I0(sr[8]),
        .I1(\sr_reg[5]_2 ),
        .I2(\sr_reg[5]_3 ),
        .I3(\alu/asr0 ),
        .I4(\sr[5]_i_7_n_0 ),
        .I5(\sr_reg[6]_4 ),
        .O(\sr_reg[8]_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \sr[5]_i_6 
       (.I0(sr[8]),
        .I1(\mul_a_reg[16] ),
        .I2(niho_dsp_a_15_sn_1),
        .O(\alu/asr0 ));
  LUT5 #(
    .INIT(32'h20020880)) 
    \sr[5]_i_7 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\sr_reg[6]_5 ),
        .I3(\sr[5]_i_2_0 ),
        .I4(O),
        .O(\sr[5]_i_7_n_0 ));
  LUT6 #(
    .INIT(64'hFFFFFFFF1010FF10)) 
    \sr[6]_i_11 
       (.I0(sr[8]),
        .I1(bbus_0[2]),
        .I2(\sr[6]_i_4_0 ),
        .I3(\sr[6]_i_29_n_0 ),
        .I4(\sr[6]_i_4_1 ),
        .I5(\sr[6]_i_4_2 ),
        .O(\sr[6]_i_11_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_15 
       (.I0(sr[8]),
        .I1(\mul_a_reg[19] ),
        .O(\sr[6]_i_15_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_16 
       (.I0(sr[8]),
        .I1(\mul_a_reg[18] ),
        .O(\sr[6]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_17 
       (.I0(sr[8]),
        .I1(\mul_a_reg[17] ),
        .O(\sr[6]_i_17_n_0 ));
  LUT3 #(
    .INIT(8'hF8)) 
    \sr[6]_i_18 
       (.I0(sr[8]),
        .I1(\mul_a_reg[16] ),
        .I2(niho_dsp_a_15_sn_1),
        .O(\sr[6]_i_18_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_19 
       (.I0(sr[8]),
        .I1(\mul_a_reg[19] ),
        .I2(\sr_reg[6]_i_6_0 ),
        .I3(\sr_reg[6]_5 ),
        .O(\sr[6]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_20 
       (.I0(sr[8]),
        .I1(\mul_a_reg[18] ),
        .I2(\sr_reg[6]_i_6_1 ),
        .I3(\sr_reg[6]_5 ),
        .O(\sr[6]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_21 
       (.I0(sr[8]),
        .I1(\mul_a_reg[17] ),
        .I2(\sr_reg[6]_i_6_2 ),
        .I3(\sr_reg[6]_5 ),
        .O(\sr[6]_i_21_n_0 ));
  LUT2 #(
    .INIT(4'h9)) 
    \sr[6]_i_22 
       (.I0(\alu/asr0 ),
        .I1(\sr_reg[5]_2 ),
        .O(\sr[6]_i_22_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \sr[6]_i_23 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .O(\sr[6]_i_23_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \sr[6]_i_24 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\sr_reg[6]_5 ),
        .I3(\sr[5]_i_2_0 ),
        .O(\sr[6]_i_24_n_0 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[6]_i_26 
       (.I0(\sr[6]_i_33_n_0 ),
        .I1(\tr[23]_i_6_0 ),
        .I2(\sr[6]_i_10 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_51 ),
        .O(\sr_reg[8]_106 ));
  LUT6 #(
    .INIT(64'h4444444440444000)) 
    \sr[6]_i_29 
       (.I0(\niho_dsp_b[5] ),
        .I1(sr[8]),
        .I2(\sr_reg[8]_42 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_43 ),
        .I5(\sr[6]_i_11_1 ),
        .O(\sr[6]_i_29_n_0 ));
  LUT6 #(
    .INIT(64'hAAAAAAAAEEEBBBEB)) 
    \sr[6]_i_3 
       (.I0(\sr_reg[8]_12 ),
        .I1(\sr_reg[6]_5 ),
        .I2(\alu/art/add/tout [18]),
        .I3(sr[8]),
        .I4(\alu/art/add/tout [34]),
        .I5(\sr_reg[6]_4 ),
        .O(alu_sr_flag));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[6]_i_33 
       (.I0(\mul_a_reg[22] ),
        .I1(\mul_a_reg[21] ),
        .I2(\tr[28]_i_8_0 ),
        .I3(\mul_a_reg[20] ),
        .I4(niho_dsp_b_0_sn_1),
        .I5(\mul_a_reg[19] ),
        .O(\sr[6]_i_33_n_0 ));
  LUT3 #(
    .INIT(8'hE2)) 
    \sr[6]_i_36 
       (.I0(\sr_reg[8]_104 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[15]_i_136_n_0 ),
        .O(\sr_reg[8]_42 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[6]_i_37 
       (.I0(\sr_reg[8]_105 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[15]_i_138_n_0 ),
        .O(\sr_reg[8]_43 ));
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \sr[6]_i_38 
       (.I0(\iv[15]_i_136_n_0 ),
        .I1(\iv[9]_i_28 ),
        .I2(\sr[6]_i_41_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_43 ),
        .O(\sr_reg[8]_102 ));
  LUT5 #(
    .INIT(32'h0E0E000E)) 
    \sr[6]_i_4 
       (.I0(\sr[6]_i_9_n_0 ),
        .I1(\sr[5]_i_3 ),
        .I2(\sr[6]_i_11_n_0 ),
        .I3(\sr[5]_i_3_0 ),
        .I4(\sr[5]_i_3_1 ),
        .O(\sr_reg[8]_12 ));
  LUT6 #(
    .INIT(64'h50305F3F503F5F3F)) 
    \sr[6]_i_41 
       (.I0(\mul_a_reg[29] ),
        .I1(\mul_a_reg[30] ),
        .I2(\tr[28]_i_8_0 ),
        .I3(niho_dsp_b_0_sn_1),
        .I4(\mul_a_reg[32] ),
        .I5(\sr[6]_i_38_0 ),
        .O(\sr[6]_i_41_n_0 ));
  LUT4 #(
    .INIT(16'h80FF)) 
    \sr[6]_i_9 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\sr[6]_i_4_3 ),
        .I3(\sr_reg[8]_14 ),
        .O(\sr[6]_i_9_n_0 ));
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \sr[7]_i_13 
       (.I0(\sr[7]_i_26_n_0 ),
        .I1(\sr_reg[8]_109 ),
        .I2(\sr[6]_i_11_0 ),
        .I3(\sr_reg[8]_110 ),
        .I4(\iv[9]_i_28 ),
        .I5(\sr[7]_i_30_n_0 ),
        .O(\sr_reg[8]_13 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \sr[7]_i_18 
       (.I0(\sr_reg[8]_74 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr_reg[8]_108 ),
        .O(\iv[14]_i_30_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_26 
       (.I0(\sr[7]_i_45_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\sr[7]_i_46_n_0 ),
        .O(\sr[7]_i_26_n_0 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_27 
       (.I0(\sr[7]_i_47_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\sr[7]_i_48_n_0 ),
        .O(\sr_reg[8]_109 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_28 
       (.I0(\badr[16]_INST_0_i_1 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\sr[7]_i_50_n_0 ),
        .O(\sr_reg[8]_110 ));
  LUT6 #(
    .INIT(64'hAAAEFFFBAAA20008)) 
    \sr[7]_i_30 
       (.I0(\sr[7]_i_51_n_0 ),
        .I1(niho_dsp_b_0_sn_1),
        .I2(\sr_reg[8]_80 ),
        .I3(\sr_reg[8]_79 ),
        .I4(bbus_0[0]),
        .I5(\sr[7]_i_52_n_0 ),
        .O(\sr[7]_i_30_n_0 ));
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \sr[7]_i_39 
       (.I0(sr[8]),
        .I1(\iv[15]_i_96_4 ),
        .I2(\iv[15]_i_96_5 ),
        .I3(\iv[15]_i_96_6 ),
        .I4(\iv[15]_i_96_7 ),
        .I5(\iv[15]_i_96_8 ),
        .O(\sr_reg[8]_80 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_45 
       (.I0(\mul_a_reg[25] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[24] ),
        .O(\sr[7]_i_45_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_46 
       (.I0(\mul_a_reg[27] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[26] ),
        .O(\sr[7]_i_46_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_47 
       (.I0(\mul_a_reg[29] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[28] ),
        .O(\sr[7]_i_47_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_48 
       (.I0(\mul_a_reg[32] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[30] ),
        .O(\sr[7]_i_48_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_49 
       (.I0(\mul_a_reg[17] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[16] ),
        .O(\badr[16]_INST_0_i_1 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_50 
       (.I0(\mul_a_reg[19] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[18] ),
        .O(\sr[7]_i_50_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_51 
       (.I0(\mul_a_reg[21] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[20] ),
        .O(\sr[7]_i_51_n_0 ));
  LUT6 #(
    .INIT(64'h00000001FFFFFFFD)) 
    \sr[7]_i_52 
       (.I0(\mul_a_reg[23] ),
        .I1(\iv[13]_i_45_0 ),
        .I2(\iv[13]_i_45_1 ),
        .I3(\iv[10]_i_44_1 ),
        .I4(\iv[10]_i_44_2 ),
        .I5(\mul_a_reg[22] ),
        .O(\sr[7]_i_52_n_0 ));
  LUT6 #(
    .INIT(64'h0000000E000E000E)) 
    \sr[7]_i_7 
       (.I0(\sr[7]_i_9_n_0 ),
        .I1(\sr[5]_i_3_2 ),
        .I2(\sr[5]_i_3_3 ),
        .I3(\sr[5]_i_3_4 ),
        .I4(\sr_reg[8]_13 ),
        .I5(\sr[5]_i_3_5 ),
        .O(\sr_reg[8]_1 ));
  LUT5 #(
    .INIT(32'h80FFFFFF)) 
    \sr[7]_i_9 
       (.I0(sr[8]),
        .I1(\mul_a_reg[30] ),
        .I2(\sr[6]_i_4_3 ),
        .I3(\niho_dsp_b[5] ),
        .I4(\sr[4]_i_38_0 ),
        .O(\sr[7]_i_9_n_0 ));
  LUT3 #(
    .INIT(8'h80)) 
    \sr[9]_i_1 
       (.I0(sr[9]),
        .I1(rst_n),
        .I2(\sr_reg[15]_0 ),
        .O(p_0_in__0[9]));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[0] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[0]_97 ),
        .Q(sr[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[10] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[10]_0 ),
        .Q(sr[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[11] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[11]_0 ),
        .Q(sr[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[12] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[0]),
        .Q(sr[12]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[13] 
       (.C(clk),
        .CE(\<const1> ),
        .D(D[1]),
        .Q(sr[13]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[14] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_0_in__0[14]),
        .Q(sr[14]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[15] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_0_in__0[15]),
        .Q(sr[15]),
        .R(\<const0> ));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[1] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[1]_9 ),
        .Q(sr[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[2] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[2]_0 ),
        .Q(sr[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[3] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[3]_0 ),
        .Q(sr[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[4] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[4]_2 ),
        .Q(sr[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[5] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[5]_4 ),
        .Q(sr[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[6] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[6]_6 ),
        .Q(sr[6]),
        .R(SR));
  CARRY4 \sr_reg[6]_i_6 
       (.CI(CO),
        .CO({\sr_reg[6]_i_6_n_0 ,\sr_reg[6]_i_6_n_1 ,\sr_reg[6]_i_6_n_2 ,\sr_reg[6]_i_6_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\sr[6]_i_15_n_0 ,\sr[6]_i_16_n_0 ,\sr[6]_i_17_n_0 ,\sr[6]_i_18_n_0 }),
        .O({\sr_reg[6]_i_6_n_4 ,\sr_reg[6]_i_6_n_5 ,\alu/art/add/tout [18],\sr_reg[6]_i_6_n_7 }),
        .S({\sr[6]_i_19_n_0 ,\sr[6]_i_20_n_0 ,\sr[6]_i_21_n_0 ,\sr[6]_i_22_n_0 }));
  CARRY4 \sr_reg[6]_i_7 
       (.CI(\tr_reg[31]_i_13_n_0 ),
        .CO(\alu/art/add/tout [34]),
        .CYINIT(\<const0> ),
        .DI({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_23_n_0 }),
        .S({\<const0> ,\<const0> ,\<const0> ,\sr[6]_i_24_n_0 }));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[7] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[7]_4 ),
        .Q(sr[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[8] 
       (.C(clk),
        .CE(\<const1> ),
        .D(\sr_reg[8]_228 ),
        .Q(sr[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \sr_reg[9] 
       (.C(clk),
        .CE(\<const1> ),
        .D(p_0_in__0[9]),
        .Q(sr[9]),
        .R(\<const0> ));
  LUT5 #(
    .INIT(32'hA65656A6)) 
    \stat[0]_i_17 
       (.I0(\badr[31]_INST_0_i_69 [1]),
        .I1(sr[4]),
        .I2(\badr[31]_INST_0_i_69 [4]),
        .I3(sr[5]),
        .I4(sr[7]),
        .O(\sr_reg[4]_1 ));
  LUT5 #(
    .INIT(32'hFFEEFCFF)) 
    \stat[0]_i_19 
       (.I0(sr[6]),
        .I1(\stat[0]_i_6 [1]),
        .I2(sr[5]),
        .I3(\badr[31]_INST_0_i_69 [4]),
        .I4(\badr[31]_INST_0_i_69 [3]),
        .O(\sr_reg[6]_3 ));
  LUT6 #(
    .INIT(64'h28AA2800820082AA)) 
    \stat[1]_i_4 
       (.I0(\stat_reg[1] ),
        .I1(sr[7]),
        .I2(sr[5]),
        .I3(\badr[31]_INST_0_i_69 [4]),
        .I4(sr[4]),
        .I5(\badr[31]_INST_0_i_69 [1]),
        .O(\sr_reg[7]_2 ));
  LUT6 #(
    .INIT(64'h1200120030FF3030)) 
    \stat[2]_i_10 
       (.I0(sr[7]),
        .I1(\badr[31]_INST_0_i_69 [3]),
        .I2(sr[5]),
        .I3(\badr[31]_INST_0_i_69 [4]),
        .I4(sr[6]),
        .I5(\badr[31]_INST_0_i_69 [2]),
        .O(\stat[2]_i_10_n_0 ));
  LUT6 #(
    .INIT(64'h00000000F7F0F7FC)) 
    \stat[2]_i_7 
       (.I0(sr[7]),
        .I1(\badr[31]_INST_0_i_69 [2]),
        .I2(\badr[31]_INST_0_i_69 [4]),
        .I3(\badr[31]_INST_0_i_69 [3]),
        .I4(sr[4]),
        .I5(\stat[2]_i_10_n_0 ),
        .O(\sr_reg[7]_0 ));
  LUT6 #(
    .INIT(64'h555557F7FFFF57F7)) 
    \tr[16]_i_11 
       (.I0(\sr_reg[8]_14 ),
        .I1(\tr[16]_i_25_n_0 ),
        .I2(\tr[23]_i_3 ),
        .I3(\sr_reg[8]_40 ),
        .I4(\sr[4]_i_42_0 ),
        .I5(\mul_a_reg[32] ),
        .O(\tr[16]_i_11_n_0 ));
  LUT5 #(
    .INIT(32'hAAAABABF)) 
    \tr[16]_i_14 
       (.I0(\sr[4]_i_38_0 ),
        .I1(\sr_reg[8]_53 ),
        .I2(\sr[6]_i_11_0 ),
        .I3(\sr_reg[8]_54 ),
        .I4(\sr[4]_i_91 ),
        .O(\sr_reg[8]_52 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[16]_i_20 
       (.I0(\mul_a_reg[24] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_6 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[16]_i_23 
       (.I0(sr[8]),
        .I1(\sr_reg[6]_i_6_n_7 ),
        .O(\sr_reg[8]_128 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \tr[16]_i_25 
       (.I0(\sr_reg[8]_71 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr_reg[8]_70 ),
        .O(\tr[16]_i_25_n_0 ));
  LUT4 #(
    .INIT(16'h0151)) 
    \tr[16]_i_27 
       (.I0(\tr[23]_i_3 ),
        .I1(\sr_reg[8]_54 ),
        .I2(\sr[6]_i_11_0 ),
        .I3(\sr_reg[8]_53 ),
        .O(\sr_reg[8]_133 ));
  LUT3 #(
    .INIT(8'hB8)) 
    \tr[16]_i_29 
       (.I0(\sr_reg[8]_46 ),
        .I1(\sr[6]_i_11_0 ),
        .I2(\sr_reg[8]_45 ),
        .O(\iv[0]_i_31_0 ));
  LUT5 #(
    .INIT(32'h8A88AAAA)) 
    \tr[16]_i_4 
       (.I0(\sr[4]_i_19_1 ),
        .I1(\iv[15]_i_54_n_0 ),
        .I2(\tr[16]_i_2 ),
        .I3(\tr[16]_i_2_0 ),
        .I4(\tr[16]_i_11_n_0 ),
        .O(\sr_reg[8]_39 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[17]_i_10 
       (.I0(sr[8]),
        .I1(\alu/art/add/tout [18]),
        .O(\sr_reg[8]_131 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[17]_i_14 
       (.I0(\mul_a_reg[25] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_5 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[18]_i_10 
       (.I0(sr[8]),
        .I1(\sr_reg[6]_i_6_n_5 ),
        .O(\sr_reg[8]_123 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[18]_i_14 
       (.I0(\mul_a_reg[26] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_4 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[19]_i_13 
       (.I0(\mul_a_reg[27] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_3 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[19]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\sr_reg[6]_i_6_n_4 ),
        .I2(Q[0]),
        .I3(\tr[19]_i_2 ),
        .I4(\tr[29]_i_2 [0]),
        .I5(\tr[19]_i_2_0 ),
        .O(\quo_reg[19] ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[20]_i_10 
       (.I0(sr[8]),
        .I1(\tr_reg[23]_i_11_n_7 ),
        .O(\sr_reg[8]_124 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[20]_i_13 
       (.I0(\mul_a_reg[28] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_2 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[21]_i_12 
       (.I0(\mul_a_reg[29] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_1 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[21]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[23]_i_11_n_6 ),
        .I2(\tr[29]_i_2 [1]),
        .I3(\tr[19]_i_2_0 ),
        .I4(Q[1]),
        .I5(\tr[19]_i_2 ),
        .O(\rem_reg[21] ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[22]_i_10 
       (.I0(sr[8]),
        .I1(\tr_reg[23]_i_11_n_5 ),
        .O(\sr_reg[8]_125 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[22]_i_15 
       (.I0(\mul_a_reg[30] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[23]_i_13 
       (.I0(\mul_a_reg[32] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_16 
       (.I0(sr[8]),
        .I1(\mul_a_reg[23] ),
        .O(\tr[23]_i_16_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_17 
       (.I0(sr[8]),
        .I1(\mul_a_reg[22] ),
        .O(\tr[23]_i_17_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_18 
       (.I0(sr[8]),
        .I1(\mul_a_reg[21] ),
        .O(\tr[23]_i_18_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[23]_i_19 
       (.I0(sr[8]),
        .I1(\mul_a_reg[20] ),
        .O(\tr[23]_i_19_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_20 
       (.I0(sr[8]),
        .I1(\mul_a_reg[23] ),
        .I2(\tr_reg[23]_i_11_0 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[23]_i_20_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_21 
       (.I0(sr[8]),
        .I1(\mul_a_reg[22] ),
        .I2(\tr_reg[23]_i_11_1 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[23]_i_21_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_22 
       (.I0(sr[8]),
        .I1(\mul_a_reg[21] ),
        .I2(\tr_reg[23]_i_11_2 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[23]_i_22_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[23]_i_23 
       (.I0(sr[8]),
        .I1(\mul_a_reg[20] ),
        .I2(\tr_reg[23]_i_11_3 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[23]_i_23_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[23]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[23]_i_11_n_4 ),
        .I2(Q[2]),
        .I3(\tr[19]_i_2 ),
        .I4(\tr[29]_i_2 [2]),
        .I5(\tr[19]_i_2_0 ),
        .O(\quo_reg[23] ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[23]_i_9 
       (.I0(\iv[7]_i_36_n_0 ),
        .I1(\tr[23]_i_3 ),
        .I2(\tr[28]_i_3 ),
        .O(\sr_reg[8]_11 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[24]_i_11 
       (.I0(sr[8]),
        .I1(\tr_reg[31]_i_32_n_7 ),
        .O(\sr_reg[8]_127 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[24]_i_13 
       (.I0(\mul_a_reg[16] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_13 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[25]_i_11 
       (.I0(sr[8]),
        .I1(\tr_reg[31]_i_32_n_6 ),
        .O(\sr_reg[8]_126 ));
  LUT6 #(
    .INIT(64'hFFFF0000B8FF0000)) 
    \tr[25]_i_17 
       (.I0(\sr_reg[8]_84 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[13]_i_48_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[27]_i_9 ),
        .I5(\tr[23]_i_3 ),
        .O(\sr_reg[8]_225 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[26]_i_10 
       (.I0(sr[8]),
        .I1(\tr_reg[31]_i_32_n_5 ),
        .O(\sr_reg[8]_130 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[26]_i_13 
       (.I0(\mul_a_reg[18] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_12 ));
  LUT6 #(
    .INIT(64'hFFFF0000B8FF0000)) 
    \tr[26]_i_15 
       (.I0(\sr_reg[8]_77 ),
        .I1(\iv[9]_i_28 ),
        .I2(\iv[14]_i_55_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\tr[27]_i_9 ),
        .I5(\tr[23]_i_3 ),
        .O(\sr_reg[8]_224 ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[26]_i_8 
       (.I0(\iv[10]_i_23_n_0 ),
        .I1(\tr[23]_i_3 ),
        .I2(\tr[28]_i_3 ),
        .O(\sr_reg[8]_10 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[27]_i_14 
       (.I0(\mul_a_reg[19] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_11 ));
  LUT3 #(
    .INIT(8'hA8)) 
    \tr[27]_i_16 
       (.I0(\tr[27]_i_9 ),
        .I1(\tr[27]_i_18_n_0 ),
        .I2(\tr[23]_i_3 ),
        .O(\sr_reg[8]_67 ));
  LUT6 #(
    .INIT(64'hEEEEE2EEFFFFFFFF)) 
    \tr[27]_i_18 
       (.I0(\sr_reg[8]_94 ),
        .I1(\iv[9]_i_28 ),
        .I2(niho_dsp_b_0_sn_1),
        .I3(\mul_a_reg[32] ),
        .I4(bbus_0[0]),
        .I5(\sr[6]_i_11_0 ),
        .O(\tr[27]_i_18_n_0 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[27]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[31]_i_32_n_4 ),
        .I2(Q[3]),
        .I3(\tr[19]_i_2 ),
        .I4(\tr[29]_i_2 [3]),
        .I5(\tr[19]_i_2_0 ),
        .O(\quo_reg[27] ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[27]_i_8 
       (.I0(\iv[11]_i_24_n_0 ),
        .I1(\tr[23]_i_3 ),
        .I2(\tr[28]_i_3 ),
        .O(\sr_reg[8]_9 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[28]_i_11 
       (.I0(\mul_a_reg[20] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_10 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[28]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[31]_i_13_n_7 ),
        .I2(\tr[29]_i_2 [4]),
        .I3(\tr[19]_i_2_0 ),
        .I4(Q[4]),
        .I5(\tr[19]_i_2 ),
        .O(\rem_reg[28] ));
  LUT3 #(
    .INIT(8'h0D)) 
    \tr[28]_i_8 
       (.I0(\iv[12]_i_23_n_0 ),
        .I1(\tr[23]_i_3 ),
        .I2(\tr[28]_i_3 ),
        .O(\sr_reg[8]_8 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[29]_i_10 
       (.I0(sr[8]),
        .I1(\sr_reg[6]_4 ),
        .O(\tr[29]_i_10_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[29]_i_12 
       (.I0(\mul_a_reg[21] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_9 ));
  LUT6 #(
    .INIT(64'h88F888F8FFFF88F8)) 
    \tr[29]_i_4 
       (.I0(\tr[29]_i_10_n_0 ),
        .I1(\tr_reg[31]_i_13_n_6 ),
        .I2(\tr[29]_i_2 [5]),
        .I3(\tr[19]_i_2_0 ),
        .I4(Q[5]),
        .I5(\tr[19]_i_2 ),
        .O(\rem_reg[29] ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[30]_i_11 
       (.I0(sr[8]),
        .I1(\tr_reg[31]_i_13_n_5 ),
        .O(\sr_reg[8]_129 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[30]_i_14 
       (.I0(\mul_a_reg[22] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_8 ));
  LUT5 #(
    .INIT(32'hFEFF1000)) 
    \tr[30]_i_16 
       (.I0(\iv[9]_i_28 ),
        .I1(\tr[28]_i_8_0 ),
        .I2(\iv[12]_i_39_n_0 ),
        .I3(\sr[6]_i_11_0 ),
        .I4(\sr_reg[8]_40 ),
        .O(\sr_reg[8]_62 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_33 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .O(\tr[31]_i_33_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_34 
       (.I0(sr[8]),
        .I1(\mul_a_reg[30] ),
        .O(\tr[31]_i_34_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_35 
       (.I0(sr[8]),
        .I1(\mul_a_reg[29] ),
        .O(\tr[31]_i_35_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_36 
       (.I0(sr[8]),
        .I1(\mul_a_reg[28] ),
        .O(\tr[31]_i_36_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_37 
       (.I0(sr[8]),
        .I1(\mul_a_reg[32] ),
        .I2(\sr_reg[6]_5 ),
        .I3(\sr[5]_i_2_0 ),
        .O(\tr[31]_i_37_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_38 
       (.I0(sr[8]),
        .I1(\mul_a_reg[30] ),
        .I2(\tr_reg[31]_i_13_0 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[31]_i_38_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_39 
       (.I0(sr[8]),
        .I1(\mul_a_reg[29] ),
        .I2(\tr_reg[31]_i_13_1 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[31]_i_39_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_40 
       (.I0(sr[8]),
        .I1(\mul_a_reg[28] ),
        .I2(\tr_reg[31]_i_13_2 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[31]_i_40_n_0 ));
  LUT2 #(
    .INIT(4'h2)) 
    \tr[31]_i_43 
       (.I0(\mul_a_reg[23] ),
        .I1(\tr[23]_i_5 ),
        .O(\iv[15]_i_108_7 ));
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFAAEA)) 
    \tr[31]_i_5 
       (.I0(\sr_reg[8]_1 ),
        .I1(sr[8]),
        .I2(O),
        .I3(\sr_reg[6]_4 ),
        .I4(\tr_reg[31] ),
        .I5(\tr_reg[31]_0 ),
        .O(p_2_in));
  LUT6 #(
    .INIT(64'h50AF5FA030CF30CF)) 
    \tr[31]_i_57 
       (.I0(sr[7]),
        .I1(sr[6]),
        .I2(\badr[31]_INST_0_i_69 [3]),
        .I3(\badr[31]_INST_0_i_69 [1]),
        .I4(sr[4]),
        .I5(\badr[31]_INST_0_i_69 [2]),
        .O(\sr_reg[7]_3 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_62 
       (.I0(sr[8]),
        .I1(\mul_a_reg[27] ),
        .O(\tr[31]_i_62_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_63 
       (.I0(sr[8]),
        .I1(\mul_a_reg[26] ),
        .O(\tr[31]_i_63_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_64 
       (.I0(sr[8]),
        .I1(\mul_a_reg[25] ),
        .O(\tr[31]_i_64_n_0 ));
  LUT2 #(
    .INIT(4'h8)) 
    \tr[31]_i_65 
       (.I0(sr[8]),
        .I1(\mul_a_reg[24] ),
        .O(\tr[31]_i_65_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_66 
       (.I0(sr[8]),
        .I1(\mul_a_reg[27] ),
        .I2(\tr_reg[31]_i_32_0 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[31]_i_66_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_67 
       (.I0(sr[8]),
        .I1(\mul_a_reg[26] ),
        .I2(\tr_reg[31]_i_32_1 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[31]_i_67_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_68 
       (.I0(sr[8]),
        .I1(\mul_a_reg[25] ),
        .I2(\tr_reg[31]_i_32_2 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[31]_i_68_n_0 ));
  LUT4 #(
    .INIT(16'h8228)) 
    \tr[31]_i_69 
       (.I0(sr[8]),
        .I1(\mul_a_reg[24] ),
        .I2(\tr_reg[31]_i_32_3 ),
        .I3(\sr_reg[6]_5 ),
        .O(\tr[31]_i_69_n_0 ));
  CARRY4 \tr_reg[23]_i_11 
       (.CI(\sr_reg[6]_i_6_n_0 ),
        .CO({\tr_reg[23]_i_11_n_0 ,\tr_reg[23]_i_11_n_1 ,\tr_reg[23]_i_11_n_2 ,\tr_reg[23]_i_11_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\tr[23]_i_16_n_0 ,\tr[23]_i_17_n_0 ,\tr[23]_i_18_n_0 ,\tr[23]_i_19_n_0 }),
        .O({\tr_reg[23]_i_11_n_4 ,\tr_reg[23]_i_11_n_5 ,\tr_reg[23]_i_11_n_6 ,\tr_reg[23]_i_11_n_7 }),
        .S({\tr[23]_i_20_n_0 ,\tr[23]_i_21_n_0 ,\tr[23]_i_22_n_0 ,\tr[23]_i_23_n_0 }));
  CARRY4 \tr_reg[31]_i_13 
       (.CI(\tr_reg[31]_i_32_n_0 ),
        .CO({\tr_reg[31]_i_13_n_0 ,\tr_reg[31]_i_13_n_1 ,\tr_reg[31]_i_13_n_2 ,\tr_reg[31]_i_13_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\tr[31]_i_33_n_0 ,\tr[31]_i_34_n_0 ,\tr[31]_i_35_n_0 ,\tr[31]_i_36_n_0 }),
        .O({O,\tr_reg[31]_i_13_n_5 ,\tr_reg[31]_i_13_n_6 ,\tr_reg[31]_i_13_n_7 }),
        .S({\tr[31]_i_37_n_0 ,\tr[31]_i_38_n_0 ,\tr[31]_i_39_n_0 ,\tr[31]_i_40_n_0 }));
  CARRY4 \tr_reg[31]_i_32 
       (.CI(\tr_reg[23]_i_11_n_0 ),
        .CO({\tr_reg[31]_i_32_n_0 ,\tr_reg[31]_i_32_n_1 ,\tr_reg[31]_i_32_n_2 ,\tr_reg[31]_i_32_n_3 }),
        .CYINIT(\<const0> ),
        .DI({\tr[31]_i_62_n_0 ,\tr[31]_i_63_n_0 ,\tr[31]_i_64_n_0 ,\tr[31]_i_65_n_0 }),
        .O({\tr_reg[31]_i_32_n_4 ,\tr_reg[31]_i_32_n_5 ,\tr_reg[31]_i_32_n_6 ,\tr_reg[31]_i_32_n_7 }),
        .S({\tr[31]_i_66_n_0 ,\tr[31]_i_67_n_0 ,\tr[31]_i_68_n_0 ,\tr[31]_i_69_n_0 }));
endmodule

module niho_rgf_treg
   (.\tr_reg[31]_0 ({tr[31],tr[30],tr[29],tr[28],tr[27],tr[26],tr[25],tr[24],tr[23],tr[22],tr[21],tr[20],tr[19],tr[18],tr[17],tr[16],tr[15],tr[14],tr[13],tr[12],tr[11],tr[10],tr[9],tr[8],tr[7],tr[6],tr[5],tr[4],tr[3],tr[2],tr[1],tr[0]}),
    SR,
    \tr_reg[0]_0 ,
    cbus,
    clk);
  input [0:0]SR;
  input [0:0]\tr_reg[0]_0 ;
  input [31:0]cbus;
  input clk;
     output [31:0]tr;

  wire [0:0]SR;
  wire [31:0]cbus;
  wire clk;
  (* DONT_TOUCH *) wire [31:0]tr;
  wire [0:0]\tr_reg[0]_0 ;

  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[0] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[0]),
        .Q(tr[0]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[10] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[10]),
        .Q(tr[10]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[11] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[11]),
        .Q(tr[11]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[12] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[12]),
        .Q(tr[12]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[13] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[13]),
        .Q(tr[13]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[14] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[14]),
        .Q(tr[14]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[15] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[15]),
        .Q(tr[15]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[16] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[16]),
        .Q(tr[16]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[17] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[17]),
        .Q(tr[17]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[18] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[18]),
        .Q(tr[18]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[19] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[19]),
        .Q(tr[19]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[1] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[1]),
        .Q(tr[1]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[20] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[20]),
        .Q(tr[20]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[21] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[21]),
        .Q(tr[21]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[22] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[22]),
        .Q(tr[22]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[23] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[23]),
        .Q(tr[23]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[24] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[24]),
        .Q(tr[24]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[25] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[25]),
        .Q(tr[25]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[26] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[26]),
        .Q(tr[26]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[27] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[27]),
        .Q(tr[27]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[28] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[28]),
        .Q(tr[28]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[29] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[29]),
        .Q(tr[29]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[2] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[2]),
        .Q(tr[2]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[30] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[30]),
        .Q(tr[30]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[31] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[31]),
        .Q(tr[31]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[3] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[3]),
        .Q(tr[3]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[4] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[4]),
        .Q(tr[4]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[5] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[5]),
        .Q(tr[5]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[6] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[6]),
        .Q(tr[6]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[7] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[7]),
        .Q(tr[7]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[8] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[8]),
        .Q(tr[8]),
        .R(SR));
  (* DONT_TOUCH *) 
  (* KEEP = "yes" *) 
  FDRE \tr_reg[9] 
       (.C(clk),
        .CE(\tr_reg[0]_0 ),
        .D(cbus[9]),
        .Q(tr[9]),
        .R(SR));
endmodule

(* STRUCTURAL_NETLIST = "yes" *)
module nihonium
   (clk,
    rst_n,
    brdy,
    irq,
    cpuid,
    irq_lev,
    irq_vec,
    fdat,
    bdatr,
    fadr,
    bcmd,
    badr,
    bdatw,
    crdy,
    cbus_i,
    ccmd,
    abus_o,
    bbus_o,
    niho_dsp_c,
    niho_dsp_a,
    niho_dsp_b);
//
//	Nihonium 16/32 bit CPU core
//		(c) 2022	1YEN Toru
//
//
//	2023/09/30	ver.1.16
//		change instruction fetch latency: 0 => 1
//		corresponding to Xilinx Vivado
//
//	2023/07/08	ver.1.14
//		instruction: adcz, sbbz, cmbz
//
//	2023/05/20	ver.1.12
//		instruction: divur, divsr, mulur, mulsr
//
//	2023/03/18	ver.1.10
//		instruction: jall, rtnl, pushcl, popcl
//
//	2023/03/11	ver.1.08
//		corresponding to 32 bit memory bus
//
//	2023/02/11	ver.1.06
//		instruction: fdown
//
//	2022/10/22	ver.1.04
//		corresponding to interrupt vector / level
//
//	2022/06/04	ver.1.02
//		instruction: csft, csfti
//
//	2022/04/09	ver.1.00
//		external 16 bit / internal 32 bit CPU
//		32 bit divider from divc32 ver.1.00
//		extended instructions:
//			link, unlk, brn, ldli, cendl, pushl, popl,
//			exsgl, exzrl, ldl, stl, ldlsp, stlsp
//
// ================================
//
//	2022/02/19	ver.1.10
//		corresponding to extended address
//		badrx output
//
//	2021/07/31	ver.1.08
//		sr bit field: cpu id for dual core edition
//
//	2021/07/10	ver.1.06
//		hcmp: half compare
//		cmb: compare with borrow
//		adc, sbb: condition of z flag changed
//
//	2021/06/12	ver.1.04
//		half precision fpu instruction:
//			hadd, hsub, hmul, hdiv, hneg, hhalf, huint, hfrac, hmvsg, hsat
//
//	2021/05/22	ver.1.02
//		mul/div instruction: mulu, muls, divu, divs, divlu, divls, divlq, divlr
//		co-processor control bit to sr
//		co-processor I/F
//
//	2021/05/01	ver.1.00
//		interrupt related instruction: pause, rti
//		sr bit operation instruction: sesrl, sesrh, clsrl, clsrh
//		sp relative instruction: ldwsp, stwsp
//		control register iv and tr
//		interrupt enable ie bit in sr
//
//	2021/04/10	ver.0.92
//		alu: smaller barrel shift unit
//
//	2021/03/06	ver.0.90
//
  input clk;
  input rst_n;
  input brdy;
  input irq;
  input [1:0]cpuid;
  input [1:0]irq_lev;
  input [5:0]irq_vec;
  input [15:0]fdat;
  input [31:0]bdatr;
  output [15:0]fadr;
  output [3:0]bcmd;
  output [31:0]badr;
  output [31:0]bdatw;
  input crdy;
  input [31:0]cbus_i;
  output [4:0]ccmd;
  output [31:0]abus_o;
  output [31:0]bbus_o;
  input [65:0]niho_dsp_c;
  output [32:0]niho_dsp_a;
  output [32:0]niho_dsp_b;

  wire [31:0]abus_0;
  wire [31:0]abus_o;
  wire [7:0]abus_sel_0;
  wire [5:0]abus_sel_cr;
  wire alu_n_136;
  wire alu_n_137;
  wire alu_n_138;
  wire alu_n_139;
  wire alu_n_140;
  wire alu_n_141;
  wire alu_n_142;
  wire alu_n_143;
  wire alu_n_144;
  wire alu_n_145;
  wire alu_n_146;
  wire alu_n_147;
  wire alu_n_148;
  wire alu_n_149;
  wire alu_n_150;
  wire alu_n_151;
  wire alu_n_152;
  wire alu_n_153;
  wire alu_n_154;
  wire alu_n_155;
  wire alu_n_156;
  wire alu_n_157;
  wire alu_n_158;
  wire alu_n_159;
  wire alu_n_160;
  wire alu_n_161;
  wire alu_n_162;
  wire alu_n_163;
  wire alu_n_164;
  wire alu_n_165;
  wire alu_n_166;
  wire alu_n_167;
  wire alu_n_4;
  wire alu_n_5;
  wire alu_n_6;
  wire alu_n_69;
  wire alu_n_70;
  wire alu_n_71;
  wire alu_n_72;
  wire alu_n_73;
  wire alu_n_74;
  wire alu_n_75;
  wire alu_n_76;
  wire alu_n_77;
  wire alu_n_78;
  wire alu_n_79;
  wire alu_n_80;
  wire alu_n_81;
  wire alu_n_82;
  wire alu_n_83;
  wire alu_n_84;
  wire alu_n_85;
  wire alu_n_86;
  wire [2:2]alu_sr_flag;
  wire [31:0]badr;
  wire [30:0]bbus_0;
  wire [31:0]bbus_o;
  wire [7:0]bbus_sel_0;
  wire [5:0]bbus_sel_cr;
  wire [5:0]bbus_sr;
  wire [3:0]bcmd;
  wire [31:0]bdatr;
  wire [31:0]bdatw;
  wire brdy;
  wire [31:0]cbus;
  wire [15:0]cbus_bk2;
  wire [31:0]cbus_i;
  wire [5:5]cbus_sel_0;
  wire [4:2]cbus_sel_cr;
  wire [4:0]ccmd;
  wire clk;
  wire [1:0]cpuid;
  wire crdy;
  (* DONT_TOUCH *) wire ctl_fetch;
  wire ctl_n_0;
  wire ctl_n_10;
  wire ctl_n_11;
  wire ctl_n_12;
  wire ctl_n_13;
  wire ctl_n_14;
  wire ctl_n_15;
  wire ctl_n_16;
  wire ctl_n_17;
  wire ctl_n_18;
  wire ctl_n_19;
  wire ctl_n_20;
  wire ctl_n_21;
  wire ctl_n_22;
  wire ctl_n_23;
  wire ctl_n_24;
  wire ctl_n_25;
  wire ctl_n_26;
  wire ctl_n_27;
  wire ctl_n_4;
  wire ctl_n_5;
  wire ctl_n_6;
  wire ctl_n_7;
  wire ctl_n_8;
  wire ctl_n_9;
  wire [1:1]ctl_selb_0;
  wire [1:0]ctl_selb_rn;
  wire ctl_sp_dec;
  wire ctl_sp_id4;
  wire ctl_sp_inc;
  wire \div/dctl/dctl_sign ;
  wire \div/dctl/dctl_sign_f ;
  wire [30:0]\div/quo ;
  wire [30:0]\div/rem ;
  wire div_crdy;
  wire [15:0]fadr;
  wire [15:0]fch_ir;
  wire fch_irq_req;
  wire fch_n_10;
  wire fch_n_11;
  wire fch_n_119;
  wire fch_n_12;
  wire fch_n_120;
  wire fch_n_121;
  wire fch_n_122;
  wire fch_n_123;
  wire fch_n_124;
  wire fch_n_125;
  wire fch_n_126;
  wire fch_n_127;
  wire fch_n_128;
  wire fch_n_129;
  wire fch_n_130;
  wire fch_n_131;
  wire fch_n_132;
  wire fch_n_133;
  wire fch_n_134;
  wire fch_n_135;
  wire fch_n_136;
  wire fch_n_137;
  wire fch_n_138;
  wire fch_n_139;
  wire fch_n_140;
  wire fch_n_141;
  wire fch_n_142;
  wire fch_n_143;
  wire fch_n_144;
  wire fch_n_145;
  wire fch_n_146;
  wire fch_n_147;
  wire fch_n_148;
  wire fch_n_149;
  wire fch_n_150;
  wire fch_n_151;
  wire fch_n_152;
  wire fch_n_153;
  wire fch_n_154;
  wire fch_n_155;
  wire fch_n_156;
  wire fch_n_157;
  wire fch_n_158;
  wire fch_n_159;
  wire fch_n_160;
  wire fch_n_161;
  wire fch_n_162;
  wire fch_n_163;
  wire fch_n_164;
  wire fch_n_165;
  wire fch_n_166;
  wire fch_n_167;
  wire fch_n_168;
  wire fch_n_169;
  wire fch_n_170;
  wire fch_n_171;
  wire fch_n_172;
  wire fch_n_173;
  wire fch_n_174;
  wire fch_n_175;
  wire fch_n_176;
  wire fch_n_177;
  wire fch_n_178;
  wire fch_n_179;
  wire fch_n_180;
  wire fch_n_181;
  wire fch_n_182;
  wire fch_n_183;
  wire fch_n_184;
  wire fch_n_185;
  wire fch_n_186;
  wire fch_n_187;
  wire fch_n_188;
  wire fch_n_189;
  wire fch_n_190;
  wire fch_n_191;
  wire fch_n_192;
  wire fch_n_193;
  wire fch_n_194;
  wire fch_n_195;
  wire fch_n_196;
  wire fch_n_197;
  wire fch_n_198;
  wire fch_n_199;
  wire fch_n_200;
  wire fch_n_201;
  wire fch_n_202;
  wire fch_n_203;
  wire fch_n_204;
  wire fch_n_205;
  wire fch_n_206;
  wire fch_n_207;
  wire fch_n_208;
  wire fch_n_209;
  wire fch_n_212;
  wire fch_n_213;
  wire fch_n_214;
  wire fch_n_215;
  wire fch_n_216;
  wire fch_n_217;
  wire fch_n_218;
  wire fch_n_219;
  wire fch_n_220;
  wire fch_n_221;
  wire fch_n_223;
  wire fch_n_224;
  wire fch_n_258;
  wire fch_n_261;
  wire fch_n_262;
  wire fch_n_263;
  wire fch_n_265;
  wire fch_n_266;
  wire fch_n_272;
  wire fch_n_275;
  wire fch_n_276;
  wire fch_n_277;
  wire fch_n_280;
  wire fch_n_283;
  wire fch_n_315;
  wire fch_n_316;
  wire fch_n_317;
  wire fch_n_318;
  wire fch_n_319;
  wire fch_n_320;
  wire fch_n_321;
  wire fch_n_322;
  wire fch_n_323;
  wire fch_n_324;
  wire fch_n_325;
  wire fch_n_326;
  wire fch_n_327;
  wire fch_n_328;
  wire fch_n_329;
  wire fch_n_330;
  wire fch_n_331;
  wire fch_n_332;
  wire fch_n_333;
  wire fch_n_334;
  wire fch_n_335;
  wire fch_n_336;
  wire fch_n_341;
  wire fch_n_342;
  wire fch_n_343;
  wire fch_n_344;
  wire fch_n_345;
  wire fch_n_346;
  wire fch_n_347;
  wire fch_n_348;
  wire fch_n_349;
  wire fch_n_350;
  wire fch_n_351;
  wire fch_n_352;
  wire fch_n_353;
  wire fch_n_354;
  wire fch_n_355;
  wire fch_n_356;
  wire fch_n_357;
  wire fch_n_358;
  wire fch_n_359;
  wire fch_n_360;
  wire fch_n_361;
  wire fch_n_362;
  wire fch_n_363;
  wire fch_n_364;
  wire fch_n_365;
  wire fch_n_366;
  wire fch_n_367;
  wire fch_n_368;
  wire fch_n_369;
  wire fch_n_370;
  wire fch_n_371;
  wire fch_n_372;
  wire fch_n_373;
  wire fch_n_374;
  wire fch_n_375;
  wire fch_n_376;
  wire fch_n_377;
  wire fch_n_378;
  wire fch_n_379;
  wire fch_n_38;
  wire fch_n_380;
  wire fch_n_381;
  wire fch_n_382;
  wire fch_n_383;
  wire fch_n_384;
  wire fch_n_385;
  wire fch_n_386;
  wire fch_n_387;
  wire fch_n_388;
  wire fch_n_389;
  wire fch_n_39;
  wire fch_n_390;
  wire fch_n_391;
  wire fch_n_392;
  wire fch_n_393;
  wire fch_n_394;
  wire fch_n_395;
  wire fch_n_396;
  wire fch_n_397;
  wire fch_n_398;
  wire fch_n_399;
  wire fch_n_40;
  wire fch_n_41;
  wire fch_n_42;
  wire fch_n_43;
  wire fch_n_44;
  wire fch_n_446;
  wire fch_n_447;
  wire fch_n_448;
  wire fch_n_449;
  wire fch_n_45;
  wire fch_n_450;
  wire fch_n_451;
  wire fch_n_452;
  wire fch_n_453;
  wire fch_n_454;
  wire fch_n_455;
  wire fch_n_456;
  wire fch_n_457;
  wire fch_n_458;
  wire fch_n_459;
  wire fch_n_460;
  wire fch_n_461;
  wire fch_n_462;
  wire fch_n_495;
  wire fch_n_496;
  wire fch_n_497;
  wire fch_n_498;
  wire fch_n_499;
  wire fch_n_500;
  wire fch_n_501;
  wire fch_n_502;
  wire fch_n_503;
  wire fch_n_504;
  wire fch_n_505;
  wire fch_n_506;
  wire fch_n_507;
  wire fch_n_508;
  wire fch_n_509;
  wire fch_n_510;
  wire fch_n_511;
  wire fch_n_512;
  wire fch_n_513;
  wire fch_n_514;
  wire fch_n_540;
  wire fch_n_541;
  wire fch_n_542;
  wire fch_n_543;
  wire fch_n_56;
  wire fch_n_57;
  wire fch_n_58;
  wire fch_n_59;
  wire fch_n_60;
  wire fch_n_61;
  wire fch_n_62;
  wire fch_n_63;
  wire fch_n_64;
  wire fch_n_65;
  wire fch_n_66;
  wire fch_n_67;
  wire fch_n_68;
  wire fch_n_69;
  wire fch_n_70;
  wire fch_n_71;
  wire fch_n_72;
  wire fch_n_73;
  wire fch_n_74;
  wire fch_n_75;
  wire fch_n_76;
  wire fch_n_77;
  wire fch_n_78;
  wire fch_n_79;
  wire fch_n_80;
  wire fch_n_85;
  wire fch_n_86;
  wire fch_n_87;
  wire fch_n_88;
  wire fch_n_89;
  wire [15:0]fch_pc;
  wire [15:0]fdat;
  wire irq;
  wire [1:0]irq_lev;
  wire [5:0]irq_vec;
  wire [15:1]\ivec/p_0_in ;
  wire mem_n_0;
  wire mem_n_1;
  wire mem_n_17;
  wire mem_n_18;
  wire mem_n_19;
  wire mem_n_2;
  wire mem_n_20;
  wire mem_n_21;
  wire mem_n_22;
  wire mem_n_23;
  wire mem_n_24;
  wire mem_n_25;
  wire mem_n_26;
  wire mem_n_27;
  wire mem_n_28;
  wire mem_n_29;
  wire mem_n_3;
  wire mem_n_30;
  wire mem_n_31;
  wire mem_n_32;
  wire mem_n_33;
  wire mem_n_4;
  wire mem_n_5;
  wire mem_n_6;
  wire [32:0]\mul/mul_a ;
  wire \mul/mul_b ;
  wire \mul/mul_rslt ;
  wire \mul/mul_rslt0 ;
  wire [15:0]\mul/mulh ;
  wire [30:17]mul_a_i;
  wire [32:0]niho_dsp_a;
  wire [32:0]niho_dsp_b;
  wire [65:0]niho_dsp_c;
  wire p_0_in;
  wire [31:19]p_2_in;
  wire [15:0]\pcnt/p_1_in ;
  wire [2:0]read_cyc;
  wire rgf_iv_ve;
  wire rgf_n_100;
  wire rgf_n_101;
  wire rgf_n_102;
  wire rgf_n_103;
  wire rgf_n_104;
  wire rgf_n_105;
  wire rgf_n_106;
  wire rgf_n_107;
  wire rgf_n_108;
  wire rgf_n_109;
  wire rgf_n_110;
  wire rgf_n_111;
  wire rgf_n_112;
  wire rgf_n_113;
  wire rgf_n_114;
  wire rgf_n_115;
  wire rgf_n_116;
  wire rgf_n_117;
  wire rgf_n_118;
  wire rgf_n_119;
  wire rgf_n_120;
  wire rgf_n_121;
  wire rgf_n_122;
  wire rgf_n_123;
  wire rgf_n_124;
  wire rgf_n_125;
  wire rgf_n_126;
  wire rgf_n_127;
  wire rgf_n_128;
  wire rgf_n_129;
  wire rgf_n_130;
  wire rgf_n_131;
  wire rgf_n_132;
  wire rgf_n_133;
  wire rgf_n_134;
  wire rgf_n_135;
  wire rgf_n_136;
  wire rgf_n_137;
  wire rgf_n_138;
  wire rgf_n_139;
  wire rgf_n_14;
  wire rgf_n_140;
  wire rgf_n_141;
  wire rgf_n_142;
  wire rgf_n_143;
  wire rgf_n_144;
  wire rgf_n_145;
  wire rgf_n_146;
  wire rgf_n_147;
  wire rgf_n_149;
  wire rgf_n_15;
  wire rgf_n_150;
  wire rgf_n_151;
  wire rgf_n_152;
  wire rgf_n_153;
  wire rgf_n_154;
  wire rgf_n_155;
  wire rgf_n_156;
  wire rgf_n_157;
  wire rgf_n_158;
  wire rgf_n_159;
  wire rgf_n_16;
  wire rgf_n_160;
  wire rgf_n_161;
  wire rgf_n_162;
  wire rgf_n_163;
  wire rgf_n_164;
  wire rgf_n_165;
  wire rgf_n_166;
  wire rgf_n_167;
  wire rgf_n_168;
  wire rgf_n_169;
  wire rgf_n_17;
  wire rgf_n_170;
  wire rgf_n_171;
  wire rgf_n_172;
  wire rgf_n_173;
  wire rgf_n_174;
  wire rgf_n_175;
  wire rgf_n_176;
  wire rgf_n_177;
  wire rgf_n_178;
  wire rgf_n_179;
  wire rgf_n_18;
  wire rgf_n_180;
  wire rgf_n_181;
  wire rgf_n_182;
  wire rgf_n_183;
  wire rgf_n_184;
  wire rgf_n_185;
  wire rgf_n_186;
  wire rgf_n_187;
  wire rgf_n_188;
  wire rgf_n_189;
  wire rgf_n_19;
  wire rgf_n_190;
  wire rgf_n_191;
  wire rgf_n_192;
  wire rgf_n_193;
  wire rgf_n_194;
  wire rgf_n_195;
  wire rgf_n_196;
  wire rgf_n_197;
  wire rgf_n_198;
  wire rgf_n_199;
  wire rgf_n_20;
  wire rgf_n_200;
  wire rgf_n_201;
  wire rgf_n_202;
  wire rgf_n_203;
  wire rgf_n_204;
  wire rgf_n_205;
  wire rgf_n_206;
  wire rgf_n_207;
  wire rgf_n_208;
  wire rgf_n_209;
  wire rgf_n_21;
  wire rgf_n_210;
  wire rgf_n_211;
  wire rgf_n_212;
  wire rgf_n_213;
  wire rgf_n_214;
  wire rgf_n_215;
  wire rgf_n_216;
  wire rgf_n_217;
  wire rgf_n_218;
  wire rgf_n_219;
  wire rgf_n_22;
  wire rgf_n_220;
  wire rgf_n_221;
  wire rgf_n_222;
  wire rgf_n_223;
  wire rgf_n_224;
  wire rgf_n_225;
  wire rgf_n_226;
  wire rgf_n_227;
  wire rgf_n_228;
  wire rgf_n_229;
  wire rgf_n_23;
  wire rgf_n_230;
  wire rgf_n_231;
  wire rgf_n_232;
  wire rgf_n_233;
  wire rgf_n_234;
  wire rgf_n_235;
  wire rgf_n_236;
  wire rgf_n_237;
  wire rgf_n_238;
  wire rgf_n_239;
  wire rgf_n_24;
  wire rgf_n_240;
  wire rgf_n_241;
  wire rgf_n_242;
  wire rgf_n_243;
  wire rgf_n_244;
  wire rgf_n_245;
  wire rgf_n_246;
  wire rgf_n_247;
  wire rgf_n_248;
  wire rgf_n_249;
  wire rgf_n_25;
  wire rgf_n_250;
  wire rgf_n_251;
  wire rgf_n_252;
  wire rgf_n_253;
  wire rgf_n_254;
  wire rgf_n_255;
  wire rgf_n_256;
  wire rgf_n_257;
  wire rgf_n_258;
  wire rgf_n_259;
  wire rgf_n_26;
  wire rgf_n_260;
  wire rgf_n_261;
  wire rgf_n_262;
  wire rgf_n_27;
  wire rgf_n_28;
  wire rgf_n_29;
  wire rgf_n_296;
  wire rgf_n_297;
  wire rgf_n_298;
  wire rgf_n_299;
  wire rgf_n_30;
  wire rgf_n_300;
  wire rgf_n_301;
  wire rgf_n_302;
  wire rgf_n_303;
  wire rgf_n_304;
  wire rgf_n_305;
  wire rgf_n_306;
  wire rgf_n_307;
  wire rgf_n_308;
  wire rgf_n_309;
  wire rgf_n_31;
  wire rgf_n_310;
  wire rgf_n_311;
  wire rgf_n_312;
  wire rgf_n_313;
  wire rgf_n_314;
  wire rgf_n_315;
  wire rgf_n_316;
  wire rgf_n_317;
  wire rgf_n_318;
  wire rgf_n_319;
  wire rgf_n_32;
  wire rgf_n_33;
  wire rgf_n_334;
  wire rgf_n_335;
  wire rgf_n_336;
  wire rgf_n_337;
  wire rgf_n_338;
  wire rgf_n_339;
  wire rgf_n_34;
  wire rgf_n_340;
  wire rgf_n_341;
  wire rgf_n_342;
  wire rgf_n_343;
  wire rgf_n_344;
  wire rgf_n_345;
  wire rgf_n_346;
  wire rgf_n_347;
  wire rgf_n_348;
  wire rgf_n_35;
  wire rgf_n_350;
  wire rgf_n_351;
  wire rgf_n_352;
  wire rgf_n_353;
  wire rgf_n_354;
  wire rgf_n_355;
  wire rgf_n_356;
  wire rgf_n_357;
  wire rgf_n_358;
  wire rgf_n_359;
  wire rgf_n_36;
  wire rgf_n_360;
  wire rgf_n_361;
  wire rgf_n_362;
  wire rgf_n_363;
  wire rgf_n_364;
  wire rgf_n_365;
  wire rgf_n_366;
  wire rgf_n_367;
  wire rgf_n_368;
  wire rgf_n_369;
  wire rgf_n_37;
  wire rgf_n_370;
  wire rgf_n_371;
  wire rgf_n_38;
  wire rgf_n_39;
  wire rgf_n_40;
  wire rgf_n_41;
  wire rgf_n_42;
  wire rgf_n_43;
  wire rgf_n_437;
  wire rgf_n_438;
  wire rgf_n_439;
  wire rgf_n_44;
  wire rgf_n_440;
  wire rgf_n_441;
  wire rgf_n_442;
  wire rgf_n_443;
  wire rgf_n_444;
  wire rgf_n_445;
  wire rgf_n_446;
  wire rgf_n_449;
  wire rgf_n_45;
  wire rgf_n_450;
  wire rgf_n_451;
  wire rgf_n_452;
  wire rgf_n_453;
  wire rgf_n_454;
  wire rgf_n_455;
  wire rgf_n_456;
  wire rgf_n_457;
  wire rgf_n_458;
  wire rgf_n_459;
  wire rgf_n_46;
  wire rgf_n_460;
  wire rgf_n_461;
  wire rgf_n_462;
  wire rgf_n_463;
  wire rgf_n_464;
  wire rgf_n_465;
  wire rgf_n_466;
  wire rgf_n_467;
  wire rgf_n_468;
  wire rgf_n_469;
  wire rgf_n_47;
  wire rgf_n_470;
  wire rgf_n_471;
  wire rgf_n_474;
  wire rgf_n_475;
  wire rgf_n_476;
  wire rgf_n_477;
  wire rgf_n_479;
  wire rgf_n_48;
  wire rgf_n_49;
  wire rgf_n_50;
  wire rgf_n_528;
  wire rgf_n_529;
  wire rgf_n_530;
  wire rgf_n_531;
  wire rgf_n_532;
  wire rgf_n_533;
  wire rgf_n_534;
  wire rgf_n_535;
  wire rgf_n_536;
  wire rgf_n_537;
  wire rgf_n_538;
  wire rgf_n_539;
  wire rgf_n_540;
  wire rgf_n_541;
  wire rgf_n_542;
  wire rgf_n_543;
  wire rgf_n_544;
  wire rgf_n_545;
  wire rgf_n_546;
  wire rgf_n_547;
  wire rgf_n_548;
  wire rgf_n_549;
  wire rgf_n_550;
  wire rgf_n_551;
  wire rgf_n_552;
  wire rgf_n_553;
  wire rgf_n_554;
  wire rgf_n_555;
  wire rgf_n_556;
  wire rgf_n_557;
  wire rgf_n_558;
  wire rgf_n_559;
  wire rgf_n_560;
  wire rgf_n_561;
  wire rgf_n_562;
  wire rgf_n_563;
  wire rgf_n_564;
  wire rgf_n_565;
  wire rgf_n_566;
  wire rgf_n_567;
  wire rgf_n_568;
  wire rgf_n_569;
  wire rgf_n_570;
  wire rgf_n_571;
  wire rgf_n_572;
  wire rgf_n_573;
  wire rgf_n_574;
  wire rgf_n_575;
  wire rgf_n_576;
  wire rgf_n_577;
  wire rgf_n_578;
  wire rgf_n_579;
  wire rgf_n_58;
  wire rgf_n_580;
  wire rgf_n_581;
  wire rgf_n_582;
  wire rgf_n_583;
  wire rgf_n_584;
  wire rgf_n_585;
  wire rgf_n_586;
  wire rgf_n_587;
  wire rgf_n_59;
  wire rgf_n_60;
  wire rgf_n_95;
  wire rgf_n_96;
  wire rgf_n_97;
  wire rgf_n_98;
  wire rgf_n_99;
  wire rgf_sr_dr;
  wire [3:0]rgf_sr_flag;
  wire [1:0]rgf_sr_ie;
  wire rgf_sr_ml;
  wire rgf_sr_nh;
  wire [15:0]rgf_tr;
  wire rst_n;
  wire [0:0]\sptr/p_0_in ;
  wire [1:0]sr_bank;
  wire [13:12]\sreg/p_0_in ;
  wire [13:12]\sreg/p_0_in__0 ;
  wire [2:0]stat;
  wire [1:0]stat_nx;
  wire [31:16]\treg/p_0_in ;

  niho_alu alu
       (.D({rgf_n_462,rgf_n_463}),
        .Q(\div/quo ),
        .abus_0(abus_0[15:0]),
        .bbus_0(bbus_0),
        .\bcmd[2]_INST_0_i_1 (fch_n_261),
        .clk(clk),
        .crdy(crdy),
        .crdy_0(alu_n_85),
        .dctl_sign(\div/dctl/dctl_sign ),
        .dctl_sign_f(\div/dctl/dctl_sign_f ),
        .\dctl_stat_reg[2] (fch_n_221),
        .div_crdy(div_crdy),
        .div_crdy_reg(alu_n_4),
        .div_crdy_reg_0(alu_n_84),
        .div_crdy_reg_1(alu_n_86),
        .\dso_reg[19] (fch_n_208),
        .\dso_reg[19]_0 (fch_n_207),
        .\dso_reg[19]_1 (fch_n_206),
        .\dso_reg[19]_2 (fch_n_205),
        .\dso_reg[23] (fch_n_204),
        .\dso_reg[23]_0 (fch_n_203),
        .\dso_reg[23]_1 (fch_n_202),
        .\dso_reg[23]_2 (fch_n_201),
        .\dso_reg[27] (fch_n_200),
        .\dso_reg[27]_0 (fch_n_258),
        .\dso_reg[27]_1 (fch_n_199),
        .\dso_reg[27]_2 (fch_n_198),
        .\dso_reg[31] (fch_n_197),
        .\dso_reg[31]_0 (fch_n_196),
        .\dso_reg[31]_1 (fch_n_195),
        .\dso_reg[31]_2 (fch_n_121),
        .mul_a(\mul/mul_a ),
        .mul_a_i(mul_a_i),
        .\mul_a_reg[16] (rgf_n_347),
        .mul_b(\mul/mul_b ),
        .\mul_b_reg[0] (alu_n_167),
        .\mul_b_reg[0]_0 (fch_n_461),
        .\mul_b_reg[10] (alu_n_158),
        .\mul_b_reg[11] (alu_n_157),
        .\mul_b_reg[12] (alu_n_156),
        .\mul_b_reg[13] (alu_n_155),
        .\mul_b_reg[14] (alu_n_154),
        .\mul_b_reg[15] (alu_n_153),
        .\mul_b_reg[16] (alu_n_152),
        .\mul_b_reg[17] (alu_n_151),
        .\mul_b_reg[18] (alu_n_150),
        .\mul_b_reg[19] (alu_n_149),
        .\mul_b_reg[1] (alu_n_166),
        .\mul_b_reg[20] (alu_n_148),
        .\mul_b_reg[21] (alu_n_147),
        .\mul_b_reg[22] (alu_n_146),
        .\mul_b_reg[23] (alu_n_145),
        .\mul_b_reg[24] (alu_n_144),
        .\mul_b_reg[25] (alu_n_143),
        .\mul_b_reg[26] (alu_n_142),
        .\mul_b_reg[27] (alu_n_141),
        .\mul_b_reg[28] (alu_n_140),
        .\mul_b_reg[29] (alu_n_139),
        .\mul_b_reg[2] (alu_n_165),
        .\mul_b_reg[30] (alu_n_138),
        .\mul_b_reg[32] ({alu_n_136,alu_n_137}),
        .\mul_b_reg[32]_0 ({fch_n_332,fch_n_333}),
        .\mul_b_reg[3] (alu_n_164),
        .\mul_b_reg[5] (alu_n_163),
        .\mul_b_reg[6] (alu_n_162),
        .\mul_b_reg[7] (alu_n_161),
        .\mul_b_reg[8] (alu_n_160),
        .\mul_b_reg[9] (alu_n_159),
        .mul_rslt(\mul/mul_rslt ),
        .mul_rslt0(\mul/mul_rslt0 ),
        .mul_rslt_reg(alu_n_6),
        .mulh(\mul/mulh ),
        .\mulh_reg[0] (fch_n_460),
        .\niho_dsp_a[32]_INST_0_i_12 (stat[1]),
        .niho_dsp_b(niho_dsp_b[4]),
        .\niho_dsp_b[4] (fch_n_209),
        .\niho_dsp_b[4]_0 (fch_n_143),
        .niho_dsp_c(niho_dsp_c[31:16]),
        .\niho_dsp_c[31] (alu_n_5),
        .out(fch_ir[7]),
        .p_0_in(p_0_in),
        .\rem_reg[30] (\div/rem ),
        .\remden_reg[12] (alu_n_82),
        .\remden_reg[13] (alu_n_69),
        .\remden_reg[14] (alu_n_83),
        .\remden_reg[15] (alu_n_70),
        .\remden_reg[16] (alu_n_81),
        .\remden_reg[16]_0 (rgf_n_317),
        .\remden_reg[17] (alu_n_80),
        .\remden_reg[17]_0 (rgf_n_314),
        .\remden_reg[18] (alu_n_79),
        .\remden_reg[18]_0 (rgf_n_313),
        .\remden_reg[19] (alu_n_78),
        .\remden_reg[19]_0 (rgf_n_461),
        .\remden_reg[20] (alu_n_77),
        .\remden_reg[20]_0 (rgf_n_311),
        .\remden_reg[21] (alu_n_76),
        .\remden_reg[21]_0 (rgf_n_309),
        .\remden_reg[22] (alu_n_71),
        .\remden_reg[22]_0 (rgf_n_308),
        .\remden_reg[23] (alu_n_72),
        .\remden_reg[23]_0 (rgf_n_306),
        .\remden_reg[24] (alu_n_73),
        .\remden_reg[24]_0 (rgf_n_304),
        .\remden_reg[25] (alu_n_75),
        .\remden_reg[25]_0 (rgf_n_302),
        .\remden_reg[26] (alu_n_74),
        .\remden_reg[26]_0 (rgf_n_470),
        .\remden_reg[27] (rgf_n_469),
        .\remden_reg[28] (rgf_n_466),
        .\remden_reg[29] (rgf_n_297),
        .\remden_reg[30] (rgf_n_464),
        .\remden_reg[31] (rgf_n_177),
        .rgf_sr_nh(rgf_sr_nh),
        .rst_n(rst_n),
        .\tr[31]_i_5 (fch_n_215),
        .\tr[31]_i_5_0 (fch_n_214));
  niho_fsm ctl
       (.D({fch_n_272,stat_nx}),
        .Q(stat),
        .\bcmd[2] (fch_n_266),
        .\bcmd[2]_0 (alu_n_84),
        .clk(clk),
        .ctl_fetch_fl_reg(fch_n_283),
        .out({fch_ir[15:10],fch_ir[6],fch_ir[3],fch_ir[0]}),
        .p_0_in(p_0_in),
        .rgf_sr_flag(rgf_sr_flag[3:1]),
        .\sr_reg[7] (ctl_n_4),
        .\stat[2]_i_2_0 (fch_n_280),
        .\stat_reg[0]_0 (ctl_n_6),
        .\stat_reg[0]_1 (ctl_n_9),
        .\stat_reg[0]_2 (ctl_n_10),
        .\stat_reg[0]_3 (ctl_n_12),
        .\stat_reg[0]_4 (ctl_n_14),
        .\stat_reg[0]_5 (ctl_n_19),
        .\stat_reg[0]_6 (ctl_n_22),
        .\stat_reg[1]_0 (ctl_n_5),
        .\stat_reg[1]_1 (ctl_n_7),
        .\stat_reg[1]_10 (ctl_n_26),
        .\stat_reg[1]_11 (ctl_n_27),
        .\stat_reg[1]_2 (ctl_n_8),
        .\stat_reg[1]_3 (ctl_n_11),
        .\stat_reg[1]_4 (ctl_n_15),
        .\stat_reg[1]_5 (ctl_n_17),
        .\stat_reg[1]_6 (ctl_n_18),
        .\stat_reg[1]_7 (ctl_n_20),
        .\stat_reg[1]_8 (ctl_n_21),
        .\stat_reg[1]_9 (ctl_n_24),
        .\stat_reg[2]_0 (ctl_n_0),
        .\stat_reg[2]_1 (ctl_n_13),
        .\stat_reg[2]_2 (ctl_n_16),
        .\stat_reg[2]_3 (ctl_n_23),
        .\stat_reg[2]_4 (ctl_n_25));
  niho_fch fch
       (.D(\sreg/p_0_in__0 ),
        .E(fch_n_373),
        .O(rgf_n_45),
        .Q({\div/quo [30],\div/quo [26:24],\div/quo [22],\div/quo [20],\div/quo [18:0]}),
        .S({fch_n_501,fch_n_502,fch_n_503,fch_n_504}),
        .abus_0(abus_0),
        .abus_sel_0(abus_sel_0),
        .abus_sel_cr({abus_sel_cr[5],abus_sel_cr[2:0]}),
        .alu_sr_flag(alu_sr_flag),
        .badr(badr),
        .\badr[0]_INST_0_i_1 (fch_n_194),
        .\badr[2]_INST_0_i_1 (fch_n_193),
        .\badr[31]_INST_0_i_1 ({\treg/p_0_in ,rgf_tr}),
        .\badr[31]_INST_0_i_36_0 (rgf_n_439),
        .\badr[5]_INST_0_i_1 (fch_n_192),
        .\badr[6]_INST_0_i_1 (fch_n_191),
        .bbus_0({bbus_0[30:6],bbus_0[4:1]}),
        .bbus_o({bbus_o[31:6],bbus_o[4:1]}),
        .\bbus_o[16]_0 (rgf_n_568),
        .\bbus_o[17]_0 (rgf_n_567),
        .\bbus_o[18]_0 (rgf_n_566),
        .\bbus_o[19]_0 (rgf_n_565),
        .\bbus_o[20]_0 (rgf_n_564),
        .\bbus_o[21]_0 (rgf_n_563),
        .\bbus_o[22]_0 (rgf_n_562),
        .\bbus_o[23]_0 (rgf_n_561),
        .\bbus_o[24]_0 (rgf_n_560),
        .\bbus_o[25]_0 (rgf_n_559),
        .\bbus_o[26]_0 (rgf_n_558),
        .\bbus_o[27]_0 (rgf_n_557),
        .\bbus_o[28]_0 (rgf_n_556),
        .\bbus_o[29]_0 (rgf_n_555),
        .\bbus_o[30] (rgf_n_570),
        .\bbus_o[30]_0 (rgf_n_554),
        .bbus_o_16_sp_1(rgf_n_584),
        .bbus_o_17_sp_1(rgf_n_583),
        .bbus_o_18_sp_1(rgf_n_582),
        .bbus_o_19_sp_1(rgf_n_581),
        .bbus_o_20_sp_1(rgf_n_580),
        .bbus_o_21_sp_1(rgf_n_579),
        .bbus_o_22_sp_1(rgf_n_578),
        .bbus_o_23_sp_1(rgf_n_577),
        .bbus_o_24_sp_1(rgf_n_576),
        .bbus_o_25_sp_1(rgf_n_575),
        .bbus_o_26_sp_1(rgf_n_574),
        .bbus_o_27_sp_1(rgf_n_573),
        .bbus_o_28_sp_1(rgf_n_572),
        .bbus_o_29_sp_1(rgf_n_571),
        .bbus_sel_0(bbus_sel_0),
        .bbus_sel_cr(bbus_sel_cr),
        .bbus_sr({bbus_sr[5],bbus_sr[0]}),
        .\bcmd[0] (ctl_n_25),
        .\bcmd[2] (ctl_n_8),
        .\bcmd[3] (ctl_n_9),
        .bdatr({bdatr[30],bdatr[26:24],bdatr[22],bdatr[20],bdatr[18:8]}),
        .bdatw(bdatw),
        .\bdatw[10]_INST_0_i_1_0 (fch_n_189),
        .\bdatw[11]_INST_0_i_1_0 ({fch_n_512,fch_n_513,fch_n_514}),
        .\bdatw[11]_INST_0_i_2_0 ({fch_n_505,fch_n_506,fch_n_507,fch_n_508}),
        .\bdatw[12]_INST_0_i_1_0 (fch_n_159),
        .\bdatw[12]_INST_0_i_1_1 (fch_n_179),
        .\bdatw[12]_INST_0_i_1_2 (fch_n_182),
        .\bdatw[15]_INST_0_i_1_0 ({fch_n_509,fch_n_510,fch_n_511}),
        .\bdatw[31]_INST_0_i_7_0 (rgf_n_455),
        .\bdatw[31]_INST_0_i_7_1 (ctl_n_12),
        .\bdatw[5] ({bbus_0[5],bbus_0[0]}),
        .\bdatw[8]_INST_0_i_1 (fch_n_190),
        .brdy(brdy),
        .brdy_0(fch_n_280),
        .brdy_1(fch_n_462),
        .cbus({cbus[30],cbus[26:24],cbus[22],cbus[20],cbus[18:0]}),
        .cbus_i({cbus_i[30],cbus_i[26:24],cbus_i[22],cbus_i[20],cbus_i[18:0]}),
        .\cbus_i[30] ({fch_n_56,fch_n_57,fch_n_58,fch_n_59,fch_n_60,fch_n_61,fch_n_62,fch_n_63,fch_n_64,fch_n_65,fch_n_66,fch_n_67,fch_n_68,fch_n_69,fch_n_70,fch_n_71,fch_n_72,fch_n_73,fch_n_74,fch_n_75,fch_n_76,fch_n_77,fch_n_78,fch_n_79,fch_n_80}),
        .cbus_sel_0(cbus_sel_0),
        .ccmd(ccmd[3:0]),
        .\ccmd[0]_INST_0_i_4_0 (ctl_n_17),
        .\ccmd[1]_INST_0_i_1_0 (ctl_n_24),
        .\ccmd[2]_INST_0_i_2_0 (ctl_n_0),
        .\ccmd[2]_INST_0_i_2_1 (ctl_n_21),
        .ccmd_2_sp_1(ctl_n_26),
        .clk(clk),
        .cpuid(cpuid),
        .crdy(crdy),
        .ctl_fetch_fl_reg_0(ctl_fetch),
        .ctl_fetch_fl_reg_1(ctl_n_6),
        .ctl_fetch_fl_reg_2(alu_n_84),
        .ctl_fetch_inferred_i_11_0(rgf_n_446),
        .ctl_fetch_inferred_i_21_0(ctl_n_11),
        .ctl_fetch_inferred_i_29_0(rgf_n_437),
        .ctl_fetch_inferred_i_5_0(rgf_n_441),
        .ctl_fetch_inferred_i_6_0(rgf_n_457),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .ctl_sp_dec(ctl_sp_dec),
        .ctl_sp_id4(ctl_sp_id4),
        .ctl_sp_inc(ctl_sp_inc),
        .dctl_sign(\div/dctl/dctl_sign ),
        .dctl_sign_f(\div/dctl/dctl_sign_f ),
        .div_crdy(div_crdy),
        .div_crdy_reg(fch_n_214),
        .div_crdy_reg_0(fch_n_215),
        .div_crdy_reg_1(fch_n_283),
        .\eir_fl_reg[31]_0 (rgf_n_456),
        .\eir_fl_reg[31]_1 (ctl_n_13),
        .\fch_irq_lev[1]_i_2_0 (ctl_n_14),
        .fch_irq_req(fch_irq_req),
        .fch_pc(fch_pc),
        .fdat(fdat),
        .in0(ctl_fetch),
        .irq(irq),
        .irq_lev(irq_lev),
        .irq_vec(irq_vec),
        .\iv[0]_i_21 (rgf_n_146),
        .\iv[0]_i_21_0 (rgf_n_239),
        .\iv[0]_i_27_0 (fch_n_152),
        .\iv[0]_i_9 (rgf_n_230),
        .\iv[10]_i_21 (fch_n_166),
        .\iv[10]_i_2_0 (rgf_n_118),
        .\iv[10]_i_2_1 (rgf_n_192),
        .\iv[10]_i_34 (fch_n_185),
        .\iv[10]_i_5 (rgf_n_120),
        .\iv[10]_i_6_0 (rgf_n_222),
        .\iv[11]_i_3_0 ({rgf_n_359,rgf_n_360,rgf_n_361,rgf_n_362}),
        .\iv[11]_i_7_0 (rgf_n_459),
        .\iv[11]_i_7_1 (rgf_n_221),
        .\iv[11]_i_7_2 (rgf_n_249),
        .\iv[12]_i_10 (fch_n_135),
        .\iv[12]_i_22_0 (fch_n_164),
        .\iv[12]_i_2_0 (rgf_n_190),
        .\iv[12]_i_34 (fch_n_186),
        .\iv[12]_i_4_0 (rgf_n_155),
        .\iv[12]_i_4_1 (rgf_n_174),
        .\iv[12]_i_6_0 (rgf_n_217),
        .\iv[13]_i_23 (fch_n_162),
        .\iv[13]_i_2_0 (rgf_n_189),
        .\iv[13]_i_5 (rgf_n_114),
        .\iv[13]_i_6_0 (rgf_n_475),
        .\iv[13]_i_6_1 (rgf_n_218),
        .\iv[13]_i_8_0 (rgf_n_60),
        .\iv[14]_i_2_0 (rgf_n_130),
        .\iv[14]_i_2_1 (rgf_n_129),
        .\iv[14]_i_7_0 (rgf_n_219),
        .\iv[14]_i_7_1 (rgf_n_460),
        .\iv[14]_i_7_2 (rgf_n_241),
        .\iv[15]_i_103 (fch_n_188),
        .\iv[15]_i_122_0 (ctl_n_19),
        .\iv[15]_i_13_0 (ctl_n_7),
        .\iv[15]_i_19_0 (fch_n_136),
        .\iv[15]_i_19_1 (fch_n_219),
        .\iv[15]_i_22 (rgf_n_152),
        .\iv[15]_i_22_0 (rgf_n_198),
        .\iv[15]_i_28_0 (rgf_n_307),
        .\iv[15]_i_38_0 (ctl_n_18),
        .\iv[15]_i_9_0 ({rgf_n_47,rgf_n_48,rgf_n_49,rgf_n_50}),
        .\iv[1]_i_21 (rgf_n_193),
        .\iv[1]_i_21_0 (rgf_n_458),
        .\iv[1]_i_21_1 (rgf_n_248),
        .\iv[3]_i_16 (fch_n_134),
        .\iv[3]_i_21 (rgf_n_191),
        .\iv[3]_i_2_0 (rgf_n_468),
        .\iv[3]_i_2_1 ({rgf_n_355,rgf_n_356,rgf_n_357,rgf_n_358}),
        .\iv[3]_i_8_0 (rgf_n_176),
        .\iv[4]_i_8 (rgf_n_257),
        .\iv[4]_i_8_0 (rgf_n_231),
        .\iv[5]_i_8 (rgf_n_234),
        .\iv[5]_i_8_0 (rgf_n_247),
        .\iv[6]_i_10_0 (rgf_n_197),
        .\iv[6]_i_22 (rgf_n_186),
        .\iv[6]_i_2_0 (rgf_n_465),
        .\iv[6]_i_3_0 (rgf_n_136),
        .\iv[6]_i_3_1 (rgf_n_196),
        .\iv[6]_i_8_0 (rgf_n_101),
        .\iv[6]_i_8_1 (rgf_n_167),
        .\iv[7]_i_10 (rgf_n_102),
        .\iv[7]_i_10_0 (rgf_n_254),
        .\iv[7]_i_11_0 (rgf_n_250),
        .\iv[7]_i_11_1 (rgf_n_187),
        .\iv[7]_i_2_0 ({rgf_n_351,rgf_n_352,rgf_n_353,rgf_n_354}),
        .\iv[8]_i_2_0 (rgf_n_169),
        .\iv[8]_i_34_0 (fch_n_153),
        .\iv[8]_i_35 (fch_n_500),
        .\iv[8]_i_4_0 (rgf_n_170),
        .\iv[8]_i_7_0 (rgf_n_182),
        .\iv[8]_i_7_1 (rgf_n_252),
        .\iv[9]_i_35 (fch_n_155),
        .\iv[9]_i_7_0 (rgf_n_181),
        .\iv_reg[0] (ctl_n_16),
        .\iv_reg[0]_0 (ctl_n_20),
        .\iv_reg[0]_1 (ctl_n_10),
        .\mul_a_reg[15] ({\ivec/p_0_in ,rgf_iv_ve}),
        .mul_b(\mul/mul_b ),
        .\mul_b_reg[10] (rgf_n_532),
        .\mul_b_reg[10]_0 (rgf_n_545),
        .\mul_b_reg[11] (rgf_n_531),
        .\mul_b_reg[11]_0 (rgf_n_544),
        .\mul_b_reg[12] (rgf_n_530),
        .\mul_b_reg[12]_0 (rgf_n_543),
        .\mul_b_reg[13] (rgf_n_529),
        .\mul_b_reg[13]_0 (rgf_n_542),
        .\mul_b_reg[14] (rgf_n_528),
        .\mul_b_reg[14]_0 (rgf_n_541),
        .\mul_b_reg[15] (rgf_n_479),
        .\mul_b_reg[15]_0 (rgf_n_540),
        .\mul_b_reg[15]_1 (rgf_n_440),
        .\mul_b_reg[1] (rgf_n_539),
        .\mul_b_reg[1]_0 (rgf_n_552),
        .\mul_b_reg[1]_1 (rgf_n_585),
        .\mul_b_reg[2] (rgf_n_538),
        .\mul_b_reg[2]_0 (rgf_n_551),
        .\mul_b_reg[2]_1 (rgf_n_586),
        .\mul_b_reg[31] (rgf_n_569),
        .\mul_b_reg[31]_0 (rgf_n_553),
        .\mul_b_reg[3] (rgf_n_537),
        .\mul_b_reg[3]_0 (rgf_n_550),
        .\mul_b_reg[3]_1 (rgf_n_587),
        .\mul_b_reg[4] (rgf_n_261),
        .\mul_b_reg[4]_0 (rgf_n_260),
        .\mul_b_reg[4]_1 (rgf_n_259),
        .\mul_b_reg[6] (rgf_n_536),
        .\mul_b_reg[6]_0 (rgf_n_549),
        .\mul_b_reg[7] (rgf_n_535),
        .\mul_b_reg[7]_0 (rgf_n_548),
        .\mul_b_reg[8] (rgf_n_534),
        .\mul_b_reg[8]_0 (rgf_n_547),
        .\mul_b_reg[9] (rgf_n_533),
        .\mul_b_reg[9]_0 (rgf_n_546),
        .mul_rslt(\mul/mul_rslt ),
        .mulh(\mul/mulh ),
        .\niho_dsp_a[15]_INST_0_i_2_0 (fch_n_127),
        .\niho_dsp_a[32]_INST_0_i_5_0 (fch_n_129),
        .\niho_dsp_a[32]_INST_0_i_5_1 (fch_n_130),
        .\niho_dsp_a[32]_INST_0_i_5_2 (fch_n_209),
        .\niho_dsp_a[32]_INST_0_i_5_3 (fch_n_212),
        .\niho_dsp_a[32]_INST_0_i_5_4 (fch_n_217),
        .\niho_dsp_a[32]_INST_0_i_6_0 (ctl_n_27),
        .\niho_dsp_a[32]_INST_0_i_7_0 (fch_n_133),
        .\niho_dsp_a[32]_INST_0_i_9_0 (alu_n_86),
        .niho_dsp_b({niho_dsp_b[32:6],niho_dsp_b[3:1]}),
        .\niho_dsp_b[30] (alu_n_138),
        .\niho_dsp_b[32] ({alu_n_136,alu_n_137}),
        .niho_dsp_b_10_sp_1(alu_n_158),
        .niho_dsp_b_11_sp_1(alu_n_157),
        .niho_dsp_b_12_sp_1(alu_n_156),
        .niho_dsp_b_13_sp_1(alu_n_155),
        .niho_dsp_b_14_sp_1(alu_n_154),
        .niho_dsp_b_15_sp_1(alu_n_153),
        .niho_dsp_b_16_sp_1(alu_n_152),
        .niho_dsp_b_17_sp_1(alu_n_151),
        .niho_dsp_b_18_sp_1(alu_n_150),
        .niho_dsp_b_19_sp_1(alu_n_149),
        .niho_dsp_b_1_sp_1(alu_n_166),
        .niho_dsp_b_20_sp_1(alu_n_148),
        .niho_dsp_b_21_sp_1(alu_n_147),
        .niho_dsp_b_22_sp_1(alu_n_146),
        .niho_dsp_b_23_sp_1(alu_n_145),
        .niho_dsp_b_24_sp_1(alu_n_144),
        .niho_dsp_b_25_sp_1(alu_n_143),
        .niho_dsp_b_26_sp_1(alu_n_142),
        .niho_dsp_b_27_sp_1(alu_n_141),
        .niho_dsp_b_28_sp_1(alu_n_140),
        .niho_dsp_b_29_sp_1(alu_n_139),
        .niho_dsp_b_2_sp_1(alu_n_165),
        .niho_dsp_b_3_sp_1(alu_n_164),
        .niho_dsp_b_6_sp_1(alu_n_162),
        .niho_dsp_b_7_sp_1(alu_n_161),
        .niho_dsp_b_8_sp_1(alu_n_160),
        .niho_dsp_b_9_sp_1(alu_n_159),
        .niho_dsp_c({niho_dsp_c[30],niho_dsp_c[26:24],niho_dsp_c[22],niho_dsp_c[20],niho_dsp_c[18:0]}),
        .out({fch_ir[15:10],fch_ir[7:6],fch_ir[3],fch_ir[0]}),
        .p_0_in(p_0_in),
        .\pc_reg[15] (\pcnt/p_1_in ),
        .read_cyc(read_cyc),
        .rgf_pc(fadr),
        .rst_n(rst_n),
        .rst_n_0({fch_n_332,fch_n_333}),
        .rst_n_1(fch_n_460),
        .rst_n_2(fch_n_461),
        .rst_n_fl_reg_0(fch_n_121),
        .rst_n_fl_reg_1(fch_n_195),
        .rst_n_fl_reg_10(fch_n_204),
        .rst_n_fl_reg_11(fch_n_205),
        .rst_n_fl_reg_12(fch_n_206),
        .rst_n_fl_reg_13(fch_n_207),
        .rst_n_fl_reg_14(fch_n_208),
        .rst_n_fl_reg_15(fch_n_224),
        .rst_n_fl_reg_16(fch_n_258),
        .rst_n_fl_reg_17(fch_n_261),
        .rst_n_fl_reg_18(fch_n_262),
        .rst_n_fl_reg_19(fch_n_265),
        .rst_n_fl_reg_2(fch_n_196),
        .rst_n_fl_reg_20(fch_n_266),
        .rst_n_fl_reg_21(fch_n_275),
        .rst_n_fl_reg_22(fch_n_276),
        .rst_n_fl_reg_23(fch_n_277),
        .rst_n_fl_reg_3(fch_n_197),
        .rst_n_fl_reg_4(fch_n_198),
        .rst_n_fl_reg_5(fch_n_199),
        .rst_n_fl_reg_6(fch_n_200),
        .rst_n_fl_reg_7(fch_n_201),
        .rst_n_fl_reg_8(fch_n_202),
        .rst_n_fl_reg_9(fch_n_203),
        .\sp[0]_i_13_0 (ctl_n_23),
        .\sp_reg[0] (\sptr/p_0_in ),
        .\sp_reg[10] (rgf_n_23),
        .\sp_reg[11] (rgf_n_24),
        .\sp_reg[12] (rgf_n_25),
        .\sp_reg[13] (rgf_n_26),
        .\sp_reg[14] (rgf_n_27),
        .\sp_reg[15] (rgf_n_28),
        .\sp_reg[16] (rgf_n_29),
        .\sp_reg[17] (rgf_n_30),
        .\sp_reg[18] (rgf_n_31),
        .\sp_reg[1] (rgf_n_14),
        .\sp_reg[20] (rgf_n_33),
        .\sp_reg[22] (rgf_n_35),
        .\sp_reg[24] (rgf_n_37),
        .\sp_reg[25] (rgf_n_38),
        .\sp_reg[26] (rgf_n_39),
        .\sp_reg[2] (rgf_n_15),
        .\sp_reg[30] (rgf_n_43),
        .\sp_reg[3] (rgf_n_16),
        .\sp_reg[4] (rgf_n_17),
        .\sp_reg[5] (rgf_n_18),
        .\sp_reg[6] (rgf_n_19),
        .\sp_reg[7] (rgf_n_20),
        .\sp_reg[8] (rgf_n_21),
        .\sp_reg[9] (rgf_n_22),
        .\sr[4]_i_10_0 (rgf_n_336),
        .\sr[4]_i_10_1 (rgf_n_334),
        .\sr[4]_i_18_0 (rgf_n_452),
        .\sr[4]_i_18_1 (rgf_n_125),
        .\sr[4]_i_18_2 (rgf_n_161),
        .\sr[4]_i_18_3 (rgf_n_453),
        .\sr[4]_i_18_4 (rgf_n_127),
        .\sr[4]_i_18_5 (rgf_n_163),
        .\sr[4]_i_18_6 (rgf_n_454),
        .\sr[4]_i_18_7 (rgf_n_133),
        .\sr[4]_i_18_8 (rgf_n_165),
        .\sr[4]_i_18_9 (rgf_n_166),
        .\sr[4]_i_19 (rgf_n_451),
        .\sr[4]_i_19_0 (rgf_n_105),
        .\sr[4]_i_19_1 (rgf_n_154),
        .\sr[4]_i_20 (rgf_n_173),
        .\sr[4]_i_21 (rgf_n_175),
        .\sr[4]_i_24_0 (rgf_n_467),
        .\sr[4]_i_24_1 (rgf_n_471),
        .\sr[4]_i_24_2 (rgf_n_316),
        .\sr[4]_i_37_0 (rgf_n_134),
        .\sr[4]_i_37_1 (rgf_n_132),
        .\sr[4]_i_38 (rgf_n_109),
        .\sr[4]_i_38_0 (rgf_n_210),
        .\sr[4]_i_39_0 (rgf_n_124),
        .\sr[4]_i_40_0 (fch_n_137),
        .\sr[4]_i_40_1 (rgf_n_128),
        .\sr[4]_i_41 (rgf_n_212),
        .\sr[4]_i_43_0 (rgf_n_107),
        .\sr[4]_i_43_1 (rgf_n_104),
        .\sr[4]_i_44 (rgf_n_477),
        .\sr[4]_i_44_0 (rgf_n_216),
        .\sr[4]_i_45 (rgf_n_476),
        .\sr[4]_i_45_0 (rgf_n_220),
        .\sr[4]_i_46 (rgf_n_474),
        .\sr[4]_i_46_0 (rgf_n_211),
        .\sr[4]_i_5 (rgf_n_117),
        .\sr[4]_i_5_0 (rgf_n_158),
        .\sr[4]_i_5_1 (rgf_n_450),
        .\sr[4]_i_66_0 (rgf_n_98),
        .\sr[4]_i_66_1 (rgf_n_184),
        .\sr[4]_i_66_2 (rgf_n_244),
        .\sr[4]_i_69 (rgf_n_214),
        .\sr[4]_i_74_0 (rgf_n_229),
        .\sr[4]_i_74_1 (rgf_n_228),
        .\sr[4]_i_77 (rgf_n_183),
        .\sr[4]_i_78_0 (rgf_n_237),
        .\sr[4]_i_78_1 (rgf_n_240),
        .\sr[4]_i_7_0 (rgf_n_96),
        .\sr[4]_i_7_1 (rgf_n_310),
        .\sr[4]_i_7_2 (rgf_n_258),
        .\sr[4]_i_7_3 (rgf_n_318),
        .\sr[4]_i_7_4 (rgf_n_262),
        .\sr[4]_i_80 (rgf_n_213),
        .\sr[4]_i_81 (rgf_n_215),
        .\sr[4]_i_81_0 (rgf_n_243),
        .\sr[4]_i_81_1 (rgf_n_246),
        .\sr[4]_i_85 (rgf_n_236),
        .\sr[4]_i_85_0 (rgf_n_235),
        .\sr[4]_i_85_1 (rgf_n_223),
        .\sr[4]_i_8_0 (rgf_n_95),
        .\sr[4]_i_91_0 (rgf_n_224),
        .\sr[4]_i_91_1 (rgf_n_179),
        .\sr[4]_i_91_2 (rgf_n_253),
        .\sr[4]_i_91_3 (rgf_n_255),
        .\sr[4]_i_98 (rgf_n_256),
        .\sr[6]_i_25_0 (fch_n_86),
        .\sr[7]_i_20_0 (fch_n_154),
        .\sr[7]_i_21 (fch_n_147),
        .\sr[7]_i_4_0 (rgf_n_59),
        .\sr[7]_i_7 (rgf_n_226),
        .\sr[7]_i_7_0 (rgf_n_227),
        .\sr_reg[0] (fch_n_45),
        .\sr_reg[10] (fch_n_40),
        .\sr_reg[11] (fch_n_38),
        .\sr_reg[13] ({\sreg/p_0_in ,rgf_sr_ml,rgf_sr_dr,rgf_sr_nh,rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .\sr_reg[1] (fch_n_42),
        .\sr_reg[1]_0 (fch_n_375),
        .\sr_reg[1]_1 (fch_n_376),
        .\sr_reg[1]_10 (fch_n_385),
        .\sr_reg[1]_11 (fch_n_386),
        .\sr_reg[1]_12 (fch_n_387),
        .\sr_reg[1]_13 (fch_n_388),
        .\sr_reg[1]_14 (fch_n_389),
        .\sr_reg[1]_15 (fch_n_390),
        .\sr_reg[1]_16 (fch_n_391),
        .\sr_reg[1]_17 (fch_n_392),
        .\sr_reg[1]_18 (fch_n_393),
        .\sr_reg[1]_19 (fch_n_394),
        .\sr_reg[1]_2 (fch_n_377),
        .\sr_reg[1]_20 (fch_n_395),
        .\sr_reg[1]_21 (fch_n_396),
        .\sr_reg[1]_22 (fch_n_397),
        .\sr_reg[1]_3 (fch_n_378),
        .\sr_reg[1]_4 (fch_n_379),
        .\sr_reg[1]_5 (fch_n_380),
        .\sr_reg[1]_6 (fch_n_381),
        .\sr_reg[1]_7 (fch_n_382),
        .\sr_reg[1]_8 (fch_n_383),
        .\sr_reg[1]_9 (fch_n_384),
        .\sr_reg[2] (fch_n_43),
        .\sr_reg[3] (fch_n_44),
        .\sr_reg[4] (fch_n_11),
        .\sr_reg[4]_0 (fch_n_218),
        .\sr_reg[4]_1 (rgf_n_449),
        .\sr_reg[4]_2 (rgf_n_99),
        .\sr_reg[4]_3 (rgf_n_350),
        .\sr_reg[5] (fch_n_12),
        .\sr_reg[5]_0 (rgf_n_46),
        .\sr_reg[5]_1 (rgf_n_149),
        .\sr_reg[6] (fch_n_184),
        .\sr_reg[6]_0 (fch_n_187),
        .\sr_reg[6]_1 (fch_n_213),
        .\sr_reg[6]_2 (fch_n_223),
        .\sr_reg[6]_3 (fch_n_315),
        .\sr_reg[6]_4 (fch_n_321),
        .\sr_reg[6]_5 (fch_n_398),
        .\sr_reg[7] (fch_n_399),
        .\sr_reg[7]_0 (rgf_n_58),
        .\sr_reg[8] (fch_n_10),
        .\sr_reg[8]_0 (fch_n_41),
        .\sr_reg[8]_1 (fch_n_132),
        .\sr_reg[8]_10 (fch_n_146),
        .\sr_reg[8]_11 (fch_n_148),
        .\sr_reg[8]_12 (fch_n_149),
        .\sr_reg[8]_13 (fch_n_150),
        .\sr_reg[8]_14 (fch_n_151),
        .\sr_reg[8]_15 (fch_n_156),
        .\sr_reg[8]_16 (fch_n_157),
        .\sr_reg[8]_17 (fch_n_158),
        .\sr_reg[8]_18 (fch_n_160),
        .\sr_reg[8]_19 (fch_n_161),
        .\sr_reg[8]_2 (fch_n_138),
        .\sr_reg[8]_20 (fch_n_163),
        .\sr_reg[8]_21 (fch_n_165),
        .\sr_reg[8]_22 (fch_n_167),
        .\sr_reg[8]_23 (fch_n_168),
        .\sr_reg[8]_24 (fch_n_169),
        .\sr_reg[8]_25 (fch_n_170),
        .\sr_reg[8]_26 (fch_n_171),
        .\sr_reg[8]_27 (fch_n_172),
        .\sr_reg[8]_28 (fch_n_173),
        .\sr_reg[8]_29 (fch_n_174),
        .\sr_reg[8]_3 (fch_n_139),
        .\sr_reg[8]_30 (fch_n_175),
        .\sr_reg[8]_31 (fch_n_176),
        .\sr_reg[8]_32 (fch_n_177),
        .\sr_reg[8]_33 (fch_n_178),
        .\sr_reg[8]_34 (fch_n_180),
        .\sr_reg[8]_35 (fch_n_181),
        .\sr_reg[8]_36 (fch_n_183),
        .\sr_reg[8]_37 (fch_n_220),
        .\sr_reg[8]_38 (fch_n_316),
        .\sr_reg[8]_39 (fch_n_317),
        .\sr_reg[8]_4 (fch_n_140),
        .\sr_reg[8]_40 (fch_n_318),
        .\sr_reg[8]_41 (fch_n_319),
        .\sr_reg[8]_42 (fch_n_320),
        .\sr_reg[8]_43 (fch_n_322),
        .\sr_reg[8]_44 (fch_n_323),
        .\sr_reg[8]_45 (fch_n_324),
        .\sr_reg[8]_46 (fch_n_325),
        .\sr_reg[8]_47 (fch_n_326),
        .\sr_reg[8]_48 (fch_n_327),
        .\sr_reg[8]_49 (fch_n_328),
        .\sr_reg[8]_5 (fch_n_141),
        .\sr_reg[8]_50 (fch_n_329),
        .\sr_reg[8]_51 (fch_n_330),
        .\sr_reg[8]_52 (fch_n_331),
        .\sr_reg[8]_53 (fch_n_446),
        .\sr_reg[8]_54 (fch_n_447),
        .\sr_reg[8]_55 (fch_n_448),
        .\sr_reg[8]_56 (fch_n_449),
        .\sr_reg[8]_57 (fch_n_450),
        .\sr_reg[8]_58 (fch_n_451),
        .\sr_reg[8]_59 (fch_n_452),
        .\sr_reg[8]_6 (fch_n_142),
        .\sr_reg[8]_60 (fch_n_453),
        .\sr_reg[8]_61 (fch_n_454),
        .\sr_reg[8]_62 (fch_n_455),
        .\sr_reg[8]_63 (fch_n_456),
        .\sr_reg[8]_64 (fch_n_457),
        .\sr_reg[8]_65 (fch_n_458),
        .\sr_reg[8]_66 (fch_n_459),
        .\sr_reg[8]_67 (fch_n_495),
        .\sr_reg[8]_68 (fch_n_496),
        .\sr_reg[8]_69 (fch_n_497),
        .\sr_reg[8]_7 (fch_n_143),
        .\sr_reg[8]_70 (fch_n_498),
        .\sr_reg[8]_71 (fch_n_499),
        .\sr_reg[8]_72 ({cbus_bk2[14],cbus_bk2[10:8],cbus_bk2[6],cbus_bk2[4],cbus_bk2[2:0]}),
        .\sr_reg[8]_8 (fch_n_144),
        .\sr_reg[8]_9 (fch_n_145),
        .\stat[0]_i_2_0 (rgf_n_444),
        .\stat[1]_i_10_0 (alu_n_85),
        .\stat[1]_i_6_0 (ctl_n_5),
        .\stat_reg[0] (fch_n_87),
        .\stat_reg[0]_0 (fch_n_88),
        .\stat_reg[0]_1 (fch_n_89),
        .\stat_reg[0]_10 (ctl_n_15),
        .\stat_reg[0]_11 (rgf_n_443),
        .\stat_reg[0]_2 (fch_n_123),
        .\stat_reg[0]_3 (ccmd[4]),
        .\stat_reg[0]_4 (bcmd[3]),
        .\stat_reg[0]_5 (fch_n_263),
        .\stat_reg[0]_6 (bcmd[0]),
        .\stat_reg[0]_7 (fch_n_335),
        .\stat_reg[0]_8 (fch_n_540),
        .\stat_reg[0]_9 (fch_n_542),
        .\stat_reg[1] (bcmd[2]),
        .\stat_reg[1]_0 (rgf_n_442),
        .\stat_reg[1]_1 (ctl_n_22),
        .\stat_reg[2] (fch_n_39),
        .\stat_reg[2]_0 (cbus_sel_cr),
        .\stat_reg[2]_1 (fch_n_122),
        .\stat_reg[2]_10 (fch_n_541),
        .\stat_reg[2]_11 (fch_n_543),
        .\stat_reg[2]_12 (stat),
        .\stat_reg[2]_13 (rgf_n_438),
        .\stat_reg[2]_14 (ctl_n_4),
        .\stat_reg[2]_2 (fch_n_131),
        .\stat_reg[2]_3 (fch_n_216),
        .\stat_reg[2]_4 (fch_n_221),
        .\stat_reg[2]_5 ({fch_n_272,stat_nx}),
        .\stat_reg[2]_6 (bcmd[1]),
        .\stat_reg[2]_7 (fch_n_334),
        .\stat_reg[2]_8 (fch_n_336),
        .\stat_reg[2]_9 (fch_n_374),
        .\tr[16]_i_3_0 (rgf_n_368),
        .\tr[16]_i_7_0 (rgf_n_348),
        .\tr[16]_i_7_1 (rgf_n_305),
        .\tr[17]_i_2_0 (rgf_n_371),
        .\tr[17]_i_3 (rgf_n_208),
        .\tr[17]_i_3_0 (rgf_n_209),
        .\tr[17]_i_5_0 (rgf_n_303),
        .\tr[18]_i_2_0 (rgf_n_338),
        .\tr[18]_i_2_1 (rgf_n_363),
        .\tr[18]_i_3 (rgf_n_204),
        .\tr[18]_i_3_0 (rgf_n_205),
        .\tr[18]_i_5_0 (rgf_n_346),
        .\tr[18]_i_5_1 (rgf_n_301),
        .\tr[19]_i_14_0 (fch_n_128),
        .\tr[19]_i_3 (rgf_n_202),
        .\tr[19]_i_3_0 (rgf_n_203),
        .\tr[19]_i_5_0 (rgf_n_345),
        .\tr[19]_i_5_1 (rgf_n_300),
        .\tr[19]_i_9 (rgf_n_177),
        .\tr[20]_i_2_0 (rgf_n_364),
        .\tr[20]_i_3 (rgf_n_171),
        .\tr[20]_i_5_0 (rgf_n_344),
        .\tr[20]_i_5_1 (rgf_n_299),
        .\tr[20]_i_7 (rgf_n_232),
        .\tr[21]_i_14_0 (fch_n_124),
        .\tr[21]_i_2 (rgf_n_335),
        .\tr[21]_i_3 (rgf_n_172),
        .\tr[21]_i_5_0 (rgf_n_343),
        .\tr[21]_i_5_1 (rgf_n_298),
        .\tr[21]_i_7 (rgf_n_233),
        .\tr[22]_i_2_0 (rgf_n_365),
        .\tr[22]_i_3 (rgf_n_168),
        .\tr[22]_i_5_0 (rgf_n_342),
        .\tr[22]_i_5_1 (rgf_n_296),
        .\tr[22]_i_7_0 (rgf_n_242),
        .\tr[23]_i_15_0 (fch_n_125),
        .\tr[23]_i_2 (rgf_n_319),
        .\tr[23]_i_3 (rgf_n_199),
        .\tr[23]_i_3_0 (rgf_n_200),
        .\tr[23]_i_5_0 (rgf_n_341),
        .\tr[24]_i_2_0 (rgf_n_367),
        .\tr[24]_i_3 (rgf_n_150),
        .\tr[24]_i_5_0 (rgf_n_340),
        .\tr[24]_i_7 (rgf_n_147),
        .\tr[25]_i_2_0 (rgf_n_366),
        .\tr[25]_i_5_0 (rgf_n_339),
        .\tr[25]_i_5_1 (rgf_n_315),
        .\tr[26]_i_2_0 (rgf_n_370),
        .\tr[27]_i_14 (fch_n_126),
        .\tr[27]_i_5_0 (rgf_n_337),
        .\tr[27]_i_5_1 (rgf_n_312),
        .\tr[28]_i_13_0 (fch_n_120),
        .\tr[28]_i_3 (rgf_n_106),
        .\tr[28]_i_9_0 (rgf_n_251),
        .\tr[29]_i_14_0 (fch_n_119),
        .\tr[29]_i_7 (rgf_n_245),
        .\tr[30]_i_2_0 ({\div/rem [30],\div/rem [26:24],\div/rem [22],\div/rem [20],\div/rem [18:0]}),
        .\tr[30]_i_2_1 (rgf_n_369),
        .\tr[30]_i_8 (rgf_n_238),
        .\tr[31]_i_12_0 (rgf_n_445),
        .\tr[31]_i_44_0 (fch_n_85),
        .\tr_reg[0] (fch_n_341),
        .\tr_reg[0]_0 (rgf_n_156),
        .\tr_reg[0]_1 (rgf_n_180),
        .\tr_reg[0]_2 (rgf_n_116),
        .\tr_reg[0]_3 (mem_n_17),
        .\tr_reg[0]_4 (mem_n_26),
        .\tr_reg[10] (fch_n_351),
        .\tr_reg[10]_0 (rgf_n_157),
        .\tr_reg[10]_1 (rgf_n_119),
        .\tr_reg[11] (fch_n_352),
        .\tr_reg[11]_0 (rgf_n_153),
        .\tr_reg[11]_1 (rgf_n_103),
        .\tr_reg[11]_2 (rgf_n_201),
        .\tr_reg[12] (fch_n_353),
        .\tr_reg[12]_0 (rgf_n_115),
        .\tr_reg[13] (fch_n_354),
        .\tr_reg[13]_0 (rgf_n_112),
        .\tr_reg[13]_1 (rgf_n_113),
        .\tr_reg[14] (fch_n_355),
        .\tr_reg[14]_0 (rgf_n_162),
        .\tr_reg[14]_1 (rgf_n_126),
        .\tr_reg[15] (fch_n_356),
        .\tr_reg[15]_0 (rgf_n_178),
        .\tr_reg[15]_1 (rgf_n_145),
        .\tr_reg[15]_2 (rgf_n_185),
        .\tr_reg[15]_3 (mem_n_25),
        .\tr_reg[16] (fch_n_372),
        .\tr_reg[16]_0 (rgf_n_97),
        .\tr_reg[17] (fch_n_371),
        .\tr_reg[17]_0 (rgf_n_137),
        .\tr_reg[18] (fch_n_370),
        .\tr_reg[18]_0 (rgf_n_142),
        .\tr_reg[19] (fch_n_369),
        .\tr_reg[1] (fch_n_342),
        .\tr_reg[1]_0 (rgf_n_108),
        .\tr_reg[1]_1 (mem_n_18),
        .\tr_reg[1]_2 (mem_n_27),
        .\tr_reg[20] (fch_n_368),
        .\tr_reg[20]_0 (rgf_n_140),
        .\tr_reg[21] (fch_n_367),
        .\tr_reg[22] (fch_n_366),
        .\tr_reg[22]_0 (rgf_n_141),
        .\tr_reg[23] (fch_n_365),
        .\tr_reg[24] (fch_n_364),
        .\tr_reg[24]_0 (rgf_n_138),
        .\tr_reg[25] (fch_n_363),
        .\tr_reg[25]_0 (rgf_n_144),
        .\tr_reg[26] (fch_n_362),
        .\tr_reg[26]_0 (rgf_n_143),
        .\tr_reg[27] (fch_n_361),
        .\tr_reg[28] (fch_n_360),
        .\tr_reg[29] (fch_n_359),
        .\tr_reg[2] (fch_n_343),
        .\tr_reg[2]_0 (rgf_n_110),
        .\tr_reg[2]_1 (mem_n_19),
        .\tr_reg[2]_2 (mem_n_28),
        .\tr_reg[30] (fch_n_358),
        .\tr_reg[30]_0 (rgf_n_139),
        .\tr_reg[30]_1 (alu_n_6),
        .\tr_reg[31] (fch_n_357),
        .\tr_reg[3] (fch_n_344),
        .\tr_reg[3]_0 (rgf_n_111),
        .\tr_reg[3]_1 (rgf_n_188),
        .\tr_reg[3]_2 (mem_n_20),
        .\tr_reg[3]_3 (mem_n_29),
        .\tr_reg[4] (fch_n_345),
        .\tr_reg[4]_0 (mem_n_30),
        .\tr_reg[4]_1 (mem_n_21),
        .\tr_reg[4]_2 (rgf_n_160),
        .\tr_reg[4]_3 (rgf_n_122),
        .\tr_reg[4]_4 (rgf_n_195),
        .\tr_reg[5] (fch_n_346),
        .\tr_reg[5]_0 (rgf_n_159),
        .\tr_reg[5]_1 (rgf_n_121),
        .\tr_reg[5]_2 (rgf_n_194),
        .\tr_reg[5]_3 (mem_n_22),
        .\tr_reg[5]_4 (mem_n_31),
        .\tr_reg[6] (fch_n_347),
        .\tr_reg[6]_0 (rgf_n_135),
        .\tr_reg[6]_1 (mem_n_23),
        .\tr_reg[6]_2 (mem_n_32),
        .\tr_reg[7] (fch_n_348),
        .\tr_reg[7]_0 (rgf_n_151),
        .\tr_reg[7]_1 (rgf_n_100),
        .\tr_reg[7]_2 (rgf_n_225),
        .\tr_reg[7]_3 (mem_n_24),
        .\tr_reg[7]_4 (mem_n_33),
        .\tr_reg[8] (fch_n_349),
        .\tr_reg[8]_0 (rgf_n_123),
        .\tr_reg[8]_1 (rgf_n_206),
        .\tr_reg[9] (fch_n_350),
        .\tr_reg[9]_0 (rgf_n_164),
        .\tr_reg[9]_1 (rgf_n_131),
        .\tr_reg[9]_2 (rgf_n_207));
  niho_mem mem
       (.D({mem_n_0,mem_n_1,mem_n_2,mem_n_3,mem_n_4,mem_n_5,mem_n_6}),
        .bcmd({bcmd[2],bcmd[0]}),
        .bdatr({bdatr[31],bdatr[29:27],bdatr[23],bdatr[21],bdatr[19],bdatr[15:0]}),
        .bdatr_0_sp_1(mem_n_17),
        .bdatr_10_sp_1(mem_n_28),
        .bdatr_11_sp_1(mem_n_29),
        .bdatr_12_sp_1(mem_n_30),
        .bdatr_13_sp_1(mem_n_31),
        .bdatr_14_sp_1(mem_n_32),
        .bdatr_15_sp_1(mem_n_33),
        .bdatr_1_sp_1(mem_n_18),
        .bdatr_2_sp_1(mem_n_19),
        .bdatr_3_sp_1(mem_n_20),
        .bdatr_4_sp_1(mem_n_21),
        .bdatr_5_sp_1(mem_n_22),
        .bdatr_6_sp_1(mem_n_23),
        .bdatr_7_sp_1(mem_n_24),
        .bdatr_8_sp_1(mem_n_26),
        .bdatr_9_sp_1(mem_n_27),
        .brdy(brdy),
        .cbus_i({cbus_i[31],cbus_i[29:27],cbus_i[23],cbus_i[21],cbus_i[19]}),
        .\cbus_i[31] ({cbus[31],cbus[29:27],cbus[23],cbus[21],cbus[19]}),
        .clk(clk),
        .\grn_reg[15] ({cbus[15],cbus[13:11],cbus[7],cbus[5],cbus[3]}),
        .out(rgf_sr_nh),
        .p_0_in(p_0_in),
        .p_2_in({p_2_in[31],p_2_in[29:27],p_2_in[23],p_2_in[21],p_2_in[19]}),
        .read_cyc(read_cyc),
        .\read_cyc_reg[0] (fch_n_462),
        .\read_cyc_reg[1] (mem_n_25),
        .\sp_reg[19] (rgf_n_32),
        .\sp_reg[21] (rgf_n_34),
        .\sp_reg[23] (rgf_n_36),
        .\sp_reg[27] (cbus_sel_cr[2]),
        .\sp_reg[27]_0 (rgf_n_40),
        .\sp_reg[28] (rgf_n_41),
        .\sp_reg[29] (rgf_n_42),
        .\sp_reg[31] (rgf_n_44),
        .\sr_reg[8] ({cbus_bk2[15],cbus_bk2[13:11],cbus_bk2[7],cbus_bk2[5],cbus_bk2[3]}),
        .\tr_reg[27] (ccmd[4]));
  niho_rgf rgf
       (.D(\sreg/p_0_in__0 ),
        .E(fch_n_378),
        .O(rgf_n_45),
        .Q({\div/quo [29:27],\div/quo [23],\div/quo [21],\div/quo [19]}),
        .S({fch_n_501,fch_n_502,fch_n_503,fch_n_504}),
        .abus_0(abus_0),
        .abus_o(abus_o),
        .abus_o_16_sp_1(ccmd[4]),
        .abus_sel_0(abus_sel_0),
        .abus_sel_cr({abus_sel_cr[5],abus_sel_cr[2:0]}),
        .alu_sr_flag(alu_sr_flag),
        .\art/add/iv[7]_i_32 ({rgf_n_351,rgf_n_352,rgf_n_353,rgf_n_354}),
        .\art/add/sr[5]_i_14 ({rgf_n_47,rgf_n_48,rgf_n_49,rgf_n_50}),
        .\art/add/sr[5]_i_18 ({rgf_n_359,rgf_n_360,rgf_n_361,rgf_n_362}),
        .\badr[0]_INST_0_i_1 (rgf_n_231),
        .\badr[0]_INST_0_i_1_0 (rgf_n_318),
        .\badr[1]_INST_0_i_1 (rgf_n_316),
        .\badr[21]_INST_0_i_1 (rgf_n_60),
        .\badr[2]_INST_0_i_1 (rgf_n_471),
        .\badr[31]_INST_0_i_69 ({fch_ir[15:11],fch_ir[7]}),
        .\badr[4]_INST_0_i_1 (rgf_n_467),
        .\badr[5]_INST_0_i_1 (rgf_n_258),
        .\badr[5]_INST_0_i_1_0 (rgf_n_310),
        .\badr[6]_INST_0_i_1 (rgf_n_465),
        .bbus_0({bbus_0[13],bbus_0[8],bbus_0[4:3],bbus_0[1]}),
        .bbus_o({bbus_o[5],bbus_o[0]}),
        .bbus_sel_0(bbus_sel_0),
        .bbus_sel_cr(bbus_sel_cr),
        .bbus_sr({bbus_sr[5],bbus_sr[0]}),
        .\bdatw[8]_INST_0_i_2 (rgf_n_95),
        .cbus(cbus),
        .cbus_sel_0(cbus_sel_0),
        .clk(clk),
        .ctl_selb_0(ctl_selb_0),
        .ctl_selb_rn(ctl_selb_rn),
        .ctl_sp_dec(ctl_sp_dec),
        .ctl_sp_id4(ctl_sp_id4),
        .ctl_sp_inc(ctl_sp_inc),
        .fch_irq_req(fch_irq_req),
        .fch_pc(fch_pc),
        .\grn_reg[0] (fch_n_334),
        .\grn_reg[0]_0 (fch_n_374),
        .\grn_reg[15] (fch_n_385),
        .\grn_reg[15]_0 (fch_n_389),
        .\grn_reg[15]_1 (fch_n_393),
        .\grn_reg[15]_10 (fch_n_375),
        .\grn_reg[15]_11 (fch_n_381),
        .\grn_reg[15]_12 (fch_n_382),
        .\grn_reg[15]_13 (fch_n_386),
        .\grn_reg[15]_14 (fch_n_390),
        .\grn_reg[15]_15 (fch_n_394),
        .\grn_reg[15]_16 (fch_n_373),
        .\grn_reg[15]_17 (fch_n_379),
        .\grn_reg[15]_18 (fch_n_384),
        .\grn_reg[15]_19 (fch_n_388),
        .\grn_reg[15]_2 (fch_n_397),
        .\grn_reg[15]_20 (fch_n_392),
        .\grn_reg[15]_21 (fch_n_396),
        .\grn_reg[15]_22 (fch_n_376),
        .\grn_reg[15]_3 (fch_n_377),
        .\grn_reg[15]_4 (fch_n_380),
        .\grn_reg[15]_5 (cbus_bk2),
        .\grn_reg[15]_6 (fch_n_383),
        .\grn_reg[15]_7 (fch_n_387),
        .\grn_reg[15]_8 (fch_n_391),
        .\grn_reg[15]_9 (fch_n_395),
        .\grn_reg[1] (rgf_n_539),
        .\grn_reg[2] (rgf_n_538),
        .\grn_reg[3] (rgf_n_537),
        .\grn_reg[4] (rgf_n_261),
        .\i_/bdatw[15]_INST_0_i_27 (fch_n_336),
        .\i_/bdatw[15]_INST_0_i_27_0 (fch_n_540),
        .\i_/bdatw[15]_INST_0_i_65 (fch_n_541),
        .\i_/bdatw[15]_INST_0_i_65_0 (fch_n_223),
        .\i_/bdatw[15]_INST_0_i_65_1 (fch_n_263),
        .\i_/bdatw[15]_INST_0_i_65_2 (fch_n_543),
        .\i_/bdatw[15]_INST_0_i_67 (fch_n_542),
        .\i_/bdatw[15]_INST_0_i_67_0 (fch_n_335),
        .irq(irq),
        .irq_lev(irq_lev),
        .irq_lev_0_sp_1(rgf_n_437),
        .irq_lev_1_sp_1(rgf_n_456),
        .\iv[0]_i_10 (fch_n_148),
        .\iv[0]_i_10_0 (fch_n_153),
        .\iv[0]_i_10_1 (fch_n_159),
        .\iv[0]_i_19 (fch_n_150),
        .\iv[0]_i_25 (rgf_n_170),
        .\iv[0]_i_3 (fch_n_315),
        .\iv[0]_i_3_0 (fch_n_152),
        .\iv[0]_i_3_1 (fch_n_181),
        .\iv[0]_i_6 (fch_n_213),
        .\iv[0]_i_6_0 ({fch_n_512,fch_n_513,fch_n_514}),
        .\iv[0]_i_7 (fch_n_88),
        .\iv[10]_i_10 (rgf_n_157),
        .\iv[10]_i_2 (fch_n_166),
        .\iv[10]_i_5 (fch_n_455),
        .\iv[10]_i_9 (rgf_n_158),
        .\iv[11]_i_11 (rgf_n_153),
        .\iv[12]_i_2 (fch_n_164),
        .\iv[13]_i_10 (rgf_n_112),
        .\iv[13]_i_17 (fch_n_89),
        .\iv[13]_i_17_0 (fch_n_123),
        .\iv[13]_i_2 (fch_n_162),
        .\iv[13]_i_27 (rgf_n_125),
        .\iv[14]_i_11 (rgf_n_162),
        .\iv[14]_i_35 (rgf_n_129),
        .\iv[14]_i_49 (rgf_n_167),
        .\iv[14]_i_5 (fch_n_327),
        .\iv[15]_i_108 (rgf_n_296),
        .\iv[15]_i_108_0 (rgf_n_298),
        .\iv[15]_i_108_1 (rgf_n_299),
        .\iv[15]_i_108_10 (rgf_n_334),
        .\iv[15]_i_108_11 (rgf_n_335),
        .\iv[15]_i_108_12 (rgf_n_336),
        .\iv[15]_i_108_13 (rgf_n_337),
        .\iv[15]_i_108_14 (rgf_n_338),
        .\iv[15]_i_108_15 (rgf_n_339),
        .\iv[15]_i_108_16 (rgf_n_340),
        .\iv[15]_i_108_17 (rgf_n_341),
        .\iv[15]_i_108_18 (rgf_n_342),
        .\iv[15]_i_108_19 (rgf_n_343),
        .\iv[15]_i_108_2 (rgf_n_300),
        .\iv[15]_i_108_20 (rgf_n_344),
        .\iv[15]_i_108_21 (rgf_n_345),
        .\iv[15]_i_108_22 (rgf_n_346),
        .\iv[15]_i_108_23 (rgf_n_348),
        .\iv[15]_i_108_3 (rgf_n_301),
        .\iv[15]_i_108_4 (rgf_n_303),
        .\iv[15]_i_108_5 (rgf_n_305),
        .\iv[15]_i_108_6 (rgf_n_307),
        .\iv[15]_i_108_7 (rgf_n_312),
        .\iv[15]_i_108_8 (rgf_n_315),
        .\iv[15]_i_108_9 (rgf_n_319),
        .\iv[15]_i_8 (fch_n_449),
        .\iv[15]_i_8_0 (fch_n_322),
        .\iv[15]_i_8_1 (fch_n_158),
        .\iv[15]_i_8_2 (fch_n_448),
        .\iv[15]_i_96 (fch_n_224),
        .\iv[15]_i_96_0 (fch_n_265),
        .\iv[1]_i_10 (fch_n_317),
        .\iv[1]_i_10_0 (fch_n_185),
        .\iv[1]_i_10_1 (fch_n_194),
        .\iv[1]_i_9 (fch_n_329),
        .\iv[2]_i_9 (fch_n_459),
        .\iv[3]_i_10 (fch_n_319),
        .\iv[3]_i_10_0 (fch_n_186),
        .\iv[3]_i_10_1 (fch_n_193),
        .\iv[3]_i_9 (fch_n_328),
        .\iv[4]_i_3 (fch_n_498),
        .\iv[4]_i_35 (rgf_n_171),
        .\iv[4]_i_6 ({fch_n_509,fch_n_510,fch_n_511}),
        .\iv[4]_i_9 (fch_n_458),
        .\iv[5]_i_3 (fch_n_499),
        .\iv[5]_i_9 (fch_n_457),
        .\iv[6]_i_10 (fch_n_321),
        .\iv[6]_i_10_0 (fch_n_188),
        .\iv[6]_i_10_1 (fch_n_192),
        .\iv[7]_i_17 (rgf_n_151),
        .\iv[7]_i_25 (rgf_n_225),
        .\iv[7]_i_3 (fch_n_187),
        .\iv[7]_i_33 (rgf_n_96),
        .\iv[7]_i_7 (fch_n_130),
        .\iv[7]_i_7_0 (fch_n_217),
        .\iv[7]_i_7_1 (fch_n_129),
        .\iv[7]_i_9 (fch_n_331),
        .\iv[8]_i_2 (fch_n_154),
        .\iv[8]_i_20 (rgf_n_127),
        .\iv[8]_i_34 (rgf_n_200),
        .\iv[8]_i_5 (fch_n_456),
        .\iv[8]_i_8 ({fch_n_505,fch_n_506,fch_n_507,fch_n_508}),
        .\iv[9]_i_11 (rgf_n_164),
        .\iv[9]_i_5 (fch_n_326),
        .\iv_reg[10] (rgf_n_532),
        .\iv_reg[11] (rgf_n_531),
        .\iv_reg[12] (rgf_n_530),
        .\iv_reg[13] (rgf_n_529),
        .\iv_reg[14] (rgf_n_528),
        .\iv_reg[15] (rgf_n_479),
        .\iv_reg[15]_0 ({\ivec/p_0_in ,rgf_iv_ve}),
        .\iv_reg[6] (rgf_n_536),
        .\iv_reg[7] (rgf_n_535),
        .\iv_reg[8] (rgf_n_534),
        .\iv_reg[9] (rgf_n_533),
        .mul_a(\mul/mul_a ),
        .mul_a_i(mul_a_i),
        .\mul_a_reg[0] (fch_n_341),
        .\mul_a_reg[10] (fch_n_351),
        .\mul_a_reg[11] (fch_n_352),
        .\mul_a_reg[12] (fch_n_353),
        .\mul_a_reg[13] (fch_n_354),
        .\mul_a_reg[14] (fch_n_355),
        .\mul_a_reg[15] (fch_n_356),
        .\mul_a_reg[16] (fch_n_372),
        .\mul_a_reg[17] (fch_n_371),
        .\mul_a_reg[18] (fch_n_370),
        .\mul_a_reg[19] (fch_n_369),
        .\mul_a_reg[1] (fch_n_342),
        .\mul_a_reg[20] (fch_n_368),
        .\mul_a_reg[21] (fch_n_367),
        .\mul_a_reg[22] (fch_n_366),
        .\mul_a_reg[23] (fch_n_365),
        .\mul_a_reg[24] (fch_n_364),
        .\mul_a_reg[25] (fch_n_363),
        .\mul_a_reg[26] (fch_n_362),
        .\mul_a_reg[27] (fch_n_361),
        .\mul_a_reg[28] (fch_n_360),
        .\mul_a_reg[29] (fch_n_359),
        .\mul_a_reg[2] (fch_n_343),
        .\mul_a_reg[30] (fch_n_358),
        .\mul_a_reg[32] (fch_n_212),
        .\mul_a_reg[32]_0 (fch_n_357),
        .\mul_a_reg[3] (fch_n_344),
        .\mul_a_reg[4] (fch_n_345),
        .\mul_a_reg[5] (fch_n_346),
        .\mul_a_reg[6] (fch_n_347),
        .\mul_a_reg[7] (fch_n_348),
        .\mul_a_reg[8] (fch_n_349),
        .\mul_a_reg[9] (fch_n_350),
        .\mul_b_reg[0] (fch_n_262),
        .\mul_b_reg[0]_0 (fch_n_275),
        .\mul_b_reg[5] (fch_n_276),
        .\mul_b_reg[5]_0 (fch_n_277),
        .mul_rslt(\mul/mul_rslt ),
        .mul_rslt0(\mul/mul_rslt0 ),
        .niho_dsp_a(niho_dsp_a),
        .\niho_dsp_a[15]_INST_0_i_3 (rgf_n_262),
        .niho_dsp_b({niho_dsp_b[5],niho_dsp_b[0]}),
        .\niho_dsp_b[5] (fch_n_209),
        .\niho_dsp_b[5]_0 (alu_n_163),
        .niho_dsp_b_0_sp_1(alu_n_167),
        .niho_dsp_c({niho_dsp_c[29:27],niho_dsp_c[23],niho_dsp_c[21],niho_dsp_c[19]}),
        .out({\sreg/p_0_in ,rgf_sr_ml,rgf_sr_dr,rgf_sr_nh,rgf_sr_flag,rgf_sr_ie,sr_bank}),
        .p_0_in(p_0_in),
        .p_2_in({p_2_in[31],p_2_in[29:27],p_2_in[23],p_2_in[21],p_2_in[19]}),
        .\pc_reg[15] (\pcnt/p_1_in ),
        .\remden_reg[16] (alu_n_82),
        .\remden_reg[17] (alu_n_69),
        .\remden_reg[18] (alu_n_83),
        .\remden_reg[19] (alu_n_70),
        .\remden_reg[20] (alu_n_81),
        .\remden_reg[21] (alu_n_80),
        .\remden_reg[22] (alu_n_79),
        .\remden_reg[23] (alu_n_78),
        .\remden_reg[24] (alu_n_77),
        .\remden_reg[25] (alu_n_76),
        .\remden_reg[26] (alu_n_4),
        .\remden_reg[26]_0 (alu_n_71),
        .\remden_reg[27] (alu_n_72),
        .\remden_reg[28] (alu_n_73),
        .\remden_reg[29] (alu_n_75),
        .\remden_reg[30] (alu_n_74),
        .rgf_pc(fadr),
        .rst_n(rst_n),
        .\sp_reg[0] (\sptr/p_0_in ),
        .\sp_reg[10] (rgf_n_23),
        .\sp_reg[11] (rgf_n_24),
        .\sp_reg[12] (rgf_n_25),
        .\sp_reg[13] (rgf_n_26),
        .\sp_reg[14] (rgf_n_27),
        .\sp_reg[15] (rgf_n_28),
        .\sp_reg[16] (rgf_n_29),
        .\sp_reg[16]_0 (rgf_n_568),
        .\sp_reg[17] (rgf_n_30),
        .\sp_reg[17]_0 (rgf_n_567),
        .\sp_reg[18] (rgf_n_31),
        .\sp_reg[18]_0 (rgf_n_566),
        .\sp_reg[19] (rgf_n_32),
        .\sp_reg[19]_0 (rgf_n_565),
        .\sp_reg[1] (rgf_n_14),
        .\sp_reg[1]_0 (rgf_n_585),
        .\sp_reg[20] (rgf_n_33),
        .\sp_reg[20]_0 (rgf_n_564),
        .\sp_reg[21] (rgf_n_34),
        .\sp_reg[21]_0 (rgf_n_563),
        .\sp_reg[22] (rgf_n_35),
        .\sp_reg[22]_0 (rgf_n_562),
        .\sp_reg[23] (rgf_n_36),
        .\sp_reg[23]_0 (rgf_n_561),
        .\sp_reg[24] (rgf_n_37),
        .\sp_reg[24]_0 (rgf_n_560),
        .\sp_reg[25] (rgf_n_38),
        .\sp_reg[25]_0 (rgf_n_559),
        .\sp_reg[26] (rgf_n_39),
        .\sp_reg[26]_0 (rgf_n_558),
        .\sp_reg[27] (rgf_n_40),
        .\sp_reg[27]_0 (rgf_n_557),
        .\sp_reg[28] (rgf_n_41),
        .\sp_reg[28]_0 (rgf_n_556),
        .\sp_reg[29] (rgf_n_42),
        .\sp_reg[29]_0 (rgf_n_555),
        .\sp_reg[2] (rgf_n_15),
        .\sp_reg[2]_0 (rgf_n_586),
        .\sp_reg[30] (rgf_n_43),
        .\sp_reg[30]_0 (rgf_n_554),
        .\sp_reg[31] (rgf_n_44),
        .\sp_reg[31]_0 (rgf_n_553),
        .\sp_reg[31]_1 ({mem_n_0,fch_n_56,mem_n_1,mem_n_2,mem_n_3,fch_n_57,fch_n_58,fch_n_59,mem_n_4,fch_n_60,mem_n_5,fch_n_61,mem_n_6,fch_n_62,fch_n_63,fch_n_64,fch_n_65,fch_n_66,fch_n_67,fch_n_68,fch_n_69,fch_n_70,fch_n_71,fch_n_72,fch_n_73,fch_n_74,fch_n_75,fch_n_76,fch_n_77,fch_n_78,fch_n_79,fch_n_80}),
        .\sp_reg[3] (rgf_n_16),
        .\sp_reg[3]_0 (rgf_n_587),
        .\sp_reg[4] (rgf_n_17),
        .\sp_reg[4]_0 (rgf_n_259),
        .\sp_reg[5] (rgf_n_18),
        .\sp_reg[6] (rgf_n_19),
        .\sp_reg[7] (rgf_n_20),
        .\sp_reg[8] (rgf_n_21),
        .\sp_reg[9] (rgf_n_22),
        .\sr[4]_i_116 (rgf_n_133),
        .\sr[4]_i_139 (fch_n_190),
        .\sr[4]_i_147 (rgf_n_105),
        .\sr[4]_i_16 (fch_n_133),
        .\sr[4]_i_16_0 (fch_n_179),
        .\sr[4]_i_18 (fch_n_320),
        .\sr[4]_i_19 (fch_n_316),
        .\sr[4]_i_20 (fch_n_169),
        .\sr[4]_i_20_0 (fch_n_163),
        .\sr[4]_i_20_1 (fch_n_170),
        .\sr[4]_i_20_2 (fch_n_165),
        .\sr[4]_i_21 (rgf_n_99),
        .\sr[4]_i_21_0 (fch_n_318),
        .\sr[4]_i_21_1 (fch_n_182),
        .\sr[4]_i_3 (fch_n_218),
        .\sr[4]_i_33 (fch_n_180),
        .\sr[4]_i_35 (fch_n_454),
        .\sr[4]_i_36 (fch_n_143),
        .\sr[4]_i_37 (fch_n_155),
        .\sr[4]_i_38 (fch_n_325),
        .\sr[4]_i_39 (fch_n_167),
        .\sr[4]_i_39_0 (fch_n_500),
        .\sr[4]_i_40 (fch_n_168),
        .\sr[4]_i_40_0 (fch_n_497),
        .\sr[4]_i_41 (fch_n_184),
        .\sr[4]_i_42 (fch_n_147),
        .\sr[4]_i_43 (fch_n_149),
        .\sr[4]_i_43_0 (fch_n_330),
        .\sr[4]_i_44 (fch_n_145),
        .\sr[4]_i_44_0 (fch_n_452),
        .\sr[4]_i_44_1 (fch_n_453),
        .\sr[4]_i_45 (fch_n_450),
        .\sr[4]_i_45_0 (fch_n_451),
        .\sr[4]_i_5 (fch_n_10),
        .\sr[4]_i_5_0 (fch_n_132),
        .\sr[4]_i_5_1 (fch_n_134),
        .\sr[4]_i_5_2 (fch_n_135),
        .\sr[4]_i_61 (fch_n_160),
        .\sr[4]_i_65 (rgf_n_117),
        .\sr[4]_i_87 (fch_n_191),
        .\sr[4]_i_89 (fch_n_161),
        .\sr[5]_i_2 (fch_n_121),
        .\sr[5]_i_3 (fch_n_157),
        .\sr[6]_i_11 (fch_n_178),
        .\sr[6]_i_12 (fch_n_87),
        .\sr[6]_i_12_0 (fch_n_189),
        .\sr[6]_i_13 (rgf_n_468),
        .\sr[6]_i_4 (fch_n_219),
        .\sr_reg[0] (fch_n_45),
        .\sr_reg[10] (rgf_n_545),
        .\sr_reg[10]_0 (fch_n_40),
        .\sr_reg[11] (rgf_n_544),
        .\sr_reg[11]_0 (fch_n_38),
        .\sr_reg[12] (rgf_n_543),
        .\sr_reg[13] (rgf_n_542),
        .\sr_reg[14] (rgf_n_541),
        .\sr_reg[15] (rgf_n_540),
        .\sr_reg[15]_0 (fch_n_39),
        .\sr_reg[1] (rgf_n_552),
        .\sr_reg[1]_0 (fch_n_42),
        .\sr_reg[2] (rgf_n_551),
        .\sr_reg[2]_0 (fch_n_43),
        .\sr_reg[3] (rgf_n_550),
        .\sr_reg[3]_0 (fch_n_44),
        .\sr_reg[4] (rgf_n_260),
        .\sr_reg[4]_0 (rgf_n_441),
        .\sr_reg[4]_1 (rgf_n_443),
        .\sr_reg[4]_2 (fch_n_136),
        .\sr_reg[4]_3 (fch_n_137),
        .\sr_reg[4]_4 (fch_n_11),
        .\sr_reg[5] (rgf_n_439),
        .\sr_reg[5]_0 (rgf_n_457),
        .\sr_reg[5]_1 (fch_n_446),
        .\sr_reg[5]_2 (fch_n_12),
        .\sr_reg[6] (rgf_n_229),
        .\sr_reg[6]_0 (rgf_n_236),
        .\sr_reg[6]_1 (rgf_n_240),
        .\sr_reg[6]_10 (fch_n_86),
        .\sr_reg[6]_11 (fch_n_216),
        .\sr_reg[6]_12 (fch_n_398),
        .\sr_reg[6]_2 (rgf_n_253),
        .\sr_reg[6]_3 (rgf_n_255),
        .\sr_reg[6]_4 ({rgf_n_355,rgf_n_356,rgf_n_357,rgf_n_358}),
        .\sr_reg[6]_5 (rgf_n_444),
        .\sr_reg[6]_6 (rgf_n_458),
        .\sr_reg[6]_7 (rgf_n_459),
        .\sr_reg[6]_8 (rgf_n_460),
        .\sr_reg[6]_9 (rgf_n_549),
        .\sr_reg[6]_i_6 (fch_n_205),
        .\sr_reg[6]_i_6_0 (fch_n_206),
        .\sr_reg[6]_i_6_1 (fch_n_207),
        .\sr_reg[7] (rgf_n_438),
        .\sr_reg[7]_0 (rgf_n_440),
        .\sr_reg[7]_1 (rgf_n_442),
        .\sr_reg[7]_2 (rgf_n_445),
        .\sr_reg[7]_3 (rgf_n_548),
        .\sr_reg[7]_4 (fch_n_399),
        .\sr_reg[8] (rgf_n_46),
        .\sr_reg[8]_0 (rgf_n_58),
        .\sr_reg[8]_1 (rgf_n_59),
        .\sr_reg[8]_10 (rgf_n_107),
        .\sr_reg[8]_100 (rgf_n_221),
        .\sr_reg[8]_101 (rgf_n_222),
        .\sr_reg[8]_102 (rgf_n_223),
        .\sr_reg[8]_103 (rgf_n_224),
        .\sr_reg[8]_104 (rgf_n_226),
        .\sr_reg[8]_105 (rgf_n_227),
        .\sr_reg[8]_106 (rgf_n_228),
        .\sr_reg[8]_107 (rgf_n_230),
        .\sr_reg[8]_108 (rgf_n_232),
        .\sr_reg[8]_109 (rgf_n_233),
        .\sr_reg[8]_11 (rgf_n_108),
        .\sr_reg[8]_110 (rgf_n_234),
        .\sr_reg[8]_111 (rgf_n_235),
        .\sr_reg[8]_112 (rgf_n_237),
        .\sr_reg[8]_113 (rgf_n_238),
        .\sr_reg[8]_114 (rgf_n_239),
        .\sr_reg[8]_115 (rgf_n_241),
        .\sr_reg[8]_116 (rgf_n_242),
        .\sr_reg[8]_117 (rgf_n_243),
        .\sr_reg[8]_118 (rgf_n_244),
        .\sr_reg[8]_119 (rgf_n_245),
        .\sr_reg[8]_12 (rgf_n_109),
        .\sr_reg[8]_120 (rgf_n_246),
        .\sr_reg[8]_121 (rgf_n_247),
        .\sr_reg[8]_122 (rgf_n_248),
        .\sr_reg[8]_123 (rgf_n_249),
        .\sr_reg[8]_124 (rgf_n_250),
        .\sr_reg[8]_125 (rgf_n_251),
        .\sr_reg[8]_126 (rgf_n_252),
        .\sr_reg[8]_127 (rgf_n_254),
        .\sr_reg[8]_128 (rgf_n_256),
        .\sr_reg[8]_129 (rgf_n_257),
        .\sr_reg[8]_13 (rgf_n_110),
        .\sr_reg[8]_130 (rgf_n_297),
        .\sr_reg[8]_131 (rgf_n_302),
        .\sr_reg[8]_132 (rgf_n_304),
        .\sr_reg[8]_133 (rgf_n_306),
        .\sr_reg[8]_134 (rgf_n_308),
        .\sr_reg[8]_135 (rgf_n_309),
        .\sr_reg[8]_136 (rgf_n_311),
        .\sr_reg[8]_137 (rgf_n_313),
        .\sr_reg[8]_138 (rgf_n_314),
        .\sr_reg[8]_139 (rgf_n_317),
        .\sr_reg[8]_14 (rgf_n_111),
        .\sr_reg[8]_140 (rgf_n_347),
        .\sr_reg[8]_141 (rgf_n_350),
        .\sr_reg[8]_142 (rgf_n_363),
        .\sr_reg[8]_143 (rgf_n_364),
        .\sr_reg[8]_144 (rgf_n_365),
        .\sr_reg[8]_145 (rgf_n_366),
        .\sr_reg[8]_146 (rgf_n_367),
        .\sr_reg[8]_147 (rgf_n_368),
        .\sr_reg[8]_148 (rgf_n_369),
        .\sr_reg[8]_149 (rgf_n_370),
        .\sr_reg[8]_15 (rgf_n_113),
        .\sr_reg[8]_150 (rgf_n_371),
        .\sr_reg[8]_151 (rgf_n_446),
        .\sr_reg[8]_152 (rgf_n_449),
        .\sr_reg[8]_153 (rgf_n_450),
        .\sr_reg[8]_154 (rgf_n_451),
        .\sr_reg[8]_155 (rgf_n_452),
        .\sr_reg[8]_156 (rgf_n_453),
        .\sr_reg[8]_157 (rgf_n_454),
        .\sr_reg[8]_158 (rgf_n_461),
        .\sr_reg[8]_159 ({rgf_n_462,rgf_n_463}),
        .\sr_reg[8]_16 (rgf_n_114),
        .\sr_reg[8]_160 (rgf_n_464),
        .\sr_reg[8]_161 (rgf_n_466),
        .\sr_reg[8]_162 (rgf_n_469),
        .\sr_reg[8]_163 (rgf_n_470),
        .\sr_reg[8]_164 (rgf_n_474),
        .\sr_reg[8]_165 (rgf_n_475),
        .\sr_reg[8]_166 (rgf_n_476),
        .\sr_reg[8]_167 (rgf_n_477),
        .\sr_reg[8]_168 (rgf_n_547),
        .\sr_reg[8]_169 (fch_n_41),
        .\sr_reg[8]_17 (rgf_n_115),
        .\sr_reg[8]_18 (rgf_n_116),
        .\sr_reg[8]_19 (rgf_n_118),
        .\sr_reg[8]_2 (rgf_n_97),
        .\sr_reg[8]_20 (rgf_n_119),
        .\sr_reg[8]_21 (rgf_n_120),
        .\sr_reg[8]_22 (rgf_n_121),
        .\sr_reg[8]_23 (rgf_n_122),
        .\sr_reg[8]_24 (rgf_n_123),
        .\sr_reg[8]_25 (rgf_n_124),
        .\sr_reg[8]_26 (rgf_n_126),
        .\sr_reg[8]_27 (rgf_n_128),
        .\sr_reg[8]_28 (rgf_n_130),
        .\sr_reg[8]_29 (rgf_n_131),
        .\sr_reg[8]_3 (rgf_n_98),
        .\sr_reg[8]_30 (rgf_n_132),
        .\sr_reg[8]_31 (rgf_n_134),
        .\sr_reg[8]_32 (rgf_n_135),
        .\sr_reg[8]_33 (rgf_n_136),
        .\sr_reg[8]_34 (rgf_n_144),
        .\sr_reg[8]_35 (rgf_n_145),
        .\sr_reg[8]_36 (rgf_n_146),
        .\sr_reg[8]_37 (rgf_n_147),
        .\sr_reg[8]_38 (rgf_n_149),
        .\sr_reg[8]_39 (rgf_n_150),
        .\sr_reg[8]_4 (rgf_n_100),
        .\sr_reg[8]_40 (rgf_n_152),
        .\sr_reg[8]_41 (rgf_n_154),
        .\sr_reg[8]_42 (rgf_n_155),
        .\sr_reg[8]_43 (rgf_n_156),
        .\sr_reg[8]_44 (rgf_n_159),
        .\sr_reg[8]_45 (rgf_n_160),
        .\sr_reg[8]_46 (rgf_n_161),
        .\sr_reg[8]_47 (rgf_n_163),
        .\sr_reg[8]_48 (rgf_n_165),
        .\sr_reg[8]_49 (rgf_n_166),
        .\sr_reg[8]_5 (rgf_n_101),
        .\sr_reg[8]_50 (rgf_n_168),
        .\sr_reg[8]_51 (rgf_n_169),
        .\sr_reg[8]_52 (rgf_n_172),
        .\sr_reg[8]_53 (rgf_n_173),
        .\sr_reg[8]_54 (rgf_n_174),
        .\sr_reg[8]_55 (rgf_n_175),
        .\sr_reg[8]_56 (rgf_n_176),
        .\sr_reg[8]_57 (rgf_n_177),
        .\sr_reg[8]_58 (rgf_n_178),
        .\sr_reg[8]_59 (rgf_n_179),
        .\sr_reg[8]_6 (rgf_n_102),
        .\sr_reg[8]_60 (rgf_n_180),
        .\sr_reg[8]_61 (rgf_n_181),
        .\sr_reg[8]_62 (rgf_n_182),
        .\sr_reg[8]_63 (rgf_n_183),
        .\sr_reg[8]_64 (rgf_n_184),
        .\sr_reg[8]_65 (rgf_n_185),
        .\sr_reg[8]_66 (rgf_n_186),
        .\sr_reg[8]_67 (rgf_n_187),
        .\sr_reg[8]_68 (rgf_n_188),
        .\sr_reg[8]_69 (rgf_n_189),
        .\sr_reg[8]_7 (rgf_n_103),
        .\sr_reg[8]_70 (rgf_n_190),
        .\sr_reg[8]_71 (rgf_n_191),
        .\sr_reg[8]_72 (rgf_n_192),
        .\sr_reg[8]_73 (rgf_n_193),
        .\sr_reg[8]_74 (rgf_n_194),
        .\sr_reg[8]_75 (rgf_n_195),
        .\sr_reg[8]_76 (rgf_n_196),
        .\sr_reg[8]_77 (rgf_n_197),
        .\sr_reg[8]_78 (rgf_n_198),
        .\sr_reg[8]_79 (rgf_n_199),
        .\sr_reg[8]_8 (rgf_n_104),
        .\sr_reg[8]_80 (rgf_n_201),
        .\sr_reg[8]_81 (rgf_n_202),
        .\sr_reg[8]_82 (rgf_n_203),
        .\sr_reg[8]_83 (rgf_n_204),
        .\sr_reg[8]_84 (rgf_n_205),
        .\sr_reg[8]_85 (rgf_n_206),
        .\sr_reg[8]_86 (rgf_n_207),
        .\sr_reg[8]_87 (rgf_n_208),
        .\sr_reg[8]_88 (rgf_n_209),
        .\sr_reg[8]_89 (rgf_n_210),
        .\sr_reg[8]_9 (rgf_n_106),
        .\sr_reg[8]_90 (rgf_n_211),
        .\sr_reg[8]_91 (rgf_n_212),
        .\sr_reg[8]_92 (rgf_n_213),
        .\sr_reg[8]_93 (rgf_n_214),
        .\sr_reg[8]_94 (rgf_n_215),
        .\sr_reg[8]_95 (rgf_n_216),
        .\sr_reg[8]_96 (rgf_n_217),
        .\sr_reg[8]_97 (rgf_n_218),
        .\sr_reg[8]_98 (rgf_n_219),
        .\sr_reg[8]_99 (rgf_n_220),
        .\sr_reg[9] (rgf_n_546),
        .\stat[0]_i_6 ({stat[2],stat[0]}),
        .\stat_reg[0] (rgf_n_455),
        .\stat_reg[1] (ctl_n_19),
        .\tr[16]_i_6 (fch_n_323),
        .\tr[16]_i_6_0 (fch_n_447),
        .\tr[17]_i_2 (fch_n_176),
        .\tr[17]_i_9 (rgf_n_137),
        .\tr[18]_i_2 (fch_n_173),
        .\tr[18]_i_9 (rgf_n_142),
        .\tr[19]_i_2 (fch_n_171),
        .\tr[19]_i_2_0 (fch_n_215),
        .\tr[19]_i_2_1 (fch_n_214),
        .\tr[19]_i_3 (fch_n_151),
        .\tr[19]_i_3_0 (fch_n_140),
        .\tr[20]_i_2 (fch_n_138),
        .\tr[20]_i_3 (fch_n_174),
        .\tr[20]_i_9 (rgf_n_140),
        .\tr[21]_i_2 (fch_n_142),
        .\tr[21]_i_3 (fch_n_175),
        .\tr[22]_i_11 (fch_n_122),
        .\tr[22]_i_2 (fch_n_141),
        .\tr[22]_i_3 (fch_n_156),
        .\tr[22]_i_9 (rgf_n_141),
        .\tr[23]_i_2 (fch_n_177),
        .\tr[24]_i_10 (rgf_n_138),
        .\tr[24]_i_2 (fch_n_183),
        .\tr[24]_i_3 (fch_n_324),
        .\tr[24]_i_3_0 (fch_n_172),
        .\tr[25]_i_2 (fch_n_220),
        .\tr[26]_i_3 (fch_n_139),
        .\tr[26]_i_9 (rgf_n_143),
        .\tr[28]_i_2 (fch_n_144),
        .\tr[29]_i_2 ({\div/rem [29:27],\div/rem [23],\div/rem [21],\div/rem [19]}),
        .\tr[29]_i_3 (fch_n_496),
        .\tr[30]_i_10 (rgf_n_139),
        .\tr[30]_i_3 (fch_n_146),
        .\tr[30]_i_3_0 (fch_n_495),
        .\tr_reg[0] (cbus_sel_cr[4:3]),
        .\tr_reg[16] (rgf_n_584),
        .\tr_reg[17] (rgf_n_583),
        .\tr_reg[18] (rgf_n_582),
        .\tr_reg[19] (rgf_n_581),
        .\tr_reg[19]_0 (fch_n_128),
        .\tr_reg[1] (fch_n_131),
        .\tr_reg[1]_0 (fch_n_127),
        .\tr_reg[20] (rgf_n_580),
        .\tr_reg[21] (rgf_n_579),
        .\tr_reg[21]_0 (fch_n_124),
        .\tr_reg[22] (rgf_n_578),
        .\tr_reg[23] (rgf_n_577),
        .\tr_reg[23]_0 (fch_n_125),
        .\tr_reg[23]_i_11 (fch_n_201),
        .\tr_reg[23]_i_11_0 (fch_n_202),
        .\tr_reg[23]_i_11_1 (fch_n_203),
        .\tr_reg[23]_i_11_2 (fch_n_204),
        .\tr_reg[24] (rgf_n_576),
        .\tr_reg[25] (rgf_n_575),
        .\tr_reg[26] (rgf_n_574),
        .\tr_reg[27] (rgf_n_573),
        .\tr_reg[27]_0 (alu_n_6),
        .\tr_reg[27]_1 (fch_n_126),
        .\tr_reg[28] (rgf_n_572),
        .\tr_reg[28]_0 (fch_n_120),
        .\tr_reg[29] (rgf_n_571),
        .\tr_reg[29]_0 (fch_n_119),
        .\tr_reg[30] (rgf_n_570),
        .\tr_reg[31] ({\treg/p_0_in ,rgf_tr}),
        .\tr_reg[31]_0 (rgf_n_569),
        .\tr_reg[31]_1 (alu_n_5),
        .\tr_reg[31]_2 (fch_n_85),
        .\tr_reg[31]_i_13 (fch_n_195),
        .\tr_reg[31]_i_13_0 (fch_n_196),
        .\tr_reg[31]_i_13_1 (fch_n_197),
        .\tr_reg[31]_i_32 (fch_n_198),
        .\tr_reg[31]_i_32_0 (fch_n_199),
        .\tr_reg[31]_i_32_1 (fch_n_258),
        .\tr_reg[31]_i_32_2 (fch_n_200),
        .\tr_reg[5] ({bbus_0[5],bbus_0[0]}));
endmodule
